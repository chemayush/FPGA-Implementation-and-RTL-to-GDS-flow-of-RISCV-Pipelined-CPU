magic
tech sky130A
magscale 1 2
timestamp 1741991081
<< nwell >>
rect 1066 2159 126538 127313
<< obsli1 >>
rect 1104 2159 126500 127313
<< obsm1 >>
rect 474 2128 126854 127424
<< metal2 >>
rect 65706 129009 65762 129809
<< obsm2 >>
rect 478 128953 65650 129146
rect 65818 128953 126850 129146
rect 478 2139 126850 128953
<< metal3 >>
rect 0 119688 800 119808
rect 0 118328 800 118448
rect 0 114928 800 115048
rect 0 114248 800 114368
rect 0 112888 800 113008
rect 0 112208 800 112328
rect 0 111528 800 111648
rect 0 110168 800 110288
rect 0 109488 800 109608
rect 0 108808 800 108928
rect 0 108128 800 108248
rect 0 107448 800 107568
rect 0 106768 800 106888
rect 0 106088 800 106208
rect 0 105408 800 105528
rect 0 104728 800 104848
rect 0 104048 800 104168
rect 0 103368 800 103488
rect 0 102688 800 102808
rect 0 102008 800 102128
rect 0 101328 800 101448
rect 0 100648 800 100768
rect 0 99968 800 100088
rect 0 99288 800 99408
rect 0 98608 800 98728
rect 0 97928 800 98048
rect 0 97248 800 97368
rect 0 96568 800 96688
rect 0 95888 800 96008
rect 0 95208 800 95328
rect 0 94528 800 94648
rect 0 93848 800 93968
rect 126865 68008 127665 68128
rect 126865 14288 127665 14408
<< obsm3 >>
rect 422 119888 126865 127329
rect 880 119608 126865 119888
rect 422 118528 126865 119608
rect 880 118248 126865 118528
rect 422 115128 126865 118248
rect 880 114848 126865 115128
rect 422 114448 126865 114848
rect 880 114168 126865 114448
rect 422 113088 126865 114168
rect 880 112808 126865 113088
rect 422 112408 126865 112808
rect 880 112128 126865 112408
rect 422 111728 126865 112128
rect 880 111448 126865 111728
rect 422 110368 126865 111448
rect 880 110088 126865 110368
rect 422 109688 126865 110088
rect 880 109408 126865 109688
rect 422 109008 126865 109408
rect 880 108728 126865 109008
rect 422 108328 126865 108728
rect 880 108048 126865 108328
rect 422 107648 126865 108048
rect 880 107368 126865 107648
rect 422 106968 126865 107368
rect 880 106688 126865 106968
rect 422 106288 126865 106688
rect 880 106008 126865 106288
rect 422 105608 126865 106008
rect 880 105328 126865 105608
rect 422 104928 126865 105328
rect 880 104648 126865 104928
rect 422 104248 126865 104648
rect 880 103968 126865 104248
rect 422 103568 126865 103968
rect 880 103288 126865 103568
rect 422 102888 126865 103288
rect 880 102608 126865 102888
rect 422 102208 126865 102608
rect 880 101928 126865 102208
rect 422 101528 126865 101928
rect 880 101248 126865 101528
rect 422 100848 126865 101248
rect 880 100568 126865 100848
rect 422 100168 126865 100568
rect 880 99888 126865 100168
rect 422 99488 126865 99888
rect 880 99208 126865 99488
rect 422 98808 126865 99208
rect 880 98528 126865 98808
rect 422 98128 126865 98528
rect 880 97848 126865 98128
rect 422 97448 126865 97848
rect 880 97168 126865 97448
rect 422 96768 126865 97168
rect 880 96488 126865 96768
rect 422 96088 126865 96488
rect 880 95808 126865 96088
rect 422 95408 126865 95808
rect 880 95128 126865 95408
rect 422 94728 126865 95128
rect 880 94448 126865 94728
rect 422 94048 126865 94448
rect 880 93768 126865 94048
rect 422 68208 126865 93768
rect 422 67928 126785 68208
rect 422 14488 126865 67928
rect 422 14208 126785 14488
rect 422 2143 126865 14208
<< metal4 >>
rect 4208 2128 4528 127344
rect 4868 2128 5188 127344
rect 34928 2128 35248 127344
rect 35588 2128 35908 127344
rect 65648 2128 65968 127344
rect 66308 2128 66628 127344
rect 96368 2128 96688 127344
rect 97028 2128 97348 127344
<< obsm4 >>
rect 342 3979 4128 127125
rect 4608 3979 4788 127125
rect 5268 3979 34848 127125
rect 35328 3979 35508 127125
rect 35988 3979 65568 127125
rect 66048 3979 66228 127125
rect 66708 3979 96288 127125
rect 96768 3979 96948 127125
rect 97428 3979 125245 127125
<< metal5 >>
rect 1056 97914 126548 98234
rect 1056 97254 126548 97574
rect 1056 67278 126548 67598
rect 1056 66618 126548 66938
rect 1056 36642 126548 36962
rect 1056 35982 126548 36302
rect 1056 6006 126548 6326
rect 1056 5346 126548 5666
<< obsm5 >>
rect 300 98554 122612 124940
rect 300 96934 736 98554
rect 300 67918 122612 96934
rect 300 66298 736 67918
rect 300 37282 122612 66298
rect 300 35662 736 37282
rect 300 19900 122612 35662
<< labels >>
rlabel metal3 s 0 93848 800 93968 6 Instr[0]
port 1 nsew signal output
rlabel metal3 s 0 112208 800 112328 6 Instr[10]
port 2 nsew signal output
rlabel metal3 s 0 99288 800 99408 6 Instr[11]
port 3 nsew signal output
rlabel metal3 s 0 97928 800 98048 6 Instr[12]
port 4 nsew signal output
rlabel metal3 s 0 99968 800 100088 6 Instr[13]
port 5 nsew signal output
rlabel metal3 s 0 106768 800 106888 6 Instr[14]
port 6 nsew signal output
rlabel metal3 s 0 105408 800 105528 6 Instr[15]
port 7 nsew signal output
rlabel metal3 s 0 114928 800 115048 6 Instr[16]
port 8 nsew signal output
rlabel metal3 s 0 98608 800 98728 6 Instr[17]
port 9 nsew signal output
rlabel metal3 s 0 112888 800 113008 6 Instr[18]
port 10 nsew signal output
rlabel metal3 s 0 95888 800 96008 6 Instr[19]
port 11 nsew signal output
rlabel metal3 s 0 96568 800 96688 6 Instr[1]
port 12 nsew signal output
rlabel metal3 s 0 114248 800 114368 6 Instr[20]
port 13 nsew signal output
rlabel metal3 s 0 118328 800 118448 6 Instr[21]
port 14 nsew signal output
rlabel metal3 s 0 111528 800 111648 6 Instr[22]
port 15 nsew signal output
rlabel metal3 s 0 119688 800 119808 6 Instr[23]
port 16 nsew signal output
rlabel metal3 s 0 103368 800 103488 6 Instr[24]
port 17 nsew signal output
rlabel metal3 s 0 110168 800 110288 6 Instr[25]
port 18 nsew signal output
rlabel metal3 s 0 108128 800 108248 6 Instr[26]
port 19 nsew signal output
rlabel metal3 s 0 104048 800 104168 6 Instr[27]
port 20 nsew signal output
rlabel metal3 s 0 95208 800 95328 6 Instr[28]
port 21 nsew signal output
rlabel metal3 s 0 101328 800 101448 6 Instr[29]
port 22 nsew signal output
rlabel metal3 s 0 94528 800 94648 6 Instr[2]
port 23 nsew signal output
rlabel metal3 s 0 102008 800 102128 6 Instr[30]
port 24 nsew signal output
rlabel metal3 s 0 102688 800 102808 6 Instr[31]
port 25 nsew signal output
rlabel metal3 s 0 97248 800 97368 6 Instr[3]
port 26 nsew signal output
rlabel metal3 s 0 109488 800 109608 6 Instr[4]
port 27 nsew signal output
rlabel metal3 s 0 104728 800 104848 6 Instr[5]
port 28 nsew signal output
rlabel metal3 s 0 106088 800 106208 6 Instr[6]
port 29 nsew signal output
rlabel metal3 s 0 108808 800 108928 6 Instr[7]
port 30 nsew signal output
rlabel metal3 s 0 100648 800 100768 6 Instr[8]
port 31 nsew signal output
rlabel metal3 s 0 107448 800 107568 6 Instr[9]
port 32 nsew signal output
rlabel metal4 s 4868 2128 5188 127344 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 35588 2128 35908 127344 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 66308 2128 66628 127344 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 97028 2128 97348 127344 6 VGND
port 33 nsew ground bidirectional
rlabel metal5 s 1056 6006 126548 6326 6 VGND
port 33 nsew ground bidirectional
rlabel metal5 s 1056 36642 126548 36962 6 VGND
port 33 nsew ground bidirectional
rlabel metal5 s 1056 67278 126548 67598 6 VGND
port 33 nsew ground bidirectional
rlabel metal5 s 1056 97914 126548 98234 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 4208 2128 4528 127344 6 VPWR
port 34 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 127344 6 VPWR
port 34 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 127344 6 VPWR
port 34 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 127344 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1056 5346 126548 5666 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1056 35982 126548 36302 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1056 66618 126548 66938 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1056 97254 126548 97574 6 VPWR
port 34 nsew power bidirectional
rlabel metal3 s 126865 14288 127665 14408 6 clk
port 35 nsew signal input
rlabel metal3 s 126865 68008 127665 68128 6 correct
port 36 nsew signal output
rlabel metal2 s 65706 129009 65762 129809 6 reset
port 37 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 127665 129809
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 57131082
string GDS_FILE /openlane/designs/pl_riscv_cpu/runs/RUN_2025.03.14_21.47.52/results/signoff/pl_riscv_cpu.magic.gds
string GDS_START 1239800
<< end >>

