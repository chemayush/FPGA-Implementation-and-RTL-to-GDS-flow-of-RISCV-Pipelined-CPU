* NGSPICE file created from pl_riscv_cpu.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtn_1 abstract view
.subckt sky130_fd_sc_hd__dlxtn_1 D GATE_N VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_2 abstract view
.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_2 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_1 abstract view
.subckt sky130_fd_sc_hd__clkinv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_4 abstract view
.subckt sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

.subckt pl_riscv_cpu Instr[0] Instr[10] Instr[11] Instr[12] Instr[13] Instr[14] Instr[15]
+ Instr[16] Instr[17] Instr[18] Instr[19] Instr[1] Instr[20] Instr[21] Instr[22] Instr[23]
+ Instr[24] Instr[25] Instr[26] Instr[27] Instr[28] Instr[29] Instr[2] Instr[30] Instr[31]
+ Instr[3] Instr[4] Instr[5] Instr[6] Instr[7] Instr[8] Instr[9] VGND VPWR clk correct
+ reset
XFILLER_0_193_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18869_ _05473_ _05619_ VGND VGND VPWR VPWR _06212_ sky130_fd_sc_hd__or2b_1
XFILLER_0_20_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20900_ datamem.data_ram\[12\]\[22\] _07833_ VGND VGND VPWR VPWR _08190_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_2_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21880_ _08795_ _09111_ _09113_ _09115_ VGND VGND VPWR VPWR _09116_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_171_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20831_ _06796_ _08111_ _08114_ _08120_ VGND VGND VPWR VPWR _08121_ sky130_fd_sc_hd__a31o_1
X_32817_ clknet_leaf_234_clk _04239_ VGND VGND VPWR VPWR datamem.data_ram\[12\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20762_ datamem.data_ram\[1\]\[6\] _06997_ _08051_ _06604_ VGND VGND VPWR VPWR _08052_
+ sky130_fd_sc_hd__a211o_1
X_23550_ clknet_1_0__leaf__10172_ VGND VGND VPWR VPWR _10174_ sky130_fd_sc_hd__buf_1
XFILLER_0_193_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32748_ clknet_leaf_233_clk _04170_ VGND VGND VPWR VPWR datamem.data_ram\[15\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_212_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22501_ rvcpu.dp.rf.reg_file_arr\[28\]\[10\] rvcpu.dp.rf.reg_file_arr\[30\]\[10\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[10\] rvcpu.dp.rf.reg_file_arr\[31\]\[10\] _09483_
+ _09656_ VGND VGND VPWR VPWR _09657_ sky130_fd_sc_hd__mux4_1
X_20693_ datamem.data_ram\[57\]\[5\] _06949_ _07982_ _07983_ VGND VGND VPWR VPWR _07984_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_174_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32679_ clknet_leaf_183_clk _04101_ VGND VGND VPWR VPWR datamem.data_ram\[18\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_25220_ _10849_ VGND VGND VPWR VPWR _02660_ sky130_fd_sc_hd__clkbuf_1
X_22432_ _09534_ _09591_ VGND VGND VPWR VPWR _09592_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25151_ _10762_ net3278 _10802_ VGND VGND VPWR VPWR _10808_ sky130_fd_sc_hd__mux2_1
X_22363_ _09510_ _09515_ _09519_ _09524_ _09525_ VGND VGND VPWR VPWR _09526_ sky130_fd_sc_hd__a311o_2
X_23573__195 clknet_1_1__leaf__10176_ VGND VGND VPWR VPWR net321 sky130_fd_sc_hd__inv_2
XFILLER_0_27_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21314_ _08575_ VGND VGND VPWR VPWR _08576_ sky130_fd_sc_hd__clkbuf_4
X_25082_ _10772_ VGND VGND VPWR VPWR _02599_ sky130_fd_sc_hd__clkbuf_1
X_24167__9 clknet_1_0__leaf__10264_ VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__inv_2
X_22294_ _09442_ _09450_ _09455_ _09458_ VGND VGND VPWR VPWR _09459_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_14_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28910_ _12960_ VGND VGND VPWR VPWR _04239_ sky130_fd_sc_hd__clkbuf_1
Xhold340 datamem.data_ram\[60\]\[0\] VGND VGND VPWR VPWR net1490 sky130_fd_sc_hd__dlygate4sd3_1
X_21245_ _08498_ _08501_ _08504_ _08507_ VGND VGND VPWR VPWR _08508_ sky130_fd_sc_hd__or4_1
X_29890_ net268 _01625_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[17\]\[21\] sky130_fd_sc_hd__dfxtp_1
Xhold351 datamem.data_ram\[21\]\[6\] VGND VGND VPWR VPWR net1501 sky130_fd_sc_hd__dlygate4sd3_1
Xhold362 datamem.data_ram\[14\]\[5\] VGND VGND VPWR VPWR net1512 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold373 datamem.data_ram\[4\]\[4\] VGND VGND VPWR VPWR net1523 sky130_fd_sc_hd__dlygate4sd3_1
X_23037__738 clknet_1_1__leaf__10089_ VGND VGND VPWR VPWR net864 sky130_fd_sc_hd__inv_2
Xhold384 datamem.data_ram\[33\]\[7\] VGND VGND VPWR VPWR net1534 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28841_ _12734_ net3632 net69 VGND VGND VPWR VPWR _12924_ sky130_fd_sc_hd__mux2_1
X_21176_ _08408_ _08464_ _06911_ VGND VGND VPWR VPWR _08465_ sky130_fd_sc_hd__mux2_1
Xhold395 datamem.data_ram\[12\]\[3\] VGND VGND VPWR VPWR net1545 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_225_5893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20127_ datamem.data_ram\[3\]\[27\] _06863_ _06620_ datamem.data_ram\[4\]\[27\] _07419_
+ VGND VGND VPWR VPWR _07420_ sky130_fd_sc_hd__o221a_1
X_28772_ _12601_ _10960_ _12886_ VGND VGND VPWR VPWR _12887_ sky130_fd_sc_hd__a21oi_4
X_25984_ _13903_ _11268_ VGND VGND VPWR VPWR _11316_ sky130_fd_sc_hd__nand2_1
X_27723_ _12300_ VGND VGND VPWR VPWR _03712_ sky130_fd_sc_hd__clkbuf_1
X_20058_ datamem.data_ram\[46\]\[26\] _06743_ _07242_ datamem.data_ram\[41\]\[26\]
+ _07351_ VGND VGND VPWR VPWR _07352_ sky130_fd_sc_hd__o221a_1
X_24935_ _10480_ net2478 net91 VGND VGND VPWR VPWR _10686_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1040 datamem.data_ram\[45\]\[15\] VGND VGND VPWR VPWR net2190 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_137_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1051 rvcpu.dp.rf.reg_file_arr\[30\]\[29\] VGND VGND VPWR VPWR net2201 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1062 datamem.data_ram\[60\]\[31\] VGND VGND VPWR VPWR net2212 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_159_4310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27654_ _12263_ VGND VGND VPWR VPWR _03680_ sky130_fd_sc_hd__clkbuf_1
Xhold1073 datamem.data_ram\[47\]\[23\] VGND VGND VPWR VPWR net2223 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_159_4321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24866_ _10400_ net3668 _10641_ VGND VGND VPWR VPWR _10649_ sky130_fd_sc_hd__mux2_1
Xhold1084 datamem.data_ram\[3\]\[22\] VGND VGND VPWR VPWR net2234 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_202 _09482_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1095 datamem.data_ram\[37\]\[13\] VGND VGND VPWR VPWR net2245 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_213 _09725_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26605_ _10520_ _11123_ _10998_ VGND VGND VPWR VPWR _11650_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_200_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_224 _10057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27585_ _12226_ VGND VGND VPWR VPWR _03648_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_235 _10268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_4207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24797_ _10500_ VGND VGND VPWR VPWR _10611_ sky130_fd_sc_hd__buf_6
XANTENNA_246 _11972_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_0__10205_ _10205_ VGND VGND VPWR VPWR clknet_0__10205_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_95_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_4218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_257 _13200_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_1_1__f__10105_ clknet_0__10105_ VGND VGND VPWR VPWR clknet_1_1__leaf__10105_
+ sky130_fd_sc_hd__clkbuf_16
X_29324_ clknet_leaf_0_clk _01059_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD1E\[31\] sky130_fd_sc_hd__dfxtp_1
X_26536_ _11081_ _11610_ VGND VGND VPWR VPWR _11612_ sky130_fd_sc_hd__and2_1
XFILLER_0_138_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_268 _13229_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_279 _13251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__10136_ _10136_ VGND VGND VPWR VPWR clknet_0__10136_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_83_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29255_ _09255_ net3186 _13141_ VGND VGND VPWR VPWR _13148_ sky130_fd_sc_hd__mux2_1
X_26467_ _11576_ _11236_ _11540_ _06538_ _11589_ VGND VGND VPWR VPWR _11590_ sky130_fd_sc_hd__a221o_1
XFILLER_0_67_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16220_ _14465_ VGND VGND VPWR VPWR _01927_ sky130_fd_sc_hd__clkbuf_1
X_28206_ _12460_ net4247 net46 VGND VGND VPWR VPWR _12571_ sky130_fd_sc_hd__mux2_1
X_25418_ _10758_ net2283 _10961_ VGND VGND VPWR VPWR _10965_ sky130_fd_sc_hd__mux2_1
X_29186_ _13110_ VGND VGND VPWR VPWR _04365_ sky130_fd_sc_hd__clkbuf_1
X_26398_ _13517_ _11153_ _11538_ _11541_ _10780_ VGND VGND VPWR VPWR _03146_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_192_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28137_ _12534_ VGND VGND VPWR VPWR _03892_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_114_3225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16151_ _14418_ VGND VGND VPWR VPWR _01949_ sky130_fd_sc_hd__clkbuf_1
X_25349_ _10325_ _10921_ _10922_ VGND VGND VPWR VPWR _10923_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_114_3236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15102_ _13353_ _13644_ _13645_ _13646_ _13412_ VGND VGND VPWR VPWR _13647_ sky130_fd_sc_hd__a221o_1
XFILLER_0_180_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_210_52 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16082_ net2868 _13275_ _14348_ VGND VGND VPWR VPWR _14382_ sky130_fd_sc_hd__mux2_1
X_28068_ _12367_ net3061 _12492_ VGND VGND VPWR VPWR _12498_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_185_4926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_185_4937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15033_ _13573_ _13576_ _13579_ _13423_ _13466_ VGND VGND VPWR VPWR _13580_ sky130_fd_sc_hd__o221a_1
X_27019_ _07791_ _11109_ _11839_ VGND VGND VPWR VPWR _11896_ sky130_fd_sc_hd__or3_1
X_19910_ datamem.data_ram\[46\]\[17\] _06628_ _06829_ datamem.data_ram\[43\]\[17\]
+ VGND VGND VPWR VPWR _07205_ sky130_fd_sc_hd__o22a_1
XFILLER_0_146_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30030_ net392 _01765_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[13\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_19841_ _06989_ VGND VGND VPWR VPWR _07136_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_43_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_219_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24168__10 clknet_1_1__leaf__10264_ VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__inv_2
X_23860__423 clknet_1_0__leaf__10219_ VGND VGND VPWR VPWR net549 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_88_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19772_ _06967_ _07064_ _07066_ VGND VGND VPWR VPWR _07067_ sky130_fd_sc_hd__and3_1
X_16984_ _04744_ VGND VGND VPWR VPWR _01550_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_88_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18723_ _05693_ _05944_ _05820_ VGND VGND VPWR VPWR _06075_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_155_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_3955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15935_ _14303_ VGND VGND VPWR VPWR _02058_ sky130_fd_sc_hd__clkbuf_1
X_31981_ clknet_leaf_138_clk _03403_ VGND VGND VPWR VPWR datamem.data_ram\[53\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_14 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18654_ _06004_ _06008_ _06009_ VGND VGND VPWR VPWR _06010_ sky130_fd_sc_hd__and3_1
X_30932_ clknet_leaf_154_clk _02667_ VGND VGND VPWR VPWR datamem.data_ram\[40\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_24183__24 clknet_1_0__leaf__10265_ VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__inv_2
X_15866_ _14265_ VGND VGND VPWR VPWR _02089_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_188_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14817_ _13369_ VGND VGND VPWR VPWR _13370_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_203_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17605_ _13260_ net3109 _05068_ VGND VGND VPWR VPWR _05074_ sky130_fd_sc_hd__mux2_1
XFILLER_0_192_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18585_ _05676_ _05943_ VGND VGND VPWR VPWR _05944_ sky130_fd_sc_hd__or2_2
X_30863_ clknet_leaf_264_clk _02598_ VGND VGND VPWR VPWR datamem.data_ram\[43\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_188_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15797_ _14228_ VGND VGND VPWR VPWR _02129_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_188_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_47_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17536_ _05037_ VGND VGND VPWR VPWR _01275_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32602_ clknet_leaf_266_clk _04024_ VGND VGND VPWR VPWR datamem.data_ram\[20\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_14748_ _13300_ VGND VGND VPWR VPWR _13301_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_58_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_103_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30794_ clknet_leaf_180_clk _02529_ VGND VGND VPWR VPWR datamem.data_ram\[46\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_103_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32533_ clknet_leaf_244_clk _03955_ VGND VGND VPWR VPWR datamem.data_ram\[23\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_17467_ _14181_ net3401 _04996_ VGND VGND VPWR VPWR _05001_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14679_ _13243_ VGND VGND VPWR VPWR _13244_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_11_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19206_ rvcpu.dp.plde.ImmExtE\[24\] rvcpu.dp.plde.PCE\[24\] VGND VGND VPWR VPWR _06515_
+ sky130_fd_sc_hd__or2_1
X_16418_ _14575_ VGND VGND VPWR VPWR _01831_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_184_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32464_ clknet_leaf_182_clk _03886_ VGND VGND VPWR VPWR datamem.data_ram\[26\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_17398_ _04964_ VGND VGND VPWR VPWR _01340_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_884 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31415_ clknet_leaf_53_clk _03118_ VGND VGND VPWR VPWR datamem.data_ram\[15\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_19137_ _06454_ VGND VGND VPWR VPWR rvcpu.dp.lAuiPCE\[15\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16349_ net2298 _14447_ _14536_ VGND VGND VPWR VPWR _14539_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32395_ clknet_leaf_77_clk _03817_ VGND VGND VPWR VPWR datamem.data_ram\[29\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19068_ rvcpu.dp.plde.ImmExtE\[7\] rvcpu.dp.plde.PCE\[7\] VGND VGND VPWR VPWR _06394_
+ sky130_fd_sc_hd__nand2_1
X_31346_ clknet_leaf_19_clk _03049_ VGND VGND VPWR VPWR rvcpu.dp.plde.ALUControlE\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18019_ _05384_ _05385_ _05388_ VGND VGND VPWR VPWR _05389_ sky130_fd_sc_hd__nand3_1
XFILLER_0_11_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31277_ clknet_leaf_126_clk _02980_ VGND VGND VPWR VPWR datamem.data_ram\[24\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__10125_ clknet_0__10125_ VGND VGND VPWR VPWR clknet_1_0__leaf__10125_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_61_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21030_ datamem.data_ram\[17\]\[31\] _06944_ _07838_ VGND VGND VPWR VPWR _08319_
+ sky130_fd_sc_hd__o21a_1
X_30228_ net582 _01963_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[7\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_226_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30159_ net521 _01894_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[0\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_226_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24720_ _10478_ net3743 net59 VGND VGND VPWR VPWR _10568_ sky130_fd_sc_hd__mux2_1
X_21932_ _08725_ _09164_ VGND VGND VPWR VPWR _09165_ sky130_fd_sc_hd__nor2_1
XFILLER_0_179_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24651_ _10529_ VGND VGND VPWR VPWR _02411_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_195_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21863_ _08510_ _09099_ VGND VGND VPWR VPWR _09100_ sky130_fd_sc_hd__nor2_1
XFILLER_0_171_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20814_ datamem.data_ram\[56\]\[30\] _06934_ VGND VGND VPWR VPWR _08104_ sky130_fd_sc_hd__or2_1
X_27370_ _12103_ VGND VGND VPWR VPWR _03556_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21794_ rvcpu.dp.rf.reg_file_arr\[4\]\[21\] rvcpu.dp.rf.reg_file_arr\[5\]\[21\] rvcpu.dp.rf.reg_file_arr\[6\]\[21\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[21\] _08839_ _08840_ VGND VGND VPWR VPWR _09035_
+ sky130_fd_sc_hd__mux4_1
X_24582_ _10385_ net3229 _10491_ VGND VGND VPWR VPWR _10492_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26321_ _11493_ VGND VGND VPWR VPWR _03117_ sky130_fd_sc_hd__clkbuf_1
X_20745_ _08032_ _08034_ VGND VGND VPWR VPWR _08035_ sky130_fd_sc_hd__and2_1
XFILLER_0_163_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_886 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29040_ _13018_ net1812 _13030_ _13033_ VGND VGND VPWR VPWR _04296_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_189_5026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_4104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_174_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26252_ _11438_ _11458_ _11459_ net1176 VGND VGND VPWR VPWR _03082_ sky130_fd_sc_hd__a2bb2o_1
X_20676_ datamem.data_ram\[40\]\[5\] _07138_ _06977_ datamem.data_ram\[44\]\[5\] _07966_
+ VGND VGND VPWR VPWR _07967_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_189_5037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25203_ _10840_ VGND VGND VPWR VPWR _02652_ sky130_fd_sc_hd__clkbuf_1
X_22415_ rvcpu.dp.rf.reg_file_arr\[16\]\[6\] rvcpu.dp.rf.reg_file_arr\[17\]\[6\] rvcpu.dp.rf.reg_file_arr\[18\]\[6\]
+ rvcpu.dp.rf.reg_file_arr\[19\]\[6\] _09512_ _09513_ VGND VGND VPWR VPWR _09575_
+ sky130_fd_sc_hd__mux4_2
X_26183_ _11428_ VGND VGND VPWR VPWR _03044_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23395_ _10148_ VGND VGND VPWR VPWR _01536_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25134_ _10476_ net3117 net87 VGND VGND VPWR VPWR _10799_ sky130_fd_sc_hd__mux2_1
X_22346_ _09501_ _09505_ _09509_ _09491_ VGND VGND VPWR VPWR _01126_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_227_5933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_227_5944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_227_5955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25065_ _09251_ VGND VGND VPWR VPWR _10762_ sky130_fd_sc_hd__buf_2
X_29942_ net312 _01677_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[15\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_22277_ _09411_ VGND VGND VPWR VPWR _09442_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_148_4044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_4055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21228_ datamem.data_ram\[53\]\[14\] datamem.data_ram\[52\]\[14\] datamem.data_ram\[52\]\[7\]
+ datamem.data_ram\[53\]\[7\] VGND VGND VPWR VPWR _08491_ sky130_fd_sc_hd__or4_1
XFILLER_0_218_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold170 datamem.data_ram\[43\]\[2\] VGND VGND VPWR VPWR net1320 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_180_4812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold181 datamem.data_ram\[44\]\[7\] VGND VGND VPWR VPWR net1331 sky130_fd_sc_hd__dlygate4sd3_1
X_29873_ net251 _01608_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[17\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_180_4823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold192 datamem.data_ram\[4\]\[7\] VGND VGND VPWR VPWR net1342 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28824_ _12751_ net2349 _12914_ VGND VGND VPWR VPWR _12915_ sky130_fd_sc_hd__mux2_1
X_21159_ datamem.data_ram\[2\]\[23\] datamem.data_ram\[3\]\[23\] _07912_ VGND VGND
+ VPWR VPWR _08448_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_6_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23998__532 clknet_1_0__leaf__10240_ VGND VGND VPWR VPWR net658 sky130_fd_sc_hd__inv_2
X_28755_ _12687_ net3237 _12877_ VGND VGND VPWR VPWR _12878_ sky130_fd_sc_hd__mux2_1
X_25967_ net4409 _11302_ _11300_ _11306_ VGND VGND VPWR VPWR _02950_ sky130_fd_sc_hd__o211a_1
XFILLER_0_219_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27706_ _12291_ VGND VGND VPWR VPWR _03704_ sky130_fd_sc_hd__clkbuf_1
X_15720_ _14184_ VGND VGND VPWR VPWR _02162_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_107_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24918_ _10400_ net3210 _10669_ VGND VGND VPWR VPWR _10677_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28686_ _12279_ _12622_ _12795_ VGND VGND VPWR VPWR _12841_ sky130_fd_sc_hd__a21oi_1
X_25898_ net1807 _11263_ VGND VGND VPWR VPWR _11267_ sky130_fd_sc_hd__or2_1
XFILLER_0_213_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27637_ _12130_ net3135 _12251_ VGND VGND VPWR VPWR _12254_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15651_ _14137_ net4395 _14131_ VGND VGND VPWR VPWR _14138_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_178_4763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24849_ _10639_ VGND VGND VPWR VPWR _02499_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_178_4774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_201_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14602_ _13185_ VGND VGND VPWR VPWR _03202_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_200_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18370_ _05282_ _05732_ _05734_ VGND VGND VPWR VPWR _05735_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_115_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27568_ _12217_ VGND VGND VPWR VPWR _03640_ sky130_fd_sc_hd__clkbuf_1
X_15582_ _14098_ VGND VGND VPWR VPWR _02214_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_205_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29307_ clknet_leaf_0_clk _01042_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD1E\[14\] sky130_fd_sc_hd__dfxtp_1
X_17321_ _04923_ VGND VGND VPWR VPWR _01384_ sky130_fd_sc_hd__clkbuf_1
X_26519_ _10780_ _11604_ VGND VGND VPWR VPWR _11605_ sky130_fd_sc_hd__nor2_2
XFILLER_0_185_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27499_ _12145_ net2188 _12179_ VGND VGND VPWR VPWR _12181_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17252_ _04886_ VGND VGND VPWR VPWR _01416_ sky130_fd_sc_hd__clkbuf_1
X_29238_ _09325_ net3323 _13132_ VGND VGND VPWR VPWR _13139_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_3781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16203_ net3399 _14453_ _14443_ VGND VGND VPWR VPWR _14454_ sky130_fd_sc_hd__mux2_1
XFILLER_0_221_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_3792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29169_ _13101_ VGND VGND VPWR VPWR _04357_ sky130_fd_sc_hd__clkbuf_1
X_17183_ _14170_ net2793 _04840_ VGND VGND VPWR VPWR _04850_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_854 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31200_ clknet_leaf_29_clk _02903_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCPlus4D\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_3678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16134_ net1963 _13251_ _14407_ VGND VGND VPWR VPWR _14410_ sky130_fd_sc_hd__mux2_1
X_32180_ clknet_leaf_161_clk _03602_ VGND VGND VPWR VPWR datamem.data_ram\[37\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_133_3689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31131_ clknet_leaf_125_clk _02866_ VGND VGND VPWR VPWR datamem.data_ram\[25\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_16065_ _14373_ VGND VGND VPWR VPWR _01990_ sky130_fd_sc_hd__clkbuf_1
X_15016_ _13333_ _13563_ VGND VGND VPWR VPWR _13564_ sky130_fd_sc_hd__or2_1
X_31062_ clknet_leaf_273_clk _02797_ VGND VGND VPWR VPWR datamem.data_ram\[8\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_209_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_202_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30013_ net375 _01748_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[13\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_19824_ _07096_ _07118_ VGND VGND VPWR VPWR _07119_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_36_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_209_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_208_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1809 datamem.data_ram\[0\]\[27\] VGND VGND VPWR VPWR net2959 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19755_ datamem.data_ram\[56\]\[25\] _06807_ _06726_ datamem.data_ram\[63\]\[25\]
+ _07049_ VGND VGND VPWR VPWR _07050_ sky130_fd_sc_hd__o221a_1
XFILLER_0_120_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16967_ _04735_ VGND VGND VPWR VPWR _01558_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_223_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18706_ _05878_ _06058_ _05697_ VGND VGND VPWR VPWR _06059_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15918_ _14294_ VGND VGND VPWR VPWR _02066_ sky130_fd_sc_hd__clkbuf_1
X_19686_ datamem.data_ram\[61\]\[0\] _06969_ _06980_ _06981_ VGND VGND VPWR VPWR _06982_
+ sky130_fd_sc_hd__a211o_1
X_31964_ clknet_leaf_122_clk _03386_ VGND VGND VPWR VPWR datamem.data_ram\[28\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_16898_ net2243 _14449_ _04695_ VGND VGND VPWR VPWR _04699_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18637_ _05346_ _05594_ _05956_ VGND VGND VPWR VPWR _05994_ sky130_fd_sc_hd__and3_1
X_30915_ clknet_leaf_172_clk _02650_ VGND VGND VPWR VPWR datamem.data_ram\[41\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_15849_ _14256_ VGND VGND VPWR VPWR _02097_ sky130_fd_sc_hd__clkbuf_1
X_31895_ _04415_ net118 VGND VGND VPWR VPWR datamem.rd_data_mem\[0\] sky130_fd_sc_hd__dlxtn_1
XFILLER_0_189_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30846_ clknet_leaf_216_clk _02581_ VGND VGND VPWR VPWR datamem.data_ram\[43\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_18568_ _05692_ _05925_ _05927_ _05750_ VGND VGND VPWR VPWR _05928_ sky130_fd_sc_hd__a211o_1
XFILLER_0_91_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17519_ _05028_ VGND VGND VPWR VPWR _01283_ sky130_fd_sc_hd__clkbuf_1
X_18499_ _05383_ _05397_ _05238_ VGND VGND VPWR VPWR _05861_ sky130_fd_sc_hd__o21a_1
X_30777_ clknet_leaf_220_clk _02512_ VGND VGND VPWR VPWR datamem.data_ram\[46\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20530_ _07820_ VGND VGND VPWR VPWR _07821_ sky130_fd_sc_hd__buf_6
X_32516_ clknet_leaf_169_clk _03938_ VGND VGND VPWR VPWR datamem.data_ram\[24\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32447_ clknet_leaf_81_clk _03869_ VGND VGND VPWR VPWR datamem.data_ram\[27\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_20461_ datamem.data_ram\[18\]\[20\] _06611_ _06782_ datamem.data_ram\[17\]\[20\]
+ VGND VGND VPWR VPWR _07753_ sky130_fd_sc_hd__o22a_1
XFILLER_0_132_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22200_ _09273_ net2952 _09371_ VGND VGND VPWR VPWR _09373_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32378_ clknet_leaf_160_clk _03800_ VGND VGND VPWR VPWR datamem.data_ram\[2\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_20392_ datamem.data_ram\[26\]\[28\] _06689_ _06661_ datamem.data_ram\[29\]\[28\]
+ VGND VGND VPWR VPWR _07684_ sky130_fd_sc_hd__o22a_1
X_23867__429 clknet_1_1__leaf__10220_ VGND VGND VPWR VPWR net555 sky130_fd_sc_hd__inv_2
XFILLER_0_3_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22131_ _09240_ net4371 _09332_ VGND VGND VPWR VPWR _09335_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31329_ clknet_leaf_16_clk _03032_ VGND VGND VPWR VPWR rvcpu.dp.plde.RdE\[0\] sky130_fd_sc_hd__dfxtp_1
X_22062_ _09280_ VGND VGND VPWR VPWR _01071_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__10108_ clknet_0__10108_ VGND VGND VPWR VPWR clknet_1_0__leaf__10108_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_100_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21013_ datamem.data_ram\[56\]\[31\] _06811_ _06812_ datamem.data_ram\[59\]\[31\]
+ _08301_ VGND VGND VPWR VPWR _08302_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_222_5830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26870_ _11795_ net1471 _11797_ _11805_ VGND VGND VPWR VPWR _03354_ sky130_fd_sc_hd__a31o_1
XFILLER_0_227_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25821_ rvcpu.dp.pcreg.q\[21\] rvcpu.dp.pcreg.q\[20\] _11200_ VGND VGND VPWR VPWR
+ _11208_ sky130_fd_sc_hd__and3_1
XFILLER_0_215_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28540_ _09251_ VGND VGND VPWR VPWR _12762_ sky130_fd_sc_hd__buf_2
X_25752_ net2400 _11155_ VGND VGND VPWR VPWR _11156_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24703_ _10452_ net3439 _10552_ VGND VGND VPWR VPWR _10559_ sky130_fd_sc_hd__mux2_1
X_28471_ _12456_ net3193 _12713_ VGND VGND VPWR VPWR _12718_ sky130_fd_sc_hd__mux2_1
X_21915_ rvcpu.dp.rf.reg_file_arr\[28\]\[28\] rvcpu.dp.rf.reg_file_arr\[30\]\[28\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[28\] rvcpu.dp.rf.reg_file_arr\[31\]\[28\] _08533_
+ _08536_ VGND VGND VPWR VPWR _09149_ sky130_fd_sc_hd__mux4_2
X_25683_ _10268_ _11112_ _10052_ VGND VGND VPWR VPWR _11113_ sky130_fd_sc_hd__and3_2
X_22895_ _09516_ _10027_ _10029_ _09404_ VGND VGND VPWR VPWR _10030_ sky130_fd_sc_hd__o211a_1
XFILLER_0_195_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27422_ _12133_ VGND VGND VPWR VPWR _03578_ sky130_fd_sc_hd__clkbuf_1
X_24634_ _07136_ VGND VGND VPWR VPWR _10520_ sky130_fd_sc_hd__buf_8
X_21846_ rvcpu.dp.rf.reg_file_arr\[12\]\[24\] rvcpu.dp.rf.reg_file_arr\[13\]\[24\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[24\] rvcpu.dp.rf.reg_file_arr\[15\]\[24\] _08578_
+ _08684_ VGND VGND VPWR VPWR _09084_ sky130_fd_sc_hd__mux4_2
XFILLER_0_77_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27353_ _12093_ net2365 _12081_ VGND VGND VPWR VPWR _12094_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_216_5678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24565_ _10439_ net3202 _10482_ VGND VGND VPWR VPWR _10483_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_216_5689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21777_ _08695_ _09018_ VGND VGND VPWR VPWR _09019_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_176_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26304_ net1843 _11478_ VGND VGND VPWR VPWR _11485_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23516_ _10166_ VGND VGND VPWR VPWR _01639_ sky130_fd_sc_hd__clkbuf_1
X_27284_ _11965_ _12054_ VGND VGND VPWR VPWR _12055_ sky130_fd_sc_hd__and2_1
X_20728_ datamem.data_ram\[30\]\[6\] datamem.data_ram\[31\]\[6\] _07837_ VGND VGND
+ VPWR VPWR _08018_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24496_ _10438_ VGND VGND VPWR VPWR _02347_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29023_ _13023_ VGND VGND VPWR VPWR _04289_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26235_ _11379_ _03031_ _11454_ VGND VGND VPWR VPWR _03068_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_137_Right_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20659_ datamem.data_ram\[45\]\[29\] _07037_ _07948_ _07949_ VGND VGND VPWR VPWR
+ _07950_ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_12_Left_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_208_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26166_ net4449 _11408_ VGND VGND VPWR VPWR _11420_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25117_ _10735_ net3121 net88 VGND VGND VPWR VPWR _10790_ sky130_fd_sc_hd__mux2_1
X_22329_ rvcpu.dp.rf.reg_file_arr\[20\]\[2\] rvcpu.dp.rf.reg_file_arr\[21\]\[2\] rvcpu.dp.rf.reg_file_arr\[22\]\[2\]
+ rvcpu.dp.rf.reg_file_arr\[23\]\[2\] _09445_ _09447_ VGND VGND VPWR VPWR _09493_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_72_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26097_ _11383_ VGND VGND VPWR VPWR _03002_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_72_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24065__592 clknet_1_1__leaf__10247_ VGND VGND VPWR VPWR net718 sky130_fd_sc_hd__inv_2
XFILLER_0_209_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29925_ net295 _01660_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[16\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_25048_ _10750_ VGND VGND VPWR VPWR _02587_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_167_4497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_178_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_109_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17870_ rvcpu.dp.plde.Rs1E\[4\] rvcpu.dp.plem.RdM\[4\] VGND VGND VPWR VPWR _05243_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_109_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29856_ net234 _01591_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[18\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_28807_ _12687_ net3335 _12905_ VGND VGND VPWR VPWR _12906_ sky130_fd_sc_hd__mux2_1
X_16821_ net3868 _14440_ _04648_ VGND VGND VPWR VPWR _04658_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26999_ _07019_ _10918_ _10897_ VGND VGND VPWR VPWR _11884_ sky130_fd_sc_hd__or3_1
X_29787_ net1133 _01522_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[20\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_21_Left_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16752_ _04621_ VGND VGND VPWR VPWR _01667_ sky130_fd_sc_hd__clkbuf_1
X_19540_ _06753_ _06819_ _06712_ _06835_ VGND VGND VPWR VPWR _06836_ sky130_fd_sc_hd__o211a_1
X_28738_ _12734_ net3161 net41 VGND VGND VPWR VPWR _12869_ sky130_fd_sc_hd__mux2_1
XFILLER_0_191_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15703_ _14130_ VGND VGND VPWR VPWR _14173_ sky130_fd_sc_hd__buf_4
XFILLER_0_186_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19471_ datamem.data_ram\[52\]\[16\] _06766_ _06699_ datamem.data_ram\[49\]\[16\]
+ VGND VGND VPWR VPWR _06767_ sky130_fd_sc_hd__o22a_1
X_28669_ _12279_ _12612_ _12795_ VGND VGND VPWR VPWR _12832_ sky130_fd_sc_hd__a21oi_4
X_16683_ _14147_ net4289 _04576_ VGND VGND VPWR VPWR _04585_ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30700_ clknet_leaf_147_clk _02435_ VGND VGND VPWR VPWR datamem.data_ram\[4\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_18422_ _05722_ rvcpu.dp.plde.ALUControlE\[0\] rvcpu.dp.plde.ALUControlE\[1\] VGND
+ VGND VPWR VPWR _05786_ sky130_fd_sc_hd__or3b_4
X_15634_ _14125_ VGND VGND VPWR VPWR _02189_ sky130_fd_sc_hd__clkbuf_1
X_31680_ clknet_leaf_13_clk net1255 VGND VGND VPWR VPWR rvcpu.dp.plmw.ALUResultW\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_185_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_139_3821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_139_3832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18353_ _05698_ _05701_ _05703_ _05717_ VGND VGND VPWR VPWR _05718_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_139_3843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30631_ clknet_leaf_197_clk _02366_ VGND VGND VPWR VPWR datamem.data_ram\[51\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_15565_ _13573_ _13796_ _13499_ VGND VGND VPWR VPWR _14088_ sky130_fd_sc_hd__or3_1
XFILLER_0_111_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17304_ net2068 _13216_ _04913_ VGND VGND VPWR VPWR _04915_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_620 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18284_ _05648_ _05287_ VGND VGND VPWR VPWR _05649_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_135_3729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30562_ clknet_leaf_217_clk _02297_ VGND VGND VPWR VPWR datamem.data_ram\[54\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_15496_ _14021_ _14022_ _14023_ VGND VGND VPWR VPWR _14024_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32301_ clknet_leaf_166_clk _03723_ VGND VGND VPWR VPWR datamem.data_ram\[32\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_30_Left_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17235_ _14154_ net3991 _04876_ VGND VGND VPWR VPWR _04878_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_104_Right_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_226_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30493_ clknet_leaf_144_clk _02228_ VGND VGND VPWR VPWR datamem.data_ram\[57\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32232_ clknet_leaf_169_clk _03654_ VGND VGND VPWR VPWR datamem.data_ram\[35\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17166_ _04841_ VGND VGND VPWR VPWR _01457_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23254__901 clknet_1_0__leaf__10127_ VGND VGND VPWR VPWR net1027 sky130_fd_sc_hd__inv_2
Xhold906 datamem.data_ram\[38\]\[15\] VGND VGND VPWR VPWR net2056 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16117_ net2176 _13226_ _14396_ VGND VGND VPWR VPWR _14401_ sky130_fd_sc_hd__mux2_1
Xhold917 rvcpu.dp.rf.reg_file_arr\[3\]\[13\] VGND VGND VPWR VPWR net2067 sky130_fd_sc_hd__dlygate4sd3_1
Xhold928 rvcpu.dp.pcreg.q\[19\] VGND VGND VPWR VPWR net2078 sky130_fd_sc_hd__dlygate4sd3_1
X_32163_ clknet_leaf_243_clk _03585_ VGND VGND VPWR VPWR datamem.data_ram\[38\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_38_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17097_ _14151_ net2218 _04804_ VGND VGND VPWR VPWR _04805_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold939 datamem.data_ram\[44\]\[31\] VGND VGND VPWR VPWR net2089 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31114_ clknet_leaf_58_clk _02849_ VGND VGND VPWR VPWR datamem.data_ram\[43\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_16048_ _14364_ VGND VGND VPWR VPWR _01998_ sky130_fd_sc_hd__clkbuf_1
Xhold3008 datamem.data_ram\[59\]\[20\] VGND VGND VPWR VPWR net4158 sky130_fd_sc_hd__dlygate4sd3_1
X_32094_ clknet_leaf_237_clk _03516_ VGND VGND VPWR VPWR datamem.data_ram\[8\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3019 datamem.data_ram\[23\]\[10\] VGND VGND VPWR VPWR net4169 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31045_ clknet_leaf_234_clk _02780_ VGND VGND VPWR VPWR datamem.data_ram\[9\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2307 datamem.data_ram\[56\]\[13\] VGND VGND VPWR VPWR net3457 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2318 datamem.data_ram\[26\]\[28\] VGND VGND VPWR VPWR net3468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2329 rvcpu.dp.rf.reg_file_arr\[0\]\[17\] VGND VGND VPWR VPWR net3479 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1606 rvcpu.dp.rf.reg_file_arr\[17\]\[27\] VGND VGND VPWR VPWR net2756 sky130_fd_sc_hd__dlygate4sd3_1
X_19807_ datamem.data_ram\[6\]\[9\] _06719_ _06697_ datamem.data_ram\[0\]\[9\] _07101_
+ VGND VGND VPWR VPWR _07102_ sky130_fd_sc_hd__o221a_1
XFILLER_0_224_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1617 rvcpu.dp.rf.reg_file_arr\[31\]\[22\] VGND VGND VPWR VPWR net2767 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1628 datamem.data_ram\[10\]\[12\] VGND VGND VPWR VPWR net2778 sky130_fd_sc_hd__dlygate4sd3_1
X_17999_ _05276_ rvcpu.dp.plde.ImmExtE\[3\] VGND VGND VPWR VPWR _05369_ sky130_fd_sc_hd__or2_1
Xhold1639 datamem.data_ram\[16\]\[21\] VGND VGND VPWR VPWR net2789 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_224_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19738_ datamem.data_ram\[2\]\[25\] _07023_ _07030_ _07032_ VGND VGND VPWR VPWR _07033_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_212_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19669_ _06603_ _06939_ _06957_ _06964_ VGND VGND VPWR VPWR _06965_ sky130_fd_sc_hd__o31a_1
X_31947_ clknet_leaf_117_clk _03369_ VGND VGND VPWR VPWR datamem.data_ram\[32\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21700_ _08835_ _08945_ VGND VGND VPWR VPWR _08946_ sky130_fd_sc_hd__or2_1
XFILLER_0_220_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22680_ rvcpu.dp.rf.reg_file_arr\[8\]\[19\] rvcpu.dp.rf.reg_file_arr\[10\]\[19\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[19\] rvcpu.dp.rf.reg_file_arr\[11\]\[19\] _09608_
+ _09656_ VGND VGND VPWR VPWR _09827_ sky130_fd_sc_hd__mux4_1
X_31878_ clknet_leaf_113_clk _03332_ VGND VGND VPWR VPWR datamem.data_ram\[56\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21631_ _08672_ _08872_ _08876_ _08880_ VGND VGND VPWR VPWR _08881_ sky130_fd_sc_hd__and4_1
X_30829_ clknet_leaf_155_clk _02564_ VGND VGND VPWR VPWR datamem.data_ram\[44\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24350_ _10352_ VGND VGND VPWR VPWR _02287_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21562_ _08813_ _08814_ _08689_ VGND VGND VPWR VPWR _08815_ sky130_fd_sc_hd__a21o_1
XFILLER_0_142_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_211_5553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20513_ datamem.data_ram\[56\]\[21\] _06649_ _06621_ datamem.data_ram\[60\]\[21\]
+ VGND VGND VPWR VPWR _07804_ sky130_fd_sc_hd__o22a_1
XFILLER_0_144_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_211_5564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24281_ _10313_ VGND VGND VPWR VPWR _02257_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_160_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21493_ _08515_ _08747_ _08748_ VGND VGND VPWR VPWR _08749_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_209_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26020_ net1300 _11329_ _11325_ _11335_ VGND VGND VPWR VPWR _02974_ sky130_fd_sc_hd__o211a_1
XFILLER_0_7_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20444_ _06715_ _07719_ _07724_ _06860_ _07735_ VGND VGND VPWR VPWR _07736_ sky130_fd_sc_hd__o311a_1
XFILLER_0_43_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20375_ datamem.data_ram\[43\]\[28\] _06828_ _07663_ _07666_ VGND VGND VPWR VPWR
+ _07667_ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_207_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload90 clknet_leaf_71_clk VGND VGND VPWR VPWR clkload90/X sky130_fd_sc_hd__clkbuf_4
X_22114_ _09322_ net3138 _09302_ VGND VGND VPWR VPWR _09323_ sky130_fd_sc_hd__mux2_1
X_27971_ _09251_ VGND VGND VPWR VPWR _12441_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_219_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_228_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26922_ _10043_ VGND VGND VPWR VPWR _11839_ sky130_fd_sc_hd__buf_2
X_29710_ net1056 _01445_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[22\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_22045_ _09266_ VGND VGND VPWR VPWR _09267_ sky130_fd_sc_hd__buf_2
XFILLER_0_100_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2830 datamem.data_ram\[47\]\[28\] VGND VGND VPWR VPWR net3980 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26853_ _11781_ net1827 _11785_ _11794_ VGND VGND VPWR VPWR _03348_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_162_4372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29641_ net987 _01376_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[24\]\[4\] sky130_fd_sc_hd__dfxtp_1
Xhold2841 rvcpu.dp.rf.reg_file_arr\[23\]\[20\] VGND VGND VPWR VPWR net3991 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2852 rvcpu.dp.rf.reg_file_arr\[26\]\[20\] VGND VGND VPWR VPWR net4002 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_162_4383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_162_4394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2863 rvcpu.dp.rf.reg_file_arr\[29\]\[3\] VGND VGND VPWR VPWR net4013 sky130_fd_sc_hd__dlygate4sd3_1
X_25804_ rvcpu.dp.pcreg.q\[17\] _11191_ VGND VGND VPWR VPWR _11195_ sky130_fd_sc_hd__or2_1
Xhold2874 datamem.data_ram\[11\]\[24\] VGND VGND VPWR VPWR net4024 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2885 datamem.data_ram\[48\]\[18\] VGND VGND VPWR VPWR net4035 sky130_fd_sc_hd__dlygate4sd3_1
X_29572_ net926 _01307_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[26\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_26784_ _11753_ net1532 _11748_ _11754_ VGND VGND VPWR VPWR _03319_ sky130_fd_sc_hd__a31o_1
XFILLER_0_173_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2896 datamem.data_ram\[3\]\[11\] VGND VGND VPWR VPWR net4046 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28523_ _12750_ VGND VGND VPWR VPWR _04062_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_218_5718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25735_ _11141_ VGND VGND VPWR VPWR _02883_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_218_5729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22947_ _10056_ net1509 _10046_ _10074_ VGND VGND VPWR VPWR _01162_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_175_4700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_206_Right_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28454_ _12439_ net3634 _12704_ VGND VGND VPWR VPWR _12709_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25666_ _11085_ net1814 _11097_ _11101_ VGND VGND VPWR VPWR _02854_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_65_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22878_ rvcpu.dp.rf.reg_file_arr\[0\]\[30\] rvcpu.dp.rf.reg_file_arr\[1\]\[30\] rvcpu.dp.rf.reg_file_arr\[2\]\[30\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[30\] _09477_ _09383_ VGND VGND VPWR VPWR _10014_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_156_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_121_3390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27405_ _12122_ VGND VGND VPWR VPWR _03572_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_171_4608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24617_ _10209_ _10337_ _10501_ VGND VGND VPWR VPWR _10511_ sky130_fd_sc_hd__a21oi_4
X_28385_ _06591_ VGND VGND VPWR VPWR _12668_ sky130_fd_sc_hd__clkbuf_16
X_21829_ _08835_ _09067_ VGND VGND VPWR VPWR _09068_ sky130_fd_sc_hd__or2_1
X_25597_ _10416_ _11055_ VGND VGND VPWR VPWR _11062_ sky130_fd_sc_hd__and2_1
XFILLER_0_155_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_182_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15350_ _13438_ _13879_ _13882_ _13884_ _13885_ VGND VGND VPWR VPWR _13886_ sky130_fd_sc_hd__o32a_1
X_23735__326 clknet_1_0__leaf__10199_ VGND VGND VPWR VPWR net452 sky130_fd_sc_hd__inv_2
X_27336_ _12082_ VGND VGND VPWR VPWR _03543_ sky130_fd_sc_hd__clkbuf_1
X_24548_ _10471_ VGND VGND VPWR VPWR _02366_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15281_ _13816_ _13817_ _13819_ _13521_ VGND VGND VPWR VPWR _13820_ sky130_fd_sc_hd__a31o_1
X_27267_ _10814_ net3583 _12043_ VGND VGND VPWR VPWR _12045_ sky130_fd_sc_hd__mux2_1
X_24479_ _10429_ VGND VGND VPWR VPWR _02339_ sky130_fd_sc_hd__clkbuf_1
X_29006_ _10063_ _13010_ VGND VGND VPWR VPWR _13014_ sky130_fd_sc_hd__and2_1
XFILLER_0_163_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17020_ net2500 _14434_ _04757_ VGND VGND VPWR VPWR _04764_ sky130_fd_sc_hd__mux2_1
X_26218_ net1306 _11436_ _11444_ VGND VGND VPWR VPWR _11447_ sky130_fd_sc_hd__and3_1
XFILLER_0_163_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_3604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_3615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27198_ _11965_ _12008_ VGND VGND VPWR VPWR _12009_ sky130_fd_sc_hd__and2_1
XFILLER_0_22_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_4548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_3626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_169_4559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26149_ net1962 _11408_ VGND VGND VPWR VPWR _11411_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_95_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18971_ _05305_ _05555_ VGND VGND VPWR VPWR _06307_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_131_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17922_ rvcpu.dp.plem.ALUResultM\[29\] _05293_ _05294_ _13186_ VGND VGND VPWR VPWR
+ _05295_ sky130_fd_sc_hd__o22a_1
X_29908_ clknet_leaf_146_clk _01643_ VGND VGND VPWR VPWR datamem.data_ram\[59\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26514__2 clknet_1_1__leaf__10080_ VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__inv_2
XFILLER_0_186_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_3566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_3577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17853_ _13250_ rvcpu.dp.plde.RD2E\[9\] _05194_ VGND VGND VPWR VPWR _05230_ sky130_fd_sc_hd__mux2_1
X_29839_ net217 _01574_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[18\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16804_ _04649_ VGND VGND VPWR VPWR _01635_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_195_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32850_ clknet_leaf_212_clk _04272_ VGND VGND VPWR VPWR datamem.data_ram\[11\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_14996_ _13474_ _13490_ _13543_ _13327_ VGND VGND VPWR VPWR _13544_ sky130_fd_sc_hd__o211a_1
X_17784_ _05179_ _05180_ rvcpu.dp.plde.RD2E\[1\] VGND VGND VPWR VPWR _05181_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_206_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23284__927 clknet_1_1__leaf__10131_ VGND VGND VPWR VPWR net1053 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_50_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31801_ clknet_leaf_97_clk _03255_ VGND VGND VPWR VPWR datamem.data_ram\[46\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_19523_ _06776_ _06801_ _06809_ _06818_ VGND VGND VPWR VPWR _06819_ sky130_fd_sc_hd__a31o_1
XFILLER_0_163_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16735_ net4238 _14420_ _04612_ VGND VGND VPWR VPWR _04613_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32781_ clknet_leaf_163_clk _04203_ VGND VGND VPWR VPWR datamem.data_ram\[14\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_23896__455 clknet_1_0__leaf__10223_ VGND VGND VPWR VPWR net581 sky130_fd_sc_hd__inv_2
XFILLER_0_117_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_220_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19454_ _06585_ rvcpu.dp.plem.ALUResultM\[6\] VGND VGND VPWR VPWR _06750_ sky130_fd_sc_hd__nand2_8
X_16666_ _04575_ VGND VGND VPWR VPWR _04576_ sky130_fd_sc_hd__clkbuf_4
X_31732_ net181 _03190_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[9\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_24115__622 clknet_1_1__leaf__10259_ VGND VGND VPWR VPWR net748 sky130_fd_sc_hd__inv_2
X_18405_ _05683_ VGND VGND VPWR VPWR _05769_ sky130_fd_sc_hd__clkbuf_4
X_15617_ net2409 _13251_ _14114_ VGND VGND VPWR VPWR _14117_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31663_ clknet_leaf_67_clk net1286 VGND VGND VPWR VPWR rvcpu.dp.plmw.ALUResultW\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_16597_ _04538_ _04465_ VGND VGND VPWR VPWR _04539_ sky130_fd_sc_hd__nand2_2
X_19385_ _06680_ VGND VGND VPWR VPWR _06681_ sky130_fd_sc_hd__buf_6
XFILLER_0_186_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_227_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15548_ _13501_ _14029_ VGND VGND VPWR VPWR _14073_ sky130_fd_sc_hd__nor2_1
X_30614_ clknet_leaf_148_clk _02349_ VGND VGND VPWR VPWR datamem.data_ram\[52\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_18336_ _05699_ _05700_ _05677_ VGND VGND VPWR VPWR _05701_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31594_ clknet_leaf_52_clk net1231 VGND VGND VPWR VPWR rvcpu.dp.plmw.PCPlus4W\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18267_ rvcpu.dp.plde.RD1E\[25\] _05564_ _05526_ VGND VGND VPWR VPWR _05632_ sky130_fd_sc_hd__o21ai_1
X_30545_ clknet_leaf_146_clk _02280_ VGND VGND VPWR VPWR datamem.data_ram\[55\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_15479_ _13690_ _13292_ _13693_ VGND VGND VPWR VPWR _14008_ sky130_fd_sc_hd__or3b_1
XFILLER_0_142_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_150_clk clknet_5_28__leaf_clk VGND VGND VPWR VPWR clknet_leaf_150_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_72_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17218_ _14137_ net3218 _04865_ VGND VGND VPWR VPWR _04869_ sky130_fd_sc_hd__mux2_1
X_18198_ _05486_ _05487_ VGND VGND VPWR VPWR _05563_ sky130_fd_sc_hd__or2b_1
X_30476_ net154 _02211_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[19\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold703 datamem.data_ram\[9\]\[2\] VGND VGND VPWR VPWR net1853 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold714 rvcpu.dp.plfd.InstrD\[7\] VGND VGND VPWR VPWR net1864 sky130_fd_sc_hd__dlygate4sd3_1
X_17149_ _04832_ VGND VGND VPWR VPWR _01465_ sky130_fd_sc_hd__clkbuf_1
X_32215_ clknet_leaf_269_clk _03637_ VGND VGND VPWR VPWR datamem.data_ram\[36\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold725 datamem.data_ram\[62\]\[15\] VGND VGND VPWR VPWR net1875 sky130_fd_sc_hd__dlygate4sd3_1
Xhold736 rvcpu.dp.rf.reg_file_arr\[19\]\[30\] VGND VGND VPWR VPWR net1886 sky130_fd_sc_hd__dlygate4sd3_1
Xhold747 rvcpu.dp.plfd.PCPlus4D\[26\] VGND VGND VPWR VPWR net1897 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20160_ datamem.data_ram\[29\]\[27\] _06724_ _06810_ _07452_ VGND VGND VPWR VPWR
+ _07453_ sky130_fd_sc_hd__o211a_1
X_32146_ clknet_leaf_229_clk _03568_ VGND VGND VPWR VPWR datamem.data_ram\[38\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold758 rvcpu.dp.rf.reg_file_arr\[17\]\[28\] VGND VGND VPWR VPWR net1908 sky130_fd_sc_hd__dlygate4sd3_1
Xhold769 rvcpu.dp.rf.reg_file_arr\[7\]\[0\] VGND VGND VPWR VPWR net1919 sky130_fd_sc_hd__dlygate4sd3_1
X_24161__664 clknet_1_1__leaf__10263_ VGND VGND VPWR VPWR net790 sky130_fd_sc_hd__inv_2
X_32077_ clknet_leaf_94_clk _03499_ VGND VGND VPWR VPWR datamem.data_ram\[33\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_20091_ datamem.data_ram\[58\]\[10\] _06689_ _06668_ datamem.data_ram\[63\]\[10\]
+ VGND VGND VPWR VPWR _07385_ sky130_fd_sc_hd__o22a_1
Xhold2104 datamem.data_ram\[26\]\[20\] VGND VGND VPWR VPWR net3254 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2115 rvcpu.dp.rf.reg_file_arr\[18\]\[1\] VGND VGND VPWR VPWR net3265 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2126 datamem.data_ram\[23\]\[14\] VGND VGND VPWR VPWR net3276 sky130_fd_sc_hd__dlygate4sd3_1
X_31028_ clknet_leaf_73_clk _02763_ VGND VGND VPWR VPWR datamem.data_ram\[40\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2137 datamem.data_ram\[43\]\[12\] VGND VGND VPWR VPWR net3287 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2148 datamem.data_ram\[53\]\[23\] VGND VGND VPWR VPWR net3298 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1403 rvcpu.dp.rf.reg_file_arr\[29\]\[12\] VGND VGND VPWR VPWR net2553 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1414 rvcpu.dp.rf.reg_file_arr\[17\]\[0\] VGND VGND VPWR VPWR net2564 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2159 datamem.data_ram\[58\]\[11\] VGND VGND VPWR VPWR net3309 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_204_5390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1425 datamem.data_ram\[19\]\[21\] VGND VGND VPWR VPWR net2575 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1436 datamem.data_ram\[35\]\[12\] VGND VGND VPWR VPWR net2586 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1447 rvcpu.dp.rf.reg_file_arr\[31\]\[0\] VGND VGND VPWR VPWR net2597 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1458 rvcpu.dp.rf.reg_file_arr\[0\]\[2\] VGND VGND VPWR VPWR net2608 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1469 rvcpu.dp.rf.reg_file_arr\[14\]\[28\] VGND VGND VPWR VPWR net2619 sky130_fd_sc_hd__dlygate4sd3_1
X_22801_ rvcpu.dp.rf.reg_file_arr\[24\]\[26\] rvcpu.dp.rf.reg_file_arr\[25\]\[26\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[26\] rvcpu.dp.rf.reg_file_arr\[27\]\[26\] _09484_
+ _09431_ VGND VGND VPWR VPWR _09941_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_200_5287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_200_5298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_196_5191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32979_ clknet_leaf_267_clk _04401_ VGND VGND VPWR VPWR datamem.data_ram\[63\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_20993_ _06641_ _08280_ _08281_ _06922_ VGND VGND VPWR VPWR _08282_ sky130_fd_sc_hd__o22a_1
XFILLER_0_149_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25520_ _10991_ net1505 _11009_ _11016_ VGND VGND VPWR VPWR _02793_ sky130_fd_sc_hd__a31o_1
X_22732_ rvcpu.dp.rf.reg_file_arr\[12\]\[22\] rvcpu.dp.rf.reg_file_arr\[13\]\[22\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[22\] rvcpu.dp.rf.reg_file_arr\[15\]\[22\] _09386_
+ _09419_ VGND VGND VPWR VPWR _09876_ sky130_fd_sc_hd__mux4_1
XFILLER_0_149_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_213_5604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25451_ _10061_ _10981_ _10982_ net1380 VGND VGND VPWR VPWR _02758_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_192_5099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22663_ rvcpu.dp.rf.reg_file_arr\[12\]\[18\] rvcpu.dp.rf.reg_file_arr\[13\]\[18\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[18\] rvcpu.dp.rf.reg_file_arr\[15\]\[18\] _09552_
+ _09721_ VGND VGND VPWR VPWR _09811_ sky130_fd_sc_hd__mux4_1
XFILLER_0_220_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_213_5615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24402_ _10380_ VGND VGND VPWR VPWR _02311_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21614_ _08864_ VGND VGND VPWR VPWR _01039_ sky130_fd_sc_hd__clkbuf_1
X_28170_ _12367_ net3078 _12546_ VGND VGND VPWR VPWR _12552_ sky130_fd_sc_hd__mux2_1
X_25382_ _10416_ _10936_ VGND VGND VPWR VPWR _10943_ sky130_fd_sc_hd__and2_1
X_22594_ _09743_ _09744_ _09421_ VGND VGND VPWR VPWR _09745_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27121_ _11956_ net1734 _11952_ _11959_ VGND VGND VPWR VPWR _03451_ sky130_fd_sc_hd__a31o_1
XFILLER_0_29_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24333_ _09248_ net4361 _10338_ VGND VGND VPWR VPWR _10343_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21545_ _08522_ VGND VGND VPWR VPWR _08798_ sky130_fd_sc_hd__buf_2
XFILLER_0_69_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_141_clk clknet_5_29__leaf_clk VGND VGND VPWR VPWR clknet_leaf_141_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_63_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27052_ _11904_ net1836 _11910_ _11916_ VGND VGND VPWR VPWR _03425_ sky130_fd_sc_hd__a31o_1
XFILLER_0_172_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24264_ _10304_ VGND VGND VPWR VPWR _02249_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_181_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21476_ rvcpu.dp.rf.reg_file_arr\[8\]\[5\] rvcpu.dp.rf.reg_file_arr\[10\]\[5\] rvcpu.dp.rf.reg_file_arr\[9\]\[5\]
+ rvcpu.dp.rf.reg_file_arr\[11\]\[5\] _08560_ _08561_ VGND VGND VPWR VPWR _08733_
+ sky130_fd_sc_hd__mux4_1
X_26003_ _09479_ _11315_ _11325_ _11326_ VGND VGND VPWR VPWR _02966_ sky130_fd_sc_hd__o211a_1
XFILLER_0_209_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20427_ datamem.data_ram\[6\]\[12\] _06629_ _07715_ _07718_ VGND VGND VPWR VPWR _07719_
+ sky130_fd_sc_hd__o211a_1
X_24195_ clknet_1_0__leaf__10079_ VGND VGND VPWR VPWR _10267_ sky130_fd_sc_hd__buf_1
XFILLER_0_160_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload190 clknet_leaf_224_clk VGND VGND VPWR VPWR clkload190/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_164_4423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20358_ datamem.data_ram\[8\]\[28\] _06696_ _06686_ datamem.data_ram\[12\]\[28\]
+ _07649_ VGND VGND VPWR VPWR _07650_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_164_4434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20289_ datamem.data_ram\[18\]\[19\] _06692_ _06635_ datamem.data_ram\[19\]\[19\]
+ _07031_ VGND VGND VPWR VPWR _07582_ sky130_fd_sc_hd__o221a_1
X_27954_ _12429_ VGND VGND VPWR VPWR _03814_ sky130_fd_sc_hd__clkbuf_1
X_23077_ _10100_ VGND VGND VPWR VPWR _01266_ sky130_fd_sc_hd__clkbuf_1
X_26905_ _11827_ _11823_ VGND VGND VPWR VPWR _11828_ sky130_fd_sc_hd__and2_1
X_22028_ _09252_ net3247 _09232_ VGND VGND VPWR VPWR _09253_ sky130_fd_sc_hd__mux2_1
X_27885_ _07203_ _10042_ _10918_ VGND VGND VPWR VPWR _12392_ sky130_fd_sc_hd__or3_1
Xhold30 rvcpu.dp.plde.PCPlus4E\[17\] VGND VGND VPWR VPWR net1180 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold41 rvcpu.dp.plem.PCPlus4M\[26\] VGND VGND VPWR VPWR net1191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2660 rvcpu.dp.rf.reg_file_arr\[18\]\[23\] VGND VGND VPWR VPWR net3810 sky130_fd_sc_hd__dlygate4sd3_1
X_14850_ _13287_ _13402_ VGND VGND VPWR VPWR _13403_ sky130_fd_sc_hd__nand2_4
XFILLER_0_199_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold52 rvcpu.dp.plem.lAuiPCM\[2\] VGND VGND VPWR VPWR net1202 sky130_fd_sc_hd__dlygate4sd3_1
X_29624_ net978 _01359_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[25\]\[27\] sky130_fd_sc_hd__dfxtp_1
Xhold2671 datamem.data_ram\[56\]\[15\] VGND VGND VPWR VPWR net3821 sky130_fd_sc_hd__dlygate4sd3_1
X_26836_ _11784_ VGND VGND VPWR VPWR _11785_ sky130_fd_sc_hd__clkbuf_2
Xhold63 rvcpu.dp.plde.PCPlus4E\[24\] VGND VGND VPWR VPWR net1213 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_67_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold74 rvcpu.dp.plde.PCPlus4E\[16\] VGND VGND VPWR VPWR net1224 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2682 datamem.data_ram\[24\]\[29\] VGND VGND VPWR VPWR net3832 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_67_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold85 rvcpu.dp.plem.lAuiPCM\[11\] VGND VGND VPWR VPWR net1235 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2693 datamem.data_ram\[38\]\[12\] VGND VGND VPWR VPWR net3843 sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 rvcpu.dp.plem.lAuiPCM\[15\] VGND VGND VPWR VPWR net1246 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_123_3441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_3452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1970 rvcpu.dp.rf.reg_file_arr\[2\]\[4\] VGND VGND VPWR VPWR net3120 sky130_fd_sc_hd__dlygate4sd3_1
X_26767_ _11735_ net1691 _11737_ _11743_ VGND VGND VPWR VPWR _03313_ sky130_fd_sc_hd__a31o_1
X_14781_ _13288_ _13286_ VGND VGND VPWR VPWR _13334_ sky130_fd_sc_hd__or2b_1
Xhold1981 rvcpu.dp.rf.reg_file_arr\[22\]\[6\] VGND VGND VPWR VPWR net3131 sky130_fd_sc_hd__dlygate4sd3_1
X_29555_ net909 _01290_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[27\]\[22\] sky130_fd_sc_hd__dfxtp_1
Xhold1992 datamem.data_ram\[20\]\[19\] VGND VGND VPWR VPWR net3142 sky130_fd_sc_hd__dlygate4sd3_1
X_23979_ clknet_1_1__leaf__10224_ VGND VGND VPWR VPWR _10239_ sky130_fd_sc_hd__buf_1
X_16520_ net3442 _14480_ _04489_ VGND VGND VPWR VPWR _04498_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_63_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28506_ _09275_ VGND VGND VPWR VPWR _12739_ sky130_fd_sc_hd__clkbuf_2
X_25718_ _11132_ VGND VGND VPWR VPWR _02875_ sky130_fd_sc_hd__clkbuf_1
X_26698_ _11700_ net1379 _11693_ _11703_ VGND VGND VPWR VPWR _03284_ sky130_fd_sc_hd__a31o_1
Xclkbuf_1_1__f__10267_ clknet_0__10267_ VGND VGND VPWR VPWR clknet_1_1__leaf__10267_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_58_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29486_ net848 _01221_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[2\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16451_ _04460_ VGND VGND VPWR VPWR _01815_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_196_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25649_ _10780_ _11094_ VGND VGND VPWR VPWR _11095_ sky130_fd_sc_hd__nor2_2
XFILLER_0_156_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28437_ _12698_ net2596 _12688_ VGND VGND VPWR VPWR _12699_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__10198_ clknet_0__10198_ VGND VGND VPWR VPWR clknet_1_1__leaf__10198_
+ sky130_fd_sc_hd__clkbuf_16
X_15402_ _13593_ _13764_ _13385_ _13360_ VGND VGND VPWR VPWR _13934_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_155_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19170_ _06482_ _06483_ VGND VGND VPWR VPWR _06484_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_26_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16382_ net2142 _14480_ _14547_ VGND VGND VPWR VPWR _14556_ sky130_fd_sc_hd__mux2_1
X_28368_ _12178_ _12602_ _12573_ VGND VGND VPWR VPWR _12659_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_213_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18121_ _05486_ _05487_ VGND VGND VPWR VPWR _05488_ sky130_fd_sc_hd__and2b_1
X_15333_ _13792_ _13864_ _13866_ _13869_ VGND VGND VPWR VPWR _13870_ sky130_fd_sc_hd__and4b_1
X_27319_ _12061_ net1482 _12065_ _12074_ VGND VGND VPWR VPWR _03534_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_97_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_132_clk clknet_5_30__leaf_clk VGND VGND VPWR VPWR clknet_leaf_132_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_22_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28299_ _08133_ _09268_ VGND VGND VPWR VPWR _12622_ sky130_fd_sc_hd__nor2_4
XFILLER_0_152_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18052_ rvcpu.dp.plem.ALUResultM\[8\] _05272_ _05267_ rvcpu.dp.plde.RD1E\[8\] _05420_
+ VGND VGND VPWR VPWR _05421_ sky130_fd_sc_hd__a221o_2
XFILLER_0_48_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30330_ net676 _02065_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[4\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15264_ _13355_ _13792_ _13795_ _13803_ VGND VGND VPWR VPWR _13804_ sky130_fd_sc_hd__or4b_1
XFILLER_0_152_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17003_ net1988 _14486_ _04719_ VGND VGND VPWR VPWR _04754_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_93_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_5 _02993_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_30261_ net615 _01996_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[6\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_15195_ _13282_ _13415_ VGND VGND VPWR VPWR _13737_ sky130_fd_sc_hd__or2_2
XFILLER_0_22_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32000_ clknet_leaf_134_clk _03422_ VGND VGND VPWR VPWR datamem.data_ram\[52\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30192_ net546 _01927_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[8\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18954_ _05549_ _06278_ VGND VGND VPWR VPWR _06291_ sky130_fd_sc_hd__and2_1
XFILLER_0_219_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_197_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17905_ _05277_ VGND VGND VPWR VPWR _05278_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_52_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18885_ _05467_ _05624_ _06212_ VGND VGND VPWR VPWR _06227_ sky130_fd_sc_hd__nand3_1
Xclkbuf_leaf_199_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_199_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_158_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32902_ clknet_leaf_214_clk _04324_ VGND VGND VPWR VPWR datamem.data_ram\[0\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_17836_ _05218_ VGND VGND VPWR VPWR rvcpu.dp.SrcBFW_Mux.y\[21\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_94_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_222_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_179_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32833_ clknet_leaf_254_clk _04255_ VGND VGND VPWR VPWR datamem.data_ram\[12\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_17767_ rvcpu.dp.plde.Rs2E\[1\] VGND VGND VPWR VPWR _05165_ sky130_fd_sc_hd__inv_2
X_14979_ _13414_ _13526_ _13390_ _13483_ _13304_ VGND VGND VPWR VPWR _13527_ sky130_fd_sc_hd__a311o_1
X_23603__223 clknet_1_1__leaf__10178_ VGND VGND VPWR VPWR net349 sky130_fd_sc_hd__inv_2
X_19506_ _06689_ VGND VGND VPWR VPWR _06802_ sky130_fd_sc_hd__clkbuf_8
X_16718_ _04603_ VGND VGND VPWR VPWR _01683_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32764_ clknet_leaf_256_clk _04186_ VGND VGND VPWR VPWR datamem.data_ram\[15\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17698_ _05123_ VGND VGND VPWR VPWR _01191_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23145__820 clknet_1_1__leaf__10107_ VGND VGND VPWR VPWR net946 sky130_fd_sc_hd__inv_2
X_19437_ _06732_ VGND VGND VPWR VPWR _06733_ sky130_fd_sc_hd__buf_8
X_31715_ net164 _03173_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[9\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16649_ _14181_ net3766 _04562_ VGND VGND VPWR VPWR _04567_ sky130_fd_sc_hd__mux2_1
XFILLER_0_190_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32695_ clknet_leaf_284_clk _04117_ VGND VGND VPWR VPWR datamem.data_ram\[18\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31646_ clknet_leaf_26_clk net1190 VGND VGND VPWR VPWR rvcpu.dp.plmw.lAuiPCW\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19368_ _06663_ VGND VGND VPWR VPWR _06664_ sky130_fd_sc_hd__buf_8
XFILLER_0_18_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18319_ _05683_ VGND VGND VPWR VPWR _05684_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_123_clk clknet_5_27__leaf_clk VGND VGND VPWR VPWR clknet_leaf_123_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_127_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_210_1292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31577_ clknet_leaf_74_clk datamem.rd_data_mem\[27\] VGND VGND VPWR VPWR rvcpu.dp.plmw.ReadDataW\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_19299_ _06592_ _06594_ VGND VGND VPWR VPWR _06595_ sky130_fd_sc_hd__nor2_4
XFILLER_0_5_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21330_ rvcpu.dp.plfd.InstrD\[20\] VGND VGND VPWR VPWR _08592_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_115_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30528_ clknet_leaf_268_clk _02263_ VGND VGND VPWR VPWR datamem.data_ram\[56\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold500 rvcpu.dp.plfd.PCPlus4D\[17\] VGND VGND VPWR VPWR net1650 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30459_ net137 _02194_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[19\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_21261_ _08522_ VGND VGND VPWR VPWR _08523_ sky130_fd_sc_hd__clkbuf_4
Xhold511 datamem.data_ram\[30\]\[3\] VGND VGND VPWR VPWR net1661 sky130_fd_sc_hd__dlygate4sd3_1
Xhold522 datamem.data_ram\[25\]\[0\] VGND VGND VPWR VPWR net1672 sky130_fd_sc_hd__dlygate4sd3_1
Xhold533 datamem.data_ram\[62\]\[5\] VGND VGND VPWR VPWR net1683 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20212_ _06797_ _07471_ _07482_ _07504_ VGND VGND VPWR VPWR _07505_ sky130_fd_sc_hd__a211oi_1
Xhold544 datamem.data_ram\[50\]\[6\] VGND VGND VPWR VPWR net1694 sky130_fd_sc_hd__dlygate4sd3_1
X_21192_ _08471_ _08476_ VGND VGND VPWR VPWR _08477_ sky130_fd_sc_hd__or2b_1
XFILLER_0_60_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold555 rvcpu.dp.plfd.InstrD\[11\] VGND VGND VPWR VPWR net1705 sky130_fd_sc_hd__dlygate4sd3_1
Xhold566 datamem.data_ram\[22\]\[5\] VGND VGND VPWR VPWR net1716 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_862 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold577 datamem.data_ram\[27\]\[1\] VGND VGND VPWR VPWR net1727 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_206_5430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold588 datamem.data_ram\[36\]\[1\] VGND VGND VPWR VPWR net1738 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_206_5441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20143_ datamem.data_ram\[42\]\[27\] _06611_ _07432_ _07435_ VGND VGND VPWR VPWR
+ _07436_ sky130_fd_sc_hd__o211a_1
X_32129_ clknet_leaf_229_clk _03551_ VGND VGND VPWR VPWR datamem.data_ram\[10\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold599 datamem.data_ram\[25\]\[1\] VGND VGND VPWR VPWR net1749 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24951_ _10694_ VGND VGND VPWR VPWR _02546_ sky130_fd_sc_hd__clkbuf_1
X_20074_ _07367_ VGND VGND VPWR VPWR _07368_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_202_5338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_202_5349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1200 rvcpu.dp.rf.reg_file_arr\[0\]\[25\] VGND VGND VPWR VPWR net2350 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_198_5242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23232__881 clknet_1_1__leaf__10125_ VGND VGND VPWR VPWR net1007 sky130_fd_sc_hd__inv_2
Xhold1211 datamem.data_ram\[15\]\[15\] VGND VGND VPWR VPWR net2361 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_198_5253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1222 datamem.data_ram\[38\]\[20\] VGND VGND VPWR VPWR net2372 sky130_fd_sc_hd__dlygate4sd3_1
X_27670_ _12083_ net2509 net51 VGND VGND VPWR VPWR _12272_ sky130_fd_sc_hd__mux2_1
X_24882_ _10657_ VGND VGND VPWR VPWR _02514_ sky130_fd_sc_hd__clkbuf_1
Xhold1233 datamem.data_ram\[17\]\[28\] VGND VGND VPWR VPWR net2383 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1244 datamem.data_ram\[56\]\[23\] VGND VGND VPWR VPWR net2394 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1255 rvcpu.dp.rf.reg_file_arr\[4\]\[12\] VGND VGND VPWR VPWR net2405 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1266 datamem.data_ram\[28\]\[22\] VGND VGND VPWR VPWR net2416 sky130_fd_sc_hd__dlygate4sd3_1
X_26621_ _11658_ VGND VGND VPWR VPWR _03252_ sky130_fd_sc_hd__clkbuf_1
X_23833_ _09310_ net3555 _10210_ VGND VGND VPWR VPWR _10213_ sky130_fd_sc_hd__mux2_1
Xhold1277 rvcpu.dp.rf.reg_file_arr\[5\]\[20\] VGND VGND VPWR VPWR net2427 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1288 rvcpu.dp.rf.reg_file_arr\[12\]\[30\] VGND VGND VPWR VPWR net2438 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__10221_ _10221_ VGND VGND VPWR VPWR clknet_0__10221_ sky130_fd_sc_hd__clkbuf_16
XANTENNA_406 _06643_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1299 rvcpu.dp.rf.reg_file_arr\[1\]\[4\] VGND VGND VPWR VPWR net2449 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_417 _06741_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29340_ clknet_leaf_173_clk _01075_ VGND VGND VPWR VPWR datamem.data_ram\[62\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_26552_ _10811_ net2862 _11620_ VGND VGND VPWR VPWR _11621_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_428 _06790_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_439 _06978_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20976_ datamem.data_ram\[44\]\[15\] datamem.data_ram\[45\]\[15\] _06933_ VGND VGND
+ VPWR VPWR _08265_ sky130_fd_sc_hd__mux2_1
X_23578__200 clknet_1_0__leaf__10176_ VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__inv_2
XFILLER_0_215_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__10152_ _10152_ VGND VGND VPWR VPWR clknet_0__10152_ sky130_fd_sc_hd__clkbuf_16
X_25503_ _11006_ VGND VGND VPWR VPWR _02786_ sky130_fd_sc_hd__clkbuf_1
X_22715_ rvcpu.dp.rf.reg_file_arr\[8\]\[21\] rvcpu.dp.rf.reg_file_arr\[10\]\[21\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[21\] rvcpu.dp.rf.reg_file_arr\[11\]\[21\] _09418_
+ _09485_ VGND VGND VPWR VPWR _09860_ sky130_fd_sc_hd__mux4_1
XFILLER_0_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29271_ _13156_ VGND VGND VPWR VPWR _04404_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_157_4260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_4271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28222_ _12367_ net3832 net45 VGND VGND VPWR VPWR _12580_ sky130_fd_sc_hd__mux2_1
X_25434_ _10973_ VGND VGND VPWR VPWR _02750_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__10083_ _10083_ VGND VGND VPWR VPWR clknet_0__10083_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_36_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22646_ _09437_ VGND VGND VPWR VPWR _09795_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_153_4157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_153_4168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_4179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28153_ _12458_ net3034 net73 VGND VGND VPWR VPWR _12543_ sky130_fd_sc_hd__mux2_1
X_25365_ _10876_ net1464 _10920_ _10931_ VGND VGND VPWR VPWR _02723_ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_114_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_114_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_146_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22577_ rvcpu.dp.rf.reg_file_arr\[28\]\[14\] rvcpu.dp.rf.reg_file_arr\[30\]\[14\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[14\] rvcpu.dp.rf.reg_file_arr\[31\]\[14\] _09443_
+ _09453_ VGND VGND VPWR VPWR _09729_ sky130_fd_sc_hd__mux4_1
XFILLER_0_8_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27104_ _11835_ _11941_ VGND VGND VPWR VPWR _11949_ sky130_fd_sc_hd__and2_1
X_24316_ _10333_ VGND VGND VPWR VPWR _02272_ sky130_fd_sc_hd__clkbuf_1
X_28084_ _12506_ VGND VGND VPWR VPWR _03867_ sky130_fd_sc_hd__clkbuf_1
X_21528_ _08725_ _08781_ VGND VGND VPWR VPWR _08782_ sky130_fd_sc_hd__nor2_1
X_25296_ _10758_ net2473 _10887_ VGND VGND VPWR VPWR _10891_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27035_ _11904_ net1662 _11897_ _11906_ VGND VGND VPWR VPWR _03418_ sky130_fd_sc_hd__a31o_1
XFILLER_0_107_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24247_ _09288_ net4077 _10288_ VGND VGND VPWR VPWR _10295_ sky130_fd_sc_hd__mux2_1
X_21459_ rvcpu.dp.rf.reg_file_arr\[12\]\[4\] rvcpu.dp.rf.reg_file_arr\[13\]\[4\] rvcpu.dp.rf.reg_file_arr\[14\]\[4\]
+ rvcpu.dp.rf.reg_file_arr\[15\]\[4\] _08567_ _08570_ VGND VGND VPWR VPWR _08717_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_121_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_3175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput20 net20 VGND VGND VPWR VPWR Instr[26] sky130_fd_sc_hd__buf_2
Xoutput7 net7 VGND VGND VPWR VPWR Instr[14] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_187_4990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput31 net31 VGND VGND VPWR VPWR Instr[7] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_183_4876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28986_ _13002_ VGND VGND VPWR VPWR _04273_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_183_4887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_4898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27937_ _12420_ VGND VGND VPWR VPWR _03806_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_125_3503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15951_ _14312_ VGND VGND VPWR VPWR _02051_ sky130_fd_sc_hd__clkbuf_1
Xhold3180 rvcpu.dp.rf.reg_file_arr\[24\]\[25\] VGND VGND VPWR VPWR net4330 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14902_ _13378_ _13398_ _13452_ VGND VGND VPWR VPWR _13453_ sky130_fd_sc_hd__o21ai_1
Xhold3191 rvcpu.dp.rf.reg_file_arr\[22\]\[15\] VGND VGND VPWR VPWR net4341 sky130_fd_sc_hd__dlygate4sd3_1
X_18670_ _05441_ _05421_ _05342_ _05349_ _05664_ _05669_ VGND VGND VPWR VPWR _06025_
+ sky130_fd_sc_hd__mux4_2
X_15882_ net3460 _13173_ _14275_ VGND VGND VPWR VPWR _14276_ sky130_fd_sc_hd__mux2_1
X_27868_ _12142_ net3877 net77 VGND VGND VPWR VPWR _12383_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2490 datamem.data_ram\[51\]\[29\] VGND VGND VPWR VPWR net3640 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29607_ net961 _01342_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[25\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_17621_ net2312 _13172_ _05082_ VGND VGND VPWR VPWR _05083_ sky130_fd_sc_hd__mux2_1
X_26819_ _11767_ net1635 _11773_ _11775_ VGND VGND VPWR VPWR _03333_ sky130_fd_sc_hd__a31o_1
X_14833_ _13376_ _13384_ _13385_ VGND VGND VPWR VPWR _13386_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_4_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27799_ _12341_ VGND VGND VPWR VPWR _03747_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_1078 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_204_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_142_3894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14764_ rvcpu.dp.pcreg.q\[6\] rvcpu.dp.pcreg.q\[5\] VGND VGND VPWR VPWR _13317_ sky130_fd_sc_hd__nor2_2
X_29538_ net892 _01273_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[27\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_17552_ _05045_ VGND VGND VPWR VPWR _05046_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_153_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16503_ _04466_ VGND VGND VPWR VPWR _04489_ sky130_fd_sc_hd__buf_4
XFILLER_0_156_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17483_ _14197_ _04900_ VGND VGND VPWR VPWR _05009_ sky130_fd_sc_hd__nand2_2
X_14695_ rvcpu.dp.plmw.ALUResultW\[7\] rvcpu.dp.plmw.ReadDataW\[7\] rvcpu.dp.plmw.PCPlus4W\[7\]
+ rvcpu.dp.plmw.lAuiPCW\[7\] _13192_ _13193_ VGND VGND VPWR VPWR _13256_ sky130_fd_sc_hd__mux4_2
X_29469_ net831 _01204_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[2\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_195_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19222_ _06527_ _06528_ VGND VGND VPWR VPWR _06529_ sky130_fd_sc_hd__nand2_1
X_31500_ clknet_leaf_26_clk rvcpu.dp.lAuiPCE\[26\] VGND VGND VPWR VPWR rvcpu.dp.plem.lAuiPCM\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_15_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16434_ net1905 _14463_ _04451_ VGND VGND VPWR VPWR _04452_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32480_ clknet_leaf_271_clk _03902_ VGND VGND VPWR VPWR datamem.data_ram\[26\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_15_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_4_Left_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31431_ clknet_leaf_53_clk _03134_ VGND VGND VPWR VPWR datamem.data_ram\[14\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_19153_ _06468_ rvcpu.dp.plde.ImmExtE\[17\] _06419_ VGND VGND VPWR VPWR _06469_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16365_ _14524_ VGND VGND VPWR VPWR _14547_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_105_clk clknet_5_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_105_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_183_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23060__759 clknet_1_0__leaf__10091_ VGND VGND VPWR VPWR net885 sky130_fd_sc_hd__inv_2
XFILLER_0_137_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15316_ _13494_ _13780_ VGND VGND VPWR VPWR _13853_ sky130_fd_sc_hd__nor2_1
XFILLER_0_171_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18104_ _05469_ _05470_ VGND VGND VPWR VPWR _05472_ sky130_fd_sc_hd__and2_1
XFILLER_0_171_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31362_ clknet_leaf_19_clk _03065_ VGND VGND VPWR VPWR rvcpu.dp.plde.ImmExtE\[11\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_41_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_17__f_clk clknet_2_2_0_clk VGND VGND VPWR VPWR clknet_5_17__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_42_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19084_ _06406_ _06407_ VGND VGND VPWR VPWR _06408_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16296_ _14510_ VGND VGND VPWR VPWR _01888_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_1342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30313_ net659 _02048_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[5\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15247_ _13785_ _13773_ _13786_ _13458_ VGND VGND VPWR VPWR _13787_ sky130_fd_sc_hd__a31o_1
X_18035_ _05356_ _05361_ _05404_ _05354_ VGND VGND VPWR VPWR _05405_ sky130_fd_sc_hd__a31o_1
XFILLER_0_2_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31293_ clknet_leaf_22_clk _02996_ VGND VGND VPWR VPWR rvcpu.dp.plde.JumpE sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23175__846 clknet_1_0__leaf__10111_ VGND VGND VPWR VPWR net972 sky130_fd_sc_hd__inv_2
XFILLER_0_140_968 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30244_ net598 _01979_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[7\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_15178_ _13397_ _13341_ VGND VGND VPWR VPWR _13721_ sky130_fd_sc_hd__nor2_2
X_30175_ clknet_leaf_197_clk _01910_ VGND VGND VPWR VPWR datamem.data_ram\[58\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19986_ datamem.data_ram\[14\]\[2\] _06950_ _06919_ datamem.data_ram\[13\]\[2\] _07279_
+ VGND VGND VPWR VPWR _07280_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18937_ _06269_ _06275_ VGND VGND VPWR VPWR _06276_ sky130_fd_sc_hd__or2_1
X_18868_ _05473_ _06210_ VGND VGND VPWR VPWR _06211_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_207_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_61 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17819_ _13197_ rvcpu.dp.plde.RD2E\[26\] _05196_ VGND VGND VPWR VPWR _05207_ sky130_fd_sc_hd__mux2_1
X_18799_ _05513_ _05727_ _06146_ VGND VGND VPWR VPWR _06147_ sky130_fd_sc_hd__a21o_1
XFILLER_0_222_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20830_ _08116_ _08118_ _08119_ VGND VGND VPWR VPWR _08120_ sky130_fd_sc_hd__and3_1
X_32816_ clknet_leaf_282_clk _04238_ VGND VGND VPWR VPWR datamem.data_ram\[13\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20761_ datamem.data_ram\[0\]\[6\] _07122_ _08048_ _07868_ _08050_ VGND VGND VPWR
+ VPWR _08051_ sky130_fd_sc_hd__a221o_1
X_32747_ clknet_leaf_212_clk _04169_ VGND VGND VPWR VPWR datamem.data_ram\[15\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22500_ _09385_ VGND VGND VPWR VPWR _09656_ sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_59_Left_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_174_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20692_ datamem.data_ram\[59\]\[5\] _06961_ _06926_ datamem.data_ram\[63\]\[5\] _06679_
+ VGND VGND VPWR VPWR _07983_ sky130_fd_sc_hd__a221o_1
X_32678_ clknet_leaf_245_clk _04100_ VGND VGND VPWR VPWR datamem.data_ram\[18\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24013__545 clknet_1_1__leaf__10242_ VGND VGND VPWR VPWR net671 sky130_fd_sc_hd__inv_2
XFILLER_0_147_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22431_ rvcpu.dp.rf.reg_file_arr\[12\]\[6\] rvcpu.dp.rf.reg_file_arr\[13\]\[6\] rvcpu.dp.rf.reg_file_arr\[14\]\[6\]
+ rvcpu.dp.rf.reg_file_arr\[15\]\[6\] _09552_ _09382_ VGND VGND VPWR VPWR _09591_
+ sky130_fd_sc_hd__mux4_1
X_31629_ clknet_leaf_65_clk net1214 VGND VGND VPWR VPWR rvcpu.dp.plmw.lAuiPCW\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23493__139 clknet_1_0__leaf__10160_ VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__inv_2
XFILLER_0_134_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25150_ _10807_ VGND VGND VPWR VPWR _02632_ sky130_fd_sc_hd__clkbuf_1
X_22362_ _08589_ VGND VGND VPWR VPWR _09525_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_150_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21313_ rvcpu.dp.plfd.InstrD\[19\] _08512_ VGND VGND VPWR VPWR _08575_ sky130_fd_sc_hd__nor2_4
XFILLER_0_103_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25081_ _10731_ net3288 net89 VGND VGND VPWR VPWR _10772_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22293_ _09422_ _09456_ _09457_ VGND VGND VPWR VPWR _09458_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_103_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold330 datamem.data_ram\[39\]\[3\] VGND VGND VPWR VPWR net1480 sky130_fd_sc_hd__dlygate4sd3_1
X_21244_ datamem.data_ram\[52\]\[25\] _08505_ datamem.data_ram\[53\]\[9\] _08506_
+ VGND VGND VPWR VPWR _08507_ sky130_fd_sc_hd__or4b_1
Xhold341 datamem.data_ram\[49\]\[0\] VGND VGND VPWR VPWR net1491 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold352 datamem.data_ram\[38\]\[2\] VGND VGND VPWR VPWR net1502 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold363 datamem.data_ram\[4\]\[1\] VGND VGND VPWR VPWR net1513 sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 datamem.data_ram\[14\]\[4\] VGND VGND VPWR VPWR net1524 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_68_Left_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28840_ _09225_ _11020_ _12886_ VGND VGND VPWR VPWR _12923_ sky130_fd_sc_hd__a21oi_2
Xhold385 datamem.data_ram\[48\]\[6\] VGND VGND VPWR VPWR net1535 sky130_fd_sc_hd__dlygate4sd3_1
X_21175_ _07903_ _08422_ _08436_ _08463_ VGND VGND VPWR VPWR _08464_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_229_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold396 datamem.data_ram\[37\]\[0\] VGND VGND VPWR VPWR net1546 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_225_5894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20126_ datamem.data_ram\[7\]\[27\] _06671_ _06657_ datamem.data_ram\[1\]\[27\] VGND
+ VGND VPWR VPWR _07419_ sky130_fd_sc_hd__o22a_1
X_25983_ _11143_ VGND VGND VPWR VPWR _11315_ sky130_fd_sc_hd__buf_2
X_28771_ _06591_ VGND VGND VPWR VPWR _12886_ sky130_fd_sc_hd__buf_8
X_24934_ _10685_ VGND VGND VPWR VPWR _02538_ sky130_fd_sc_hd__clkbuf_1
X_27722_ _12083_ net3631 net49 VGND VGND VPWR VPWR _12300_ sky130_fd_sc_hd__mux2_1
X_20057_ datamem.data_ram\[45\]\[26\] _06660_ _06644_ datamem.data_ram\[40\]\[26\]
+ VGND VGND VPWR VPWR _07351_ sky130_fd_sc_hd__o22a_1
Xhold1030 datamem.data_ram\[62\]\[14\] VGND VGND VPWR VPWR net2180 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1041 rvcpu.dp.rf.reg_file_arr\[1\]\[12\] VGND VGND VPWR VPWR net2191 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1052 rvcpu.dp.rf.reg_file_arr\[10\]\[18\] VGND VGND VPWR VPWR net2202 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_159_4300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24865_ _10648_ VGND VGND VPWR VPWR _02506_ sky130_fd_sc_hd__clkbuf_1
Xhold1063 rvcpu.dp.rf.reg_file_arr\[17\]\[31\] VGND VGND VPWR VPWR net2213 sky130_fd_sc_hd__dlygate4sd3_1
X_27653_ _12145_ net3373 net79 VGND VGND VPWR VPWR _12263_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_159_4311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1074 datamem.data_ram\[19\]\[14\] VGND VGND VPWR VPWR net2224 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_159_4322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1085 rvcpu.dp.rf.reg_file_arr\[0\]\[3\] VGND VGND VPWR VPWR net2235 sky130_fd_sc_hd__dlygate4sd3_1
X_26604_ _11618_ net1798 _11639_ _11649_ VGND VGND VPWR VPWR _03244_ sky130_fd_sc_hd__a31o_1
XANTENNA_203 _09482_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1096 rvcpu.dp.rf.reg_file_arr\[9\]\[18\] VGND VGND VPWR VPWR net2246 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_213_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27584_ _12128_ net2407 _12224_ VGND VGND VPWR VPWR _12226_ sky130_fd_sc_hd__mux2_1
XANTENNA_214 _09750_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_217_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_225 _10060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24796_ _10610_ VGND VGND VPWR VPWR _02475_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_236 _10268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_155_4208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__10204_ _10204_ VGND VGND VPWR VPWR clknet_0__10204_ sky130_fd_sc_hd__clkbuf_16
X_26535_ _11517_ net1670 _11608_ _11611_ VGND VGND VPWR VPWR _03213_ sky130_fd_sc_hd__a31o_1
XANTENNA_247 _11978_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_4219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29323_ clknet_leaf_12_clk _01058_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD1E\[30\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__10104_ clknet_0__10104_ VGND VGND VPWR VPWR clknet_1_1__leaf__10104_
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_258 _13201_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_269 _13229_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_81_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20959_ datamem.data_ram\[60\]\[15\] datamem.data_ram\[61\]\[15\] _06933_ VGND VGND
+ VPWR VPWR _08248_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__10135_ _10135_ VGND VGND VPWR VPWR clknet_0__10135_ sky130_fd_sc_hd__clkbuf_16
X_26484__38 clknet_1_0__leaf__10267_ VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__inv_2
X_26466_ _11535_ rvcpu.ALUResultE\[27\] _11288_ VGND VGND VPWR VPWR _11589_ sky130_fd_sc_hd__a21o_1
XFILLER_0_165_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29254_ _13147_ VGND VGND VPWR VPWR _04396_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23678_ clknet_1_0__leaf__10192_ VGND VGND VPWR VPWR _10194_ sky130_fd_sc_hd__buf_1
XFILLER_0_138_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25417_ _10964_ VGND VGND VPWR VPWR _02742_ sky130_fd_sc_hd__clkbuf_1
X_28205_ _12570_ VGND VGND VPWR VPWR _03924_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29185_ _09255_ net2339 net63 VGND VGND VPWR VPWR _13110_ sky130_fd_sc_hd__mux2_1
X_22629_ rvcpu.dp.rf.reg_file_arr\[16\]\[17\] rvcpu.dp.rf.reg_file_arr\[17\]\[17\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[17\] rvcpu.dp.rf.reg_file_arr\[19\]\[17\] _09512_
+ _09513_ VGND VGND VPWR VPWR _09778_ sky130_fd_sc_hd__mux4_2
X_26397_ _11524_ rvcpu.ALUResultE\[6\] _06392_ _11540_ VGND VGND VPWR VPWR _11541_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_192_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28136_ _12441_ net3194 _12528_ VGND VGND VPWR VPWR _12534_ sky130_fd_sc_hd__mux2_1
X_16150_ net2275 _13275_ _14384_ VGND VGND VPWR VPWR _14418_ sky130_fd_sc_hd__mux2_1
X_25348_ _08124_ _07903_ VGND VGND VPWR VPWR _10922_ sky130_fd_sc_hd__nor2_2
XFILLER_0_134_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_114_3226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_3237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15101_ _13314_ _13292_ VGND VGND VPWR VPWR _13646_ sky130_fd_sc_hd__and2_2
XFILLER_0_140_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28067_ _12497_ VGND VGND VPWR VPWR _03859_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_79_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16081_ _14381_ VGND VGND VPWR VPWR _01982_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25279_ _10731_ net4046 _10878_ VGND VGND VPWR VPWR _10882_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_185_4927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15032_ _13343_ _13578_ VGND VGND VPWR VPWR _13579_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_185_4938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27018_ _11889_ net1619 _11885_ _11895_ VGND VGND VPWR VPWR _03412_ sky130_fd_sc_hd__a31o_1
X_23239__887 clknet_1_1__leaf__10126_ VGND VGND VPWR VPWR net1013 sky130_fd_sc_hd__inv_2
XFILLER_0_107_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19840_ datamem.data_ram\[45\]\[1\] _07132_ _07133_ datamem.data_ram\[41\]\[1\] _07134_
+ VGND VGND VPWR VPWR _07135_ sky130_fd_sc_hd__a221o_1
XFILLER_0_43_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19771_ datamem.data_ram\[27\]\[25\] _06829_ _07024_ datamem.data_ram\[28\]\[25\]
+ _07065_ VGND VGND VPWR VPWR _07066_ sky130_fd_sc_hd__o221a_1
X_28969_ _10063_ _12989_ VGND VGND VPWR VPWR _12993_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_88_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16983_ net4267 _14466_ _04742_ VGND VGND VPWR VPWR _04744_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_88_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18722_ _05331_ _05974_ _06072_ _06073_ VGND VGND VPWR VPWR _06074_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_144_3945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15934_ net1902 _13260_ _14297_ VGND VGND VPWR VPWR _14303_ sky130_fd_sc_hd__mux2_1
X_31980_ clknet_leaf_138_clk _03402_ VGND VGND VPWR VPWR datamem.data_ram\[53\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_204_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30931_ clknet_leaf_156_clk _02666_ VGND VGND VPWR VPWR datamem.data_ram\[40\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_18653_ _05771_ _05862_ _05696_ VGND VGND VPWR VPWR _06009_ sky130_fd_sc_hd__a21o_1
X_15865_ net2208 _13263_ _14258_ VGND VGND VPWR VPWR _14265_ sky130_fd_sc_hd__mux2_1
XFILLER_0_203_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23975__511 clknet_1_1__leaf__10238_ VGND VGND VPWR VPWR net637 sky130_fd_sc_hd__inv_2
XFILLER_0_8_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17604_ _05073_ VGND VGND VPWR VPWR _01235_ sky130_fd_sc_hd__clkbuf_1
X_14816_ _13296_ _13281_ VGND VGND VPWR VPWR _13369_ sky130_fd_sc_hd__nand2_4
XFILLER_0_188_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18584_ _05709_ _05826_ VGND VGND VPWR VPWR _05943_ sky130_fd_sc_hd__and2_1
X_30862_ clknet_leaf_280_clk _02597_ VGND VGND VPWR VPWR datamem.data_ram\[43\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15796_ _14185_ net4016 _14221_ VGND VGND VPWR VPWR _14228_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32601_ clknet_leaf_244_clk _04023_ VGND VGND VPWR VPWR datamem.data_ram\[20\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_47_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17535_ _13257_ net2262 _05032_ VGND VGND VPWR VPWR _05037_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14747_ _13299_ VGND VGND VPWR VPWR _13300_ sky130_fd_sc_hd__buf_2
XFILLER_0_15_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30793_ clknet_leaf_264_clk _02528_ VGND VGND VPWR VPWR datamem.data_ram\[46\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_103_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32532_ clknet_leaf_245_clk _03954_ VGND VGND VPWR VPWR datamem.data_ram\[23\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14678_ rvcpu.dp.plmw.ALUResultW\[11\] rvcpu.dp.plmw.ReadDataW\[11\] rvcpu.dp.plmw.PCPlus4W\[11\]
+ rvcpu.dp.plmw.lAuiPCW\[11\] _13168_ _13170_ VGND VGND VPWR VPWR _13243_ sky130_fd_sc_hd__mux4_2
XFILLER_0_129_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17466_ _05000_ VGND VGND VPWR VPWR _01308_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19205_ rvcpu.dp.plde.ImmExtE\[24\] rvcpu.dp.plde.PCE\[24\] VGND VGND VPWR VPWR _06514_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16417_ net3306 _14447_ _14572_ VGND VGND VPWR VPWR _14575_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32463_ clknet_leaf_184_clk _03885_ VGND VGND VPWR VPWR datamem.data_ram\[26\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_17397_ _14179_ net3359 _04960_ VGND VGND VPWR VPWR _04964_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19136_ _06453_ rvcpu.dp.plde.ImmExtE\[15\] _06419_ VGND VGND VPWR VPWR _06454_ sky130_fd_sc_hd__mux2_1
X_31414_ clknet_leaf_23_clk _03117_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCE\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16348_ _14538_ VGND VGND VPWR VPWR _01864_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32394_ clknet_leaf_81_clk _03816_ VGND VGND VPWR VPWR datamem.data_ram\[29\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19067_ _06393_ VGND VGND VPWR VPWR rvcpu.dp.lAuiPCE\[6\] sky130_fd_sc_hd__clkbuf_1
X_31345_ clknet_leaf_19_clk _03048_ VGND VGND VPWR VPWR rvcpu.dp.plde.ALUControlE\[1\]
+ sky130_fd_sc_hd__dfxtp_2
X_16279_ net2428 _14445_ _14500_ VGND VGND VPWR VPWR _14502_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18018_ rvcpu.dp.plde.RD1E\[1\] _05265_ _05269_ _13274_ _05387_ VGND VGND VPWR VPWR
+ _05388_ sky130_fd_sc_hd__a221oi_4
XFILLER_0_2_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31276_ clknet_leaf_125_clk _02979_ VGND VGND VPWR VPWR datamem.data_ram\[24\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__10124_ clknet_0__10124_ VGND VGND VPWR VPWR clknet_1_0__leaf__10124_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30227_ net581 _01962_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[7\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_227_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30158_ net520 _01893_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[0\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_19969_ _06777_ _07255_ _07257_ _07262_ VGND VGND VPWR VPWR _07263_ sky130_fd_sc_hd__a31o_1
XFILLER_0_96_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_226_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30089_ net451 _01824_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[11\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_22971__679 clknet_1_0__leaf__10082_ VGND VGND VPWR VPWR net805 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_220_5780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21931_ rvcpu.dp.rf.reg_file_arr\[28\]\[29\] rvcpu.dp.rf.reg_file_arr\[30\]\[29\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[29\] rvcpu.dp.rf.reg_file_arr\[31\]\[29\] _08629_
+ _08683_ VGND VGND VPWR VPWR _09164_ sky130_fd_sc_hd__mux4_1
XFILLER_0_59_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_179_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24650_ _10400_ net2272 _10521_ VGND VGND VPWR VPWR _10529_ sky130_fd_sc_hd__mux2_1
X_21862_ _08795_ _09094_ _09096_ _09098_ VGND VGND VPWR VPWR _09099_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_210_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_118_Right_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20813_ datamem.data_ram\[63\]\[30\] _07860_ _07862_ datamem.data_ram\[61\]\[30\]
+ _08102_ VGND VGND VPWR VPWR _08103_ sky130_fd_sc_hd__o221a_1
X_24581_ _10142_ _10347_ _10366_ VGND VGND VPWR VPWR _10491_ sky130_fd_sc_hd__a21oi_4
X_21793_ _08682_ _09031_ _09033_ _08558_ VGND VGND VPWR VPWR _09034_ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23344__982 clknet_1_1__leaf__10136_ VGND VGND VPWR VPWR net1108 sky130_fd_sc_hd__inv_2
X_26320_ net1808 _11436_ VGND VGND VPWR VPWR _11493_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20744_ datamem.data_ram\[44\]\[6\] _06615_ _06642_ datamem.data_ram\[40\]\[6\] _08033_
+ VGND VGND VPWR VPWR _08034_ sky130_fd_sc_hd__a221o_1
X_23501__146 clknet_1_0__leaf__10161_ VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__inv_2
XFILLER_0_64_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_212_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_175_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26251_ _11438_ _11458_ _11459_ net1306 VGND VGND VPWR VPWR _03081_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_150_4105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_189_5027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20675_ datamem.data_ram\[46\]\[5\] _06978_ _06948_ datamem.data_ram\[41\]\[5\] VGND
+ VGND VPWR VPWR _07966_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_189_5038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25202_ _10811_ net3959 net56 VGND VGND VPWR VPWR _10840_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22414_ _09566_ _09570_ _09574_ _09491_ VGND VGND VPWR VPWR _01129_ sky130_fd_sc_hd__o31a_1
X_26182_ _08572_ _11413_ VGND VGND VPWR VPWR _11428_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23394_ _09318_ net3146 _10143_ VGND VGND VPWR VPWR _10148_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25133_ _10798_ VGND VGND VPWR VPWR _02624_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22345_ _09476_ _09506_ _09508_ _09489_ VGND VGND VPWR VPWR _09509_ sky130_fd_sc_hd__o211a_1
XFILLER_0_143_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_227_5934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_76_Left_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_227_5945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25064_ _10761_ VGND VGND VPWR VPWR _02592_ sky130_fd_sc_hd__clkbuf_1
X_29941_ net311 _01676_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[15\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22276_ _09413_ VGND VGND VPWR VPWR _09441_ sky130_fd_sc_hd__buf_2
XFILLER_0_14_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_4045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_148_4056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold160 datamem.data_ram\[44\]\[0\] VGND VGND VPWR VPWR net1310 sky130_fd_sc_hd__dlygate4sd3_1
X_21227_ _08468_ _08353_ _08489_ VGND VGND VPWR VPWR _04439_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_104_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold171 datamem.data_ram\[45\]\[3\] VGND VGND VPWR VPWR net1321 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29872_ net250 _01607_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[17\]\[3\] sky130_fd_sc_hd__dfxtp_1
Xhold182 datamem.data_ram\[41\]\[3\] VGND VGND VPWR VPWR net1332 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_180_4813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold193 datamem.data_ram\[45\]\[2\] VGND VGND VPWR VPWR net1343 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_180_4824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28823_ _09225_ _10960_ _12886_ VGND VGND VPWR VPWR _12914_ sky130_fd_sc_hd__a21oi_4
X_21158_ _08437_ _08438_ _08441_ _08446_ VGND VGND VPWR VPWR _08447_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_6_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_6_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20109_ datamem.data_ram\[19\]\[10\] _06812_ _06685_ datamem.data_ram\[20\]\[10\]
+ _06732_ VGND VGND VPWR VPWR _07403_ sky130_fd_sc_hd__o221a_1
X_28754_ _12601_ _10997_ _12795_ VGND VGND VPWR VPWR _12877_ sky130_fd_sc_hd__a21oi_4
X_21089_ datamem.data_ram\[48\]\[7\] _06935_ _06953_ datamem.data_ram\[52\]\[7\] _08377_
+ VGND VGND VPWR VPWR _08378_ sky130_fd_sc_hd__a221o_1
X_25966_ net29 _11289_ VGND VGND VPWR VPWR _11306_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_107_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27705_ _12145_ net4111 net50 VGND VGND VPWR VPWR _12291_ sky130_fd_sc_hd__mux2_1
X_24917_ _10676_ VGND VGND VPWR VPWR _02530_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_107_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25897_ _13823_ _11256_ _11258_ _11266_ VGND VGND VPWR VPWR _02920_ sky130_fd_sc_hd__o211a_1
X_28685_ _12840_ VGND VGND VPWR VPWR _04134_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_107_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_85_Left_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27636_ _12253_ VGND VGND VPWR VPWR _03672_ sky130_fd_sc_hd__clkbuf_1
X_15650_ _13189_ VGND VGND VPWR VPWR _14137_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_178_4764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24848_ _10454_ net2223 _10631_ VGND VGND VPWR VPWR _10639_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_4775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_217_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_198_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14601_ net2159 _13184_ _13181_ VGND VGND VPWR VPWR _13185_ sky130_fd_sc_hd__mux2_1
X_15581_ net2226 _13198_ _14092_ VGND VGND VPWR VPWR _14098_ sky130_fd_sc_hd__mux2_1
X_24779_ net108 _10600_ VGND VGND VPWR VPWR _10601_ sky130_fd_sc_hd__nor2_2
X_27567_ _12083_ net4113 net82 VGND VGND VPWR VPWR _12217_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_197_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29306_ clknet_leaf_0_clk _01041_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD1E\[13\] sky130_fd_sc_hd__dfxtp_1
X_17320_ net3512 _13240_ _04913_ VGND VGND VPWR VPWR _04923_ sky130_fd_sc_hd__mux2_1
X_26518_ _11603_ _10600_ VGND VGND VPWR VPWR _11604_ sky130_fd_sc_hd__nor2_4
XFILLER_0_51_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27498_ _12180_ VGND VGND VPWR VPWR _03607_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_172_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17251_ _14170_ net4324 _04876_ VGND VGND VPWR VPWR _04886_ sky130_fd_sc_hd__mux2_1
X_29237_ _13138_ VGND VGND VPWR VPWR _04388_ sky130_fd_sc_hd__clkbuf_1
X_26449_ _11576_ _11210_ _11540_ _06499_ _11577_ VGND VGND VPWR VPWR _11578_ sky130_fd_sc_hd__a221o_1
XFILLER_0_113_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_3782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16202_ _13228_ VGND VGND VPWR VPWR _14453_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_137_3793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17182_ _04849_ VGND VGND VPWR VPWR _01449_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_226_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29168_ _09255_ net3769 net64 VGND VGND VPWR VPWR _13101_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23556__180 clknet_1_1__leaf__10174_ VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_77_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16133_ _14409_ VGND VGND VPWR VPWR _01958_ sky130_fd_sc_hd__clkbuf_1
X_28119_ _12367_ net4100 net74 VGND VGND VPWR VPWR _12525_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_94_Left_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_133_3679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29099_ _13064_ VGND VGND VPWR VPWR _04324_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31130_ clknet_leaf_125_clk _02865_ VGND VGND VPWR VPWR datamem.data_ram\[25\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_16064_ net3932 _13248_ _14371_ VGND VGND VPWR VPWR _14373_ sky130_fd_sc_hd__mux2_1
X_15015_ _13559_ _13561_ _13562_ VGND VGND VPWR VPWR _13563_ sky130_fd_sc_hd__a21oi_1
X_31061_ clknet_leaf_255_clk _02796_ VGND VGND VPWR VPWR datamem.data_ram\[8\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_30012_ clknet_leaf_175_clk _01747_ VGND VGND VPWR VPWR datamem.data_ram\[59\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19823_ _06596_ _07106_ _07117_ _06797_ VGND VGND VPWR VPWR _07118_ sky130_fd_sc_hd__a22o_1
XFILLER_0_166_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24042__571 clknet_1_1__leaf__10245_ VGND VGND VPWR VPWR net697 sky130_fd_sc_hd__inv_2
XFILLER_0_120_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19754_ datamem.data_ram\[59\]\[25\] _06812_ _06765_ datamem.data_ram\[60\]\[25\]
+ VGND VGND VPWR VPWR _07049_ sky130_fd_sc_hd__o22a_1
XFILLER_0_21_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16966_ net2491 _14449_ _04731_ VGND VGND VPWR VPWR _04735_ sky130_fd_sc_hd__mux2_1
XFILLER_0_223_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18705_ _05673_ _05680_ _05677_ VGND VGND VPWR VPWR _06058_ sky130_fd_sc_hd__mux2_1
X_15917_ net2195 _13235_ _14286_ VGND VGND VPWR VPWR _14294_ sky130_fd_sc_hd__mux2_1
XFILLER_0_223_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19685_ datamem.data_ram\[58\]\[0\] _06931_ _06942_ datamem.data_ram\[59\]\[0\] _06769_
+ VGND VGND VPWR VPWR _06981_ sky130_fd_sc_hd__a221o_1
X_31963_ clknet_leaf_122_clk _03385_ VGND VGND VPWR VPWR datamem.data_ram\[28\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_16897_ _04698_ VGND VGND VPWR VPWR _01591_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18636_ _05594_ _05956_ _05346_ VGND VGND VPWR VPWR _05993_ sky130_fd_sc_hd__a21oi_1
X_30914_ clknet_leaf_181_clk _02649_ VGND VGND VPWR VPWR datamem.data_ram\[41\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_15848_ net2067 _13238_ _14247_ VGND VGND VPWR VPWR _14256_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31894_ clknet_leaf_113_clk _03348_ VGND VGND VPWR VPWR datamem.data_ram\[36\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_188_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18567_ _05692_ _05926_ VGND VGND VPWR VPWR _05927_ sky130_fd_sc_hd__nor2_1
X_30845_ clknet_leaf_220_clk _02580_ VGND VGND VPWR VPWR datamem.data_ram\[43\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_15779_ _14168_ net3301 _14210_ VGND VGND VPWR VPWR _14219_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17518_ _13232_ net3849 _05021_ VGND VGND VPWR VPWR _05028_ sky130_fd_sc_hd__mux2_1
X_18498_ _05383_ _05397_ VGND VGND VPWR VPWR _05860_ sky130_fd_sc_hd__nand2_1
X_30776_ clknet_leaf_220_clk _02511_ VGND VGND VPWR VPWR datamem.data_ram\[46\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32515_ clknet_leaf_77_clk _03937_ VGND VGND VPWR VPWR datamem.data_ram\[24\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_17449_ _04991_ VGND VGND VPWR VPWR _01316_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_1223 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32446_ clknet_leaf_82_clk _03868_ VGND VGND VPWR VPWR datamem.data_ram\[27\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_20460_ datamem.data_ram\[31\]\[20\] _06707_ _07748_ _07751_ VGND VGND VPWR VPWR
+ _07752_ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19119_ _06438_ rvcpu.dp.plde.ImmExtE\[13\] _06419_ VGND VGND VPWR VPWR _06439_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32377_ clknet_leaf_160_clk _03799_ VGND VGND VPWR VPWR datamem.data_ram\[2\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_20391_ datamem.data_ram\[18\]\[28\] _06728_ _06766_ datamem.data_ram\[20\]\[28\]
+ _07682_ VGND VGND VPWR VPWR _07683_ sky130_fd_sc_hd__o221a_1
XFILLER_0_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22130_ _09334_ VGND VGND VPWR VPWR _01085_ sky130_fd_sc_hd__clkbuf_1
X_31328_ clknet_leaf_24_clk _03031_ VGND VGND VPWR VPWR rvcpu.dp.plde.funct3E\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_28_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22061_ _09279_ net3475 _09270_ VGND VGND VPWR VPWR _09280_ sky130_fd_sc_hd__mux2_1
X_31259_ clknet_leaf_15_clk _02962_ VGND VGND VPWR VPWR rvcpu.dp.plfd.InstrD\[17\]
+ sky130_fd_sc_hd__dfxtp_4
Xclkbuf_1_0__f__10107_ clknet_0__10107_ VGND VGND VPWR VPWR clknet_1_0__leaf__10107_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_222_5820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21012_ _07859_ _08300_ VGND VGND VPWR VPWR _08301_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_222_5831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23442__93 clknet_1_0__leaf__10155_ VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__inv_2
X_25820_ _08621_ VGND VGND VPWR VPWR _11207_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_226_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_215_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25751_ _08598_ VGND VGND VPWR VPWR _11155_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_94_clk clknet_5_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_94_clk sky130_fd_sc_hd__clkbuf_8
X_24702_ _10558_ VGND VGND VPWR VPWR _02433_ sky130_fd_sc_hd__clkbuf_1
X_21914_ _08673_ _09147_ VGND VGND VPWR VPWR _09148_ sky130_fd_sc_hd__or2_1
X_25682_ _07131_ _07177_ VGND VGND VPWR VPWR _11112_ sky130_fd_sc_hd__nor2_1
XFILLER_0_168_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28470_ _12717_ VGND VGND VPWR VPWR _04042_ sky130_fd_sc_hd__clkbuf_1
X_22894_ rvcpu.dp.plfd.InstrD\[22\] _10028_ VGND VGND VPWR VPWR _10029_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24633_ _10519_ VGND VGND VPWR VPWR _02403_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27421_ _12132_ net2788 _12126_ VGND VGND VPWR VPWR _12133_ sky130_fd_sc_hd__mux2_1
X_24019__551 clknet_1_0__leaf__10242_ VGND VGND VPWR VPWR net677 sky130_fd_sc_hd__inv_2
X_21845_ _08510_ _09082_ VGND VGND VPWR VPWR _09083_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_179_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_216_5668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24564_ _10142_ _10337_ _10366_ VGND VGND VPWR VPWR _10482_ sky130_fd_sc_hd__a21oi_4
X_27352_ _09325_ VGND VGND VPWR VPWR _12093_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_216_5679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_4650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21776_ rvcpu.dp.rf.reg_file_arr\[12\]\[20\] rvcpu.dp.rf.reg_file_arr\[13\]\[20\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[20\] rvcpu.dp.rf.reg_file_arr\[15\]\[20\] _08696_
+ _08553_ VGND VGND VPWR VPWR _09018_ sky130_fd_sc_hd__mux4_1
XFILLER_0_110_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_194_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26303_ _11484_ VGND VGND VPWR VPWR _03108_ sky130_fd_sc_hd__clkbuf_1
X_23515_ _09244_ net4096 _10162_ VGND VGND VPWR VPWR _10166_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20727_ datamem.data_ram\[21\]\[6\] _07132_ _07123_ datamem.data_ram\[20\]\[6\] _08016_
+ VGND VGND VPWR VPWR _08017_ sky130_fd_sc_hd__a221o_1
X_27283_ _10325_ _11054_ _11898_ VGND VGND VPWR VPWR _12054_ sky130_fd_sc_hd__and3_1
XFILLER_0_167_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24495_ _09330_ datamem.data_ram\[52\]\[31\] _10430_ VGND VGND VPWR VPWR _10438_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26234_ _11379_ _03030_ _11454_ VGND VGND VPWR VPWR _03067_ sky130_fd_sc_hd__a21o_1
X_29022_ _12739_ net2615 net66 VGND VGND VPWR VPWR _13023_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20658_ datamem.data_ram\[43\]\[29\] _06828_ _06789_ datamem.data_ram\[41\]\[29\]
+ _06851_ VGND VGND VPWR VPWR _07949_ sky130_fd_sc_hd__o221a_1
XFILLER_0_163_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26165_ _11419_ VGND VGND VPWR VPWR _03035_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20589_ datamem.data_ram\[16\]\[13\] datamem.data_ram\[17\]\[13\] _07826_ VGND VGND
+ VPWR VPWR _07880_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25116_ _10789_ VGND VGND VPWR VPWR _02616_ sky130_fd_sc_hd__clkbuf_1
X_22328_ rvcpu.dp.rf.reg_file_arr\[16\]\[2\] rvcpu.dp.rf.reg_file_arr\[17\]\[2\] rvcpu.dp.rf.reg_file_arr\[18\]\[2\]
+ rvcpu.dp.rf.reg_file_arr\[19\]\[2\] _09416_ _09443_ VGND VGND VPWR VPWR _09492_
+ sky130_fd_sc_hd__mux4_1
X_26096_ net1594 _11372_ VGND VGND VPWR VPWR _11383_ sky130_fd_sc_hd__and2_1
XFILLER_0_103_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_72_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29924_ net294 _01659_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[16\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_25047_ _10480_ net2184 net90 VGND VGND VPWR VPWR _10750_ sky130_fd_sc_hd__mux2_1
X_22259_ rvcpu.dp.rf.reg_file_arr\[4\]\[0\] rvcpu.dp.rf.reg_file_arr\[5\]\[0\] rvcpu.dp.rf.reg_file_arr\[6\]\[0\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[0\] _09423_ _09424_ VGND VGND VPWR VPWR _09425_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_167_4498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29855_ net233 _01590_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[18\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16820_ _04657_ VGND VGND VPWR VPWR _01627_ sky130_fd_sc_hd__clkbuf_1
X_28806_ _09225_ _10997_ _12886_ VGND VGND VPWR VPWR _12905_ sky130_fd_sc_hd__a21oi_4
X_29786_ net1132 _01521_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[20\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26998_ _11883_ VGND VGND VPWR VPWR _03404_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_217_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16751_ net2624 _14438_ _04612_ VGND VGND VPWR VPWR _04621_ sky130_fd_sc_hd__mux2_1
X_28737_ _10979_ _12622_ _12795_ VGND VGND VPWR VPWR _12868_ sky130_fd_sc_hd__a21oi_1
X_25949_ net1860 _11290_ _11286_ _11296_ VGND VGND VPWR VPWR _02942_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_85_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_85_clk sky130_fd_sc_hd__clkbuf_8
X_15702_ _13243_ VGND VGND VPWR VPWR _14172_ sky130_fd_sc_hd__buf_4
X_19470_ _06765_ VGND VGND VPWR VPWR _06766_ sky130_fd_sc_hd__buf_6
X_16682_ _04584_ VGND VGND VPWR VPWR _01700_ sky130_fd_sc_hd__clkbuf_1
X_28668_ _12831_ VGND VGND VPWR VPWR _04126_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18421_ _05784_ VGND VGND VPWR VPWR _05785_ sky130_fd_sc_hd__buf_2
XFILLER_0_213_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27619_ _12244_ VGND VGND VPWR VPWR _03664_ sky130_fd_sc_hd__clkbuf_1
X_15633_ net1918 _13275_ _14091_ VGND VGND VPWR VPWR _14125_ sky130_fd_sc_hd__mux2_1
XFILLER_0_185_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28599_ _12794_ VGND VGND VPWR VPWR _04094_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_3822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_201_577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_3833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18352_ _05707_ _05712_ _05716_ VGND VGND VPWR VPWR _05717_ sky130_fd_sc_hd__a21o_1
X_30630_ clknet_leaf_217_clk _02365_ VGND VGND VPWR VPWR datamem.data_ram\[51\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_15564_ _14075_ _14076_ _14078_ _14087_ VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__a31oi_2
XFILLER_0_115_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_185_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17303_ _04914_ VGND VGND VPWR VPWR _01393_ sky130_fd_sc_hd__clkbuf_1
X_15495_ _13337_ _13474_ _13995_ _13475_ VGND VGND VPWR VPWR _14023_ sky130_fd_sc_hd__o211a_1
X_18283_ _05286_ VGND VGND VPWR VPWR _05648_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30561_ clknet_leaf_219_clk _02296_ VGND VGND VPWR VPWR datamem.data_ram\[54\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32300_ clknet_leaf_160_clk _03722_ VGND VGND VPWR VPWR datamem.data_ram\[32\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_61_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17234_ _04877_ VGND VGND VPWR VPWR _01425_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30492_ clknet_leaf_203_clk _02227_ VGND VGND VPWR VPWR datamem.data_ram\[57\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23712__305 clknet_1_0__leaf__10197_ VGND VGND VPWR VPWR net431 sky130_fd_sc_hd__inv_2
XFILLER_0_101_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32231_ clknet_leaf_86_clk _03653_ VGND VGND VPWR VPWR datamem.data_ram\[35\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17165_ _14151_ net2614 _04840_ VGND VGND VPWR VPWR _04841_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold907 rvcpu.dp.rf.reg_file_arr\[9\]\[10\] VGND VGND VPWR VPWR net2057 sky130_fd_sc_hd__dlygate4sd3_1
X_16116_ _14400_ VGND VGND VPWR VPWR _01966_ sky130_fd_sc_hd__clkbuf_1
Xhold918 rvcpu.dp.rf.reg_file_arr\[24\]\[20\] VGND VGND VPWR VPWR net2068 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32162_ clknet_leaf_272_clk _03584_ VGND VGND VPWR VPWR datamem.data_ram\[38\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold929 rvcpu.dp.rf.reg_file_arr\[9\]\[13\] VGND VGND VPWR VPWR net2079 sky130_fd_sc_hd__dlygate4sd3_1
X_17096_ _04792_ VGND VGND VPWR VPWR _04804_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_229_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31113_ clknet_leaf_58_clk _02848_ VGND VGND VPWR VPWR datamem.data_ram\[43\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16047_ net1888 _13223_ _14360_ VGND VGND VPWR VPWR _14364_ sky130_fd_sc_hd__mux2_1
XFILLER_0_228_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32093_ clknet_leaf_236_clk _03515_ VGND VGND VPWR VPWR datamem.data_ram\[8\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3009 datamem.data_ram\[24\]\[30\] VGND VGND VPWR VPWR net4159 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_62_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31044_ clknet_leaf_73_clk _02779_ VGND VGND VPWR VPWR datamem.data_ram\[41\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2308 datamem.data_ram\[11\]\[9\] VGND VGND VPWR VPWR net3458 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2319 datamem.data_ram\[36\]\[20\] VGND VGND VPWR VPWR net3469 sky130_fd_sc_hd__dlygate4sd3_1
X_19806_ datamem.data_ram\[2\]\[9\] _06691_ _06760_ datamem.data_ram\[7\]\[9\] VGND
+ VGND VPWR VPWR _07101_ sky130_fd_sc_hd__o22a_1
XFILLER_0_23_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1607 datamem.data_ram\[0\]\[10\] VGND VGND VPWR VPWR net2757 sky130_fd_sc_hd__dlygate4sd3_1
X_17998_ _05366_ _05367_ VGND VGND VPWR VPWR _05368_ sky130_fd_sc_hd__nor2b_2
Xhold1618 datamem.data_ram\[39\]\[19\] VGND VGND VPWR VPWR net2768 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1629 datamem.data_ram\[7\]\[20\] VGND VGND VPWR VPWR net2779 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19737_ datamem.data_ram\[3\]\[25\] _06738_ _06700_ datamem.data_ram\[1\]\[25\] _07031_
+ VGND VGND VPWR VPWR _07032_ sky130_fd_sc_hd__o221a_1
X_16949_ net2277 _14432_ _04720_ VGND VGND VPWR VPWR _04726_ sky130_fd_sc_hd__mux2_1
XFILLER_0_224_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_76_clk clknet_5_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_76_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31946_ clknet_leaf_116_clk _03368_ VGND VGND VPWR VPWR datamem.data_ram\[32\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_19668_ _06680_ _06960_ _06963_ VGND VGND VPWR VPWR _06964_ sky130_fd_sc_hd__or3_1
XFILLER_0_177_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18619_ _05790_ _05967_ _05969_ _05976_ VGND VGND VPWR VPWR _05977_ sky130_fd_sc_hd__o211a_1
XFILLER_0_149_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31877_ clknet_leaf_113_clk _03331_ VGND VGND VPWR VPWR datamem.data_ram\[56\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_19599_ datamem.data_ram\[52\]\[8\] _06805_ _06893_ _06894_ VGND VGND VPWR VPWR _06895_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_177_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21630_ _08682_ _08877_ _08879_ VGND VGND VPWR VPWR _08880_ sky130_fd_sc_hd__a21o_1
X_30828_ clknet_leaf_200_clk _02563_ VGND VGND VPWR VPWR datamem.data_ram\[44\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21561_ rvcpu.dp.rf.reg_file_arr\[4\]\[9\] rvcpu.dp.rf.reg_file_arr\[5\]\[9\] rvcpu.dp.rf.reg_file_arr\[6\]\[9\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[9\] _08687_ _08649_ VGND VGND VPWR VPWR _08814_ sky130_fd_sc_hd__mux4_1
XFILLER_0_191_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30759_ clknet_leaf_152_clk _02494_ VGND VGND VPWR VPWR datamem.data_ram\[47\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20512_ datamem.data_ram\[62\]\[21\] _07028_ _06659_ datamem.data_ram\[57\]\[21\]
+ _07802_ VGND VGND VPWR VPWR _07803_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_211_5554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24280_ _09252_ net3760 _10307_ VGND VGND VPWR VPWR _10313_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_211_5565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21492_ _08512_ VGND VGND VPWR VPWR _08748_ sky130_fd_sc_hd__buf_2
XFILLER_0_144_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_209_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23652__252 clknet_1_1__leaf__10181_ VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__inv_2
X_32429_ clknet_leaf_249_clk _03851_ VGND VGND VPWR VPWR datamem.data_ram\[28\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_20443_ _06751_ _07729_ _07734_ VGND VGND VPWR VPWR _07735_ sky130_fd_sc_hd__or3_1
XFILLER_0_71_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24049__577 clknet_1_1__leaf__10246_ VGND VGND VPWR VPWR net703 sky130_fd_sc_hd__inv_2
X_23162_ clknet_1_0__leaf__10108_ VGND VGND VPWR VPWR _10110_ sky130_fd_sc_hd__buf_1
Xclkload350 clknet_1_1__leaf__10091_ VGND VGND VPWR VPWR clkload350/Y sky130_fd_sc_hd__clkinvlp_4
X_20374_ datamem.data_ram\[45\]\[28\] _06722_ _06599_ _07665_ VGND VGND VPWR VPWR
+ _07666_ sky130_fd_sc_hd__o211a_1
XFILLER_0_207_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload80 clknet_leaf_42_clk VGND VGND VPWR VPWR clkload80/Y sky130_fd_sc_hd__bufinv_16
X_22113_ _09321_ VGND VGND VPWR VPWR _09322_ sky130_fd_sc_hd__clkbuf_2
Xclkload91 clknet_leaf_72_clk VGND VGND VPWR VPWR clkload91/Y sky130_fd_sc_hd__inv_6
XFILLER_0_105_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27970_ _12440_ VGND VGND VPWR VPWR _03819_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26921_ _11831_ net1595 _11821_ _11838_ VGND VGND VPWR VPWR _03372_ sky130_fd_sc_hd__a31o_1
X_22044_ rvcpu.dp.plem.WriteDataM\[0\] _09264_ _09265_ rvcpu.dp.plem.WriteDataM\[8\]
+ VGND VGND VPWR VPWR _09266_ sky130_fd_sc_hd__a22o_4
XFILLER_0_227_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_228_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2820 datamem.data_ram\[31\]\[24\] VGND VGND VPWR VPWR net3970 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_167_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29640_ net986 _01375_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[24\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_26852_ _11672_ _11786_ VGND VGND VPWR VPWR _11794_ sky130_fd_sc_hd__and2_1
Xhold2831 datamem.data_ram\[54\]\[12\] VGND VGND VPWR VPWR net3981 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_162_4373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2842 datamem.data_ram\[54\]\[19\] VGND VGND VPWR VPWR net3992 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_162_4384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2853 rvcpu.dp.rf.reg_file_arr\[14\]\[4\] VGND VGND VPWR VPWR net4003 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_162_4395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2864 datamem.data_ram\[63\]\[14\] VGND VGND VPWR VPWR net4014 sky130_fd_sc_hd__dlygate4sd3_1
X_25803_ rvcpu.dp.pcreg.q\[17\] _11191_ VGND VGND VPWR VPWR _11194_ sky130_fd_sc_hd__nand2_1
Xhold2875 datamem.data_ram\[30\]\[19\] VGND VGND VPWR VPWR net4025 sky130_fd_sc_hd__dlygate4sd3_1
X_29571_ net925 _01306_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[26\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_104_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26783_ _11681_ _11749_ VGND VGND VPWR VPWR _11754_ sky130_fd_sc_hd__and2_1
XFILLER_0_199_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2886 datamem.data_ram\[43\]\[9\] VGND VGND VPWR VPWR net4036 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_67_clk clknet_5_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_67_clk sky130_fd_sc_hd__clkbuf_8
Xhold2897 rvcpu.dp.rf.reg_file_arr\[23\]\[9\] VGND VGND VPWR VPWR net4047 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_170_Right_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28522_ _12749_ net2204 _12735_ VGND VGND VPWR VPWR _12750_ sky130_fd_sc_hd__mux2_1
X_22946_ _10073_ _10053_ VGND VGND VPWR VPWR _10074_ sky130_fd_sc_hd__and2_1
X_25734_ _10826_ net2830 _11133_ VGND VGND VPWR VPWR _11141_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_218_5719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23507__152 clknet_1_0__leaf__10161_ VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_175_4701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28453_ _12708_ VGND VGND VPWR VPWR _04034_ sky130_fd_sc_hd__clkbuf_1
X_25665_ _11083_ _11098_ VGND VGND VPWR VPWR _11101_ sky130_fd_sc_hd__and2_1
XFILLER_0_35_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22877_ _09510_ _10006_ _10008_ _10012_ _08589_ VGND VGND VPWR VPWR _10013_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_65_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_121_3391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27404_ _12091_ net3530 net85 VGND VGND VPWR VPWR _12122_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_4609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21828_ rvcpu.dp.rf.reg_file_arr\[8\]\[23\] rvcpu.dp.rf.reg_file_arr\[10\]\[23\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[23\] rvcpu.dp.rf.reg_file_arr\[11\]\[23\] _08560_
+ _08561_ VGND VGND VPWR VPWR _09067_ sky130_fd_sc_hd__mux4_1
X_24616_ _10510_ VGND VGND VPWR VPWR _02395_ sky130_fd_sc_hd__clkbuf_1
X_25596_ _11057_ net1558 _11053_ _11061_ VGND VGND VPWR VPWR _02824_ sky130_fd_sc_hd__a31o_1
X_28384_ _12667_ VGND VGND VPWR VPWR _04006_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24547_ _10470_ net4297 _10466_ VGND VGND VPWR VPWR _10471_ sky130_fd_sc_hd__mux2_1
X_27335_ _12080_ net4093 _12081_ VGND VGND VPWR VPWR _12082_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21759_ _08817_ _08999_ _09001_ _08700_ VGND VGND VPWR VPWR _09002_ sky130_fd_sc_hd__a211o_1
XFILLER_0_38_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15280_ _13412_ _13794_ _13818_ _13791_ VGND VGND VPWR VPWR _13819_ sky130_fd_sc_hd__o211a_1
Xwire101 _10706_ VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__buf_4
XFILLER_0_110_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27266_ _12044_ VGND VGND VPWR VPWR _03511_ sky130_fd_sc_hd__clkbuf_1
X_24478_ _09330_ net3737 _10421_ VGND VGND VPWR VPWR _10429_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29005_ _12995_ net1463 _13009_ _13013_ VGND VGND VPWR VPWR _04281_ sky130_fd_sc_hd__a31o_1
X_26217_ _11446_ VGND VGND VPWR VPWR _03060_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_24_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27197_ _10402_ _10980_ VGND VGND VPWR VPWR _12008_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_130_3605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_3616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_130_3627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_169_4549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26148_ _11410_ VGND VGND VPWR VPWR _03026_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_95_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18970_ _06306_ VGND VGND VPWR VPWR rvcpu.ALUResultE\[27\] sky130_fd_sc_hd__buf_1
X_26079_ _11362_ VGND VGND VPWR VPWR _11371_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_91_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29907_ clknet_leaf_140_clk _01642_ VGND VGND VPWR VPWR datamem.data_ram\[59\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_17921_ _05268_ _05263_ VGND VGND VPWR VPWR _05294_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_128_3556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17852_ _05229_ VGND VGND VPWR VPWR rvcpu.dp.SrcBFW_Mux.y\[11\] sky130_fd_sc_hd__buf_1
X_29838_ net216 _01573_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[18\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_128_3567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_3578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23421__74 clknet_1_0__leaf__10153_ VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__inv_2
XFILLER_0_205_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16803_ net2213 _14420_ _04648_ VGND VGND VPWR VPWR _04649_ sky130_fd_sc_hd__mux2_1
XFILLER_0_227_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_179_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17783_ _05161_ VGND VGND VPWR VPWR _05180_ sky130_fd_sc_hd__buf_2
X_29769_ net1115 _01504_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[20\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14995_ _13414_ _13541_ _13523_ _13542_ VGND VGND VPWR VPWR _13543_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_58_clk clknet_5_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_58_clk sky130_fd_sc_hd__clkbuf_8
X_31800_ clknet_leaf_97_clk _03254_ VGND VGND VPWR VPWR datamem.data_ram\[46\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_50_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19522_ _06810_ _06814_ _06817_ VGND VGND VPWR VPWR _06818_ sky130_fd_sc_hd__and3_1
XFILLER_0_221_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16734_ _04611_ VGND VGND VPWR VPWR _04612_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32780_ clknet_leaf_154_clk _04202_ VGND VGND VPWR VPWR datamem.data_ram\[14\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19453_ _06716_ _06736_ _06748_ VGND VGND VPWR VPWR _06749_ sky130_fd_sc_hd__or3_1
X_31731_ net180 _03189_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[9\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_16665_ _14197_ _04465_ VGND VGND VPWR VPWR _04575_ sky130_fd_sc_hd__nand2_2
X_18404_ _05689_ VGND VGND VPWR VPWR _05768_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_29_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15616_ _14116_ VGND VGND VPWR VPWR _02198_ sky130_fd_sc_hd__clkbuf_1
X_19384_ _06679_ VGND VGND VPWR VPWR _06680_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_202_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31662_ clknet_leaf_70_clk net1258 VGND VGND VPWR VPWR rvcpu.dp.plmw.ALUResultW\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_16596_ rvcpu.dp.plmw.RegWriteW _14346_ rvcpu.dp.plmw.RdW\[1\] VGND VGND VPWR VPWR
+ _04538_ sky130_fd_sc_hd__and3_4
XFILLER_0_173_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30613_ clknet_leaf_148_clk _02348_ VGND VGND VPWR VPWR datamem.data_ram\[52\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_18335_ _05484_ _05490_ _05500_ _05506_ _05666_ _05671_ VGND VGND VPWR VPWR _05700_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_45_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15547_ _14055_ _14058_ _14060_ _14072_ VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__a31oi_4
XFILLER_0_127_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31593_ clknet_leaf_51_clk net1248 VGND VGND VPWR VPWR rvcpu.dp.plmw.PCPlus4W\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30544_ clknet_leaf_141_clk _02279_ VGND VGND VPWR VPWR datamem.data_ram\[55\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_18266_ _05531_ _05537_ _05543_ _05549_ VGND VGND VPWR VPWR _05631_ sky130_fd_sc_hd__nor4_1
X_15478_ _13327_ _13697_ _14006_ _13539_ VGND VGND VPWR VPWR _14007_ sky130_fd_sc_hd__a31o_1
XFILLER_0_167_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17217_ _04868_ VGND VGND VPWR VPWR _01433_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18197_ _05561_ VGND VGND VPWR VPWR _05562_ sky130_fd_sc_hd__inv_2
X_30475_ net153 _02210_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[19\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32214_ clknet_leaf_276_clk _03636_ VGND VGND VPWR VPWR datamem.data_ram\[36\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold704 rvcpu.dp.plfd.PCD\[6\] VGND VGND VPWR VPWR net1854 sky130_fd_sc_hd__dlygate4sd3_1
X_17148_ _14135_ net2626 _04829_ VGND VGND VPWR VPWR _04832_ sky130_fd_sc_hd__mux2_1
Xhold715 rvcpu.dp.rf.reg_file_arr\[17\]\[25\] VGND VGND VPWR VPWR net1865 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold726 rvcpu.dp.rf.reg_file_arr\[17\]\[16\] VGND VGND VPWR VPWR net1876 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold737 rvcpu.dp.plem.ALUResultM\[6\] VGND VGND VPWR VPWR net1887 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32145_ clknet_leaf_226_clk _03567_ VGND VGND VPWR VPWR datamem.data_ram\[38\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold748 rvcpu.dp.rf.reg_file_arr\[9\]\[31\] VGND VGND VPWR VPWR net1898 sky130_fd_sc_hd__dlygate4sd3_1
Xhold759 rvcpu.dp.plfd.InstrD\[31\] VGND VGND VPWR VPWR net1909 sky130_fd_sc_hd__dlygate4sd3_1
X_17079_ _04795_ VGND VGND VPWR VPWR _01498_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32076_ clknet_leaf_114_clk _03498_ VGND VGND VPWR VPWR datamem.data_ram\[33\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20090_ datamem.data_ram\[62\]\[10\] _06627_ _06723_ datamem.data_ram\[61\]\[10\]
+ VGND VGND VPWR VPWR _07384_ sky130_fd_sc_hd__o22a_1
XFILLER_0_196_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2105 datamem.data_ram\[16\]\[18\] VGND VGND VPWR VPWR net3255 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2116 datamem.data_ram\[0\]\[12\] VGND VGND VPWR VPWR net3266 sky130_fd_sc_hd__dlygate4sd3_1
X_31027_ clknet_leaf_61_clk _02762_ VGND VGND VPWR VPWR datamem.data_ram\[40\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2127 datamem.data_ram\[2\]\[27\] VGND VGND VPWR VPWR net3277 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2138 datamem.data_ram\[43\]\[11\] VGND VGND VPWR VPWR net3288 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2149 datamem.data_ram\[30\]\[9\] VGND VGND VPWR VPWR net3299 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1404 rvcpu.dp.rf.reg_file_arr\[6\]\[11\] VGND VGND VPWR VPWR net2554 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1415 datamem.data_ram\[59\]\[10\] VGND VGND VPWR VPWR net2565 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_204_5380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1300 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_204_5391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23682__278 clknet_1_0__leaf__10194_ VGND VGND VPWR VPWR net404 sky130_fd_sc_hd__inv_2
Xhold1426 datamem.data_ram\[4\]\[29\] VGND VGND VPWR VPWR net2576 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1437 rvcpu.dp.rf.reg_file_arr\[14\]\[12\] VGND VGND VPWR VPWR net2587 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1448 datamem.data_ram\[29\]\[31\] VGND VGND VPWR VPWR net2598 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_49_clk clknet_5_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_49_clk sky130_fd_sc_hd__clkbuf_8
Xhold1459 rvcpu.dp.rf.reg_file_arr\[5\]\[24\] VGND VGND VPWR VPWR net2609 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22800_ _09495_ _09939_ VGND VGND VPWR VPWR _09940_ sky130_fd_sc_hd__nor2_1
XFILLER_0_224_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_200_5288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32978_ clknet_leaf_176_clk _04400_ VGND VGND VPWR VPWR datamem.data_ram\[63\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_20992_ datamem.data_ram\[6\]\[15\] datamem.data_ram\[7\]\[15\] _06651_ VGND VGND
+ VPWR VPWR _08281_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_200_5299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_196_5192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22731_ _09870_ _09874_ rvcpu.dp.plfd.InstrD\[24\] VGND VGND VPWR VPWR _09875_ sky130_fd_sc_hd__o21a_1
X_31929_ clknet_leaf_122_clk _03351_ VGND VGND VPWR VPWR datamem.data_ram\[60\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25450_ _10058_ _10981_ _10982_ net1358 VGND VGND VPWR VPWR _02757_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22662_ rvcpu.dp.rf.reg_file_arr\[8\]\[18\] rvcpu.dp.rf.reg_file_arr\[10\]\[18\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[18\] rvcpu.dp.rf.reg_file_arr\[11\]\[18\] _09608_
+ _09656_ VGND VGND VPWR VPWR _09810_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_213_5605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_213_5616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_1238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31749__126 VGND VGND VPWR VPWR _31749__126/HI net126 sky130_fd_sc_hd__conb_1
XFILLER_0_149_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24401_ _09279_ net3275 _10376_ VGND VGND VPWR VPWR _10380_ sky130_fd_sc_hd__mux2_1
X_21613_ _08672_ _08854_ _08859_ _08863_ VGND VGND VPWR VPWR _08864_ sky130_fd_sc_hd__and4_1
X_25381_ _10938_ net1394 _10934_ _10942_ VGND VGND VPWR VPWR _02728_ sky130_fd_sc_hd__a31o_1
XFILLER_0_164_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22593_ rvcpu.dp.rf.reg_file_arr\[20\]\[15\] rvcpu.dp.rf.reg_file_arr\[21\]\[15\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[15\] rvcpu.dp.rf.reg_file_arr\[23\]\[15\] _09401_
+ _09430_ VGND VGND VPWR VPWR _09744_ sky130_fd_sc_hd__mux4_1
XFILLER_0_63_703 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27120_ _11946_ _11953_ VGND VGND VPWR VPWR _11959_ sky130_fd_sc_hd__and2_1
X_24332_ _10342_ VGND VGND VPWR VPWR _02279_ sky130_fd_sc_hd__clkbuf_1
X_21544_ _08673_ _08796_ VGND VGND VPWR VPWR _08797_ sky130_fd_sc_hd__or2_1
XFILLER_0_173_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27051_ _11803_ _11911_ VGND VGND VPWR VPWR _11916_ sky130_fd_sc_hd__and2_1
XFILLER_0_105_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24263_ _09322_ net2941 _10298_ VGND VGND VPWR VPWR _10304_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21475_ rvcpu.dp.rf.reg_file_arr\[12\]\[5\] rvcpu.dp.rf.reg_file_arr\[13\]\[5\] rvcpu.dp.rf.reg_file_arr\[14\]\[5\]
+ rvcpu.dp.rf.reg_file_arr\[15\]\[5\] _08551_ _08555_ VGND VGND VPWR VPWR _08732_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_105_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26002_ net15 _11317_ VGND VGND VPWR VPWR _11326_ sky130_fd_sc_hd__or2_1
XFILLER_0_209_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23214_ clknet_1_1__leaf__10108_ VGND VGND VPWR VPWR _10124_ sky130_fd_sc_hd__buf_1
XFILLER_0_71_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20426_ datamem.data_ram\[0\]\[12\] _06647_ _07716_ _07717_ VGND VGND VPWR VPWR _07718_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20357_ datamem.data_ram\[10\]\[28\] _06690_ _06725_ datamem.data_ram\[15\]\[28\]
+ VGND VGND VPWR VPWR _07649_ sky130_fd_sc_hd__o22a_1
Xclkload180 clknet_leaf_236_clk VGND VGND VPWR VPWR clkload180/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_105_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload191 clknet_leaf_225_clk VGND VGND VPWR VPWR clkload191/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_164_4424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_164_4435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27953_ _12371_ net2598 _12421_ VGND VGND VPWR VPWR _12429_ sky130_fd_sc_hd__mux2_1
X_23076_ _09288_ net2633 _10093_ VGND VGND VPWR VPWR _10100_ sky130_fd_sc_hd__mux2_1
X_20288_ datamem.data_ram\[22\]\[19\] _06629_ _06779_ datamem.data_ram\[16\]\[19\]
+ VGND VGND VPWR VPWR _07581_ sky130_fd_sc_hd__o22a_1
XFILLER_0_11_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26904_ _10060_ VGND VGND VPWR VPWR _11827_ sky130_fd_sc_hd__clkbuf_4
X_22027_ _09251_ VGND VGND VPWR VPWR _09252_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_41_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_216_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27884_ _11918_ VGND VGND VPWR VPWR _12391_ sky130_fd_sc_hd__buf_2
Xhold20 rvcpu.dp.plem.lAuiPCM\[7\] VGND VGND VPWR VPWR net1170 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 rvcpu.dp.plem.lAuiPCM\[17\] VGND VGND VPWR VPWR net1181 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 rvcpu.dp.plem.lAuiPCM\[29\] VGND VGND VPWR VPWR net1192 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2650 datamem.data_ram\[22\]\[25\] VGND VGND VPWR VPWR net3800 sky130_fd_sc_hd__dlygate4sd3_1
X_29623_ net977 _01358_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[25\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26835_ _07182_ _10918_ _10897_ VGND VGND VPWR VPWR _11784_ sky130_fd_sc_hd__or3_1
Xhold53 rvcpu.dp.plem.lAuiPCM\[0\] VGND VGND VPWR VPWR net1203 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2661 datamem.data_ram\[9\]\[17\] VGND VGND VPWR VPWR net3811 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 rvcpu.dp.plem.lAuiPCM\[9\] VGND VGND VPWR VPWR net1214 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2672 datamem.data_ram\[16\]\[12\] VGND VGND VPWR VPWR net3822 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_67_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2683 rvcpu.dp.rf.reg_file_arr\[17\]\[4\] VGND VGND VPWR VPWR net3833 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold75 rvcpu.dp.plem.PCPlus4M\[19\] VGND VGND VPWR VPWR net1225 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_67_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2694 datamem.data_ram\[46\]\[26\] VGND VGND VPWR VPWR net3844 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 rvcpu.dp.plem.PCPlus4M\[5\] VGND VGND VPWR VPWR net1236 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1960 rvcpu.dp.rf.reg_file_arr\[14\]\[20\] VGND VGND VPWR VPWR net3110 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold97 rvcpu.dp.plem.PCPlus4M\[7\] VGND VGND VPWR VPWR net1247 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_123_3442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29554_ net908 _01289_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[27\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_26766_ _11645_ _11738_ VGND VGND VPWR VPWR _11743_ sky130_fd_sc_hd__and2_1
XFILLER_0_199_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14780_ _13332_ VGND VGND VPWR VPWR _13333_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_123_3453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1971 datamem.data_ram\[42\]\[13\] VGND VGND VPWR VPWR net3121 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1982 rvcpu.dp.rf.reg_file_arr\[14\]\[2\] VGND VGND VPWR VPWR net3132 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_199_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1993 rvcpu.dp.rf.reg_file_arr\[30\]\[12\] VGND VGND VPWR VPWR net3143 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_168_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28505_ _12738_ VGND VGND VPWR VPWR _04056_ sky130_fd_sc_hd__clkbuf_1
X_25717_ _10826_ net1996 _11124_ VGND VGND VPWR VPWR _11132_ sky130_fd_sc_hd__mux2_1
X_22929_ _10060_ VGND VGND VPWR VPWR _10061_ sky130_fd_sc_hd__buf_2
Xclkbuf_1_1__f__10266_ clknet_0__10266_ VGND VGND VPWR VPWR clknet_1_1__leaf__10266_
+ sky130_fd_sc_hd__clkbuf_16
X_29485_ net847 _01220_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[2\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_26697_ _11672_ _11694_ VGND VGND VPWR VPWR _11703_ sky130_fd_sc_hd__and2_1
XFILLER_0_196_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_711 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28436_ _09321_ VGND VGND VPWR VPWR _12698_ sky130_fd_sc_hd__clkbuf_2
X_16450_ net1980 _14480_ _04451_ VGND VGND VPWR VPWR _04460_ sky130_fd_sc_hd__mux2_1
X_25648_ _10600_ _11075_ VGND VGND VPWR VPWR _11094_ sky130_fd_sc_hd__nor2_2
X_23659__258 clknet_1_1__leaf__10191_ VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__10197_ clknet_0__10197_ VGND VGND VPWR VPWR clknet_1_1__leaf__10197_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_128_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15401_ _13496_ _13523_ _13368_ VGND VGND VPWR VPWR _13933_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_26_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16381_ _14555_ VGND VGND VPWR VPWR _01848_ sky130_fd_sc_hd__clkbuf_1
X_28367_ _12658_ VGND VGND VPWR VPWR _03998_ sky130_fd_sc_hd__clkbuf_1
X_25579_ _11018_ net1539 _11041_ _11050_ VGND VGND VPWR VPWR _02818_ sky130_fd_sc_hd__a31o_1
XFILLER_0_183_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18120_ _05484_ _05485_ VGND VGND VPWR VPWR _05487_ sky130_fd_sc_hd__nand2_1
X_15332_ _13366_ _13308_ _13598_ _13868_ VGND VGND VPWR VPWR _13869_ sky130_fd_sc_hd__o31a_1
X_27318_ _11980_ _12066_ VGND VGND VPWR VPWR _12074_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_22_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28298_ _12621_ VGND VGND VPWR VPWR _03966_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_22_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18051_ _13253_ _05271_ VGND VGND VPWR VPWR _05420_ sky130_fd_sc_hd__and2_1
X_15263_ _13366_ _13416_ _13671_ _13799_ _13802_ VGND VGND VPWR VPWR _13803_ sky130_fd_sc_hd__o311a_1
X_27249_ _12036_ net1579 _12030_ _12038_ VGND VGND VPWR VPWR _03500_ sky130_fd_sc_hd__a31o_1
XFILLER_0_163_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_227_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17002_ _04753_ VGND VGND VPWR VPWR _01541_ sky130_fd_sc_hd__clkbuf_1
X_15194_ _13539_ _13725_ _13732_ _13736_ VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__a22o_1
XANTENNA_6 _05622_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30260_ net614 _01995_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[6\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24145__649 clknet_1_1__leaf__10262_ VGND VGND VPWR VPWR net775 sky130_fd_sc_hd__inv_2
XFILLER_0_111_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30191_ net545 _01926_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[8\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18953_ _05240_ _06279_ _06281_ _06055_ _06290_ VGND VGND VPWR VPWR rvcpu.ALUResultE\[26\]
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_123_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23824__406 clknet_1_0__leaf__10208_ VGND VGND VPWR VPWR net532 sky130_fd_sc_hd__inv_2
X_17904_ _05276_ VGND VGND VPWR VPWR _05277_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_123_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18884_ _05467_ _06225_ VGND VGND VPWR VPWR _06226_ sky130_fd_sc_hd__xor2_1
XFILLER_0_158_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_52_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_271 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32901_ clknet_leaf_236_clk _04323_ VGND VGND VPWR VPWR datamem.data_ram\[0\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17835_ rvcpu.dp.plem.ALUResultM\[21\] _05217_ _05177_ VGND VGND VPWR VPWR _05218_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23904__463 clknet_1_1__leaf__10223_ VGND VGND VPWR VPWR net589 sky130_fd_sc_hd__inv_2
XFILLER_0_83_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32832_ clknet_leaf_190_clk _04254_ VGND VGND VPWR VPWR datamem.data_ram\[12\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_222_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17766_ _05162_ rvcpu.dp.plde.Rs2E\[0\] _05163_ VGND VGND VPWR VPWR _05164_ sky130_fd_sc_hd__o21ai_1
X_14978_ _13287_ _13281_ VGND VGND VPWR VPWR _13526_ sky130_fd_sc_hd__nand2_4
X_19505_ datamem.data_ram\[54\]\[24\] _06682_ _06790_ datamem.data_ram\[49\]\[24\]
+ _06800_ VGND VGND VPWR VPWR _06801_ sky130_fd_sc_hd__o221a_1
XFILLER_0_221_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16717_ _14181_ net4062 _04598_ VGND VGND VPWR VPWR _04603_ sky130_fd_sc_hd__mux2_1
X_32763_ clknet_leaf_255_clk _04185_ VGND VGND VPWR VPWR datamem.data_ram\[15\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17697_ _13195_ net3153 _05118_ VGND VGND VPWR VPWR _05123_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19436_ _06676_ VGND VGND VPWR VPWR _06732_ sky130_fd_sc_hd__buf_8
X_31714_ net163 _03172_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[9\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_16648_ _04566_ VGND VGND VPWR VPWR _01716_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32694_ clknet_leaf_283_clk _04116_ VGND VGND VPWR VPWR datamem.data_ram\[18\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23718__311 clknet_1_0__leaf__10197_ VGND VGND VPWR VPWR net437 sky130_fd_sc_hd__inv_2
XFILLER_0_85_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31645_ clknet_leaf_27_clk net1164 VGND VGND VPWR VPWR rvcpu.dp.plmw.lAuiPCW\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19367_ _06662_ VGND VGND VPWR VPWR _06663_ sky130_fd_sc_hd__buf_8
X_16579_ _04529_ VGND VGND VPWR VPWR _01756_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18318_ _05682_ VGND VGND VPWR VPWR _05683_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19298_ _06593_ VGND VGND VPWR VPWR _06594_ sky130_fd_sc_hd__buf_8
X_31576_ clknet_leaf_72_clk datamem.rd_data_mem\[26\] VGND VGND VPWR VPWR rvcpu.dp.plmw.ReadDataW\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18249_ _05318_ _05613_ VGND VGND VPWR VPWR _05614_ sky130_fd_sc_hd__or2_1
XFILLER_0_142_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30527_ clknet_leaf_266_clk _02262_ VGND VGND VPWR VPWR datamem.data_ram\[56\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21260_ rvcpu.dp.plfd.InstrD\[17\] VGND VGND VPWR VPWR _08522_ sky130_fd_sc_hd__inv_2
XFILLER_0_206_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold501 rvcpu.dp.plfd.PCD\[29\] VGND VGND VPWR VPWR net1651 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30458_ net136 _02193_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[19\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold512 datamem.data_ram\[31\]\[5\] VGND VGND VPWR VPWR net1662 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold523 datamem.data_ram\[27\]\[4\] VGND VGND VPWR VPWR net1673 sky130_fd_sc_hd__dlygate4sd3_1
X_20211_ _06716_ _07487_ _07492_ _07503_ VGND VGND VPWR VPWR _07504_ sky130_fd_sc_hd__o31a_1
Xhold534 datamem.data_ram\[50\]\[3\] VGND VGND VPWR VPWR net1684 sky130_fd_sc_hd__dlygate4sd3_1
Xhold545 datamem.data_ram\[1\]\[1\] VGND VGND VPWR VPWR net1695 sky130_fd_sc_hd__dlygate4sd3_1
X_21191_ _06915_ _07368_ _07413_ _07277_ VGND VGND VPWR VPWR _08476_ sky130_fd_sc_hd__o22a_1
XFILLER_0_29_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold556 datamem.data_ram\[62\]\[0\] VGND VGND VPWR VPWR net1706 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30389_ net727 _02124_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[31\]\[0\] sky130_fd_sc_hd__dfxtp_1
Xhold567 datamem.data_ram\[17\]\[0\] VGND VGND VPWR VPWR net1717 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_206_5431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold578 rvcpu.dp.plfd.PCPlus4D\[15\] VGND VGND VPWR VPWR net1728 sky130_fd_sc_hd__dlygate4sd3_1
X_20142_ datamem.data_ram\[43\]\[27\] _06828_ _07434_ _06851_ VGND VGND VPWR VPWR
+ _07435_ sky130_fd_sc_hd__o211a_1
X_32128_ clknet_leaf_194_clk _03550_ VGND VGND VPWR VPWR datamem.data_ram\[7\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold589 datamem.data_ram\[24\]\[2\] VGND VGND VPWR VPWR net1739 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_206_5442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23152__825 clknet_1_0__leaf__10109_ VGND VGND VPWR VPWR net951 sky130_fd_sc_hd__inv_2
X_23764__353 clknet_1_1__leaf__10201_ VGND VGND VPWR VPWR net479 sky130_fd_sc_hd__inv_2
XFILLER_0_110_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32059_ clknet_leaf_133_clk _03481_ VGND VGND VPWR VPWR datamem.data_ram\[48\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_24950_ _10452_ net2773 _10687_ VGND VGND VPWR VPWR _10694_ sky130_fd_sc_hd__mux2_1
X_20073_ _07177_ _07328_ _07333_ _07366_ VGND VGND VPWR VPWR _07367_ sky130_fd_sc_hd__o31a_4
XTAP_TAPCELL_ROW_202_5339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1201 rvcpu.dp.rf.reg_file_arr\[6\]\[16\] VGND VGND VPWR VPWR net2351 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_198_5243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1212 rvcpu.dp.rf.reg_file_arr\[16\]\[16\] VGND VGND VPWR VPWR net2362 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_198_5254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1223 rvcpu.dp.rf.reg_file_arr\[14\]\[15\] VGND VGND VPWR VPWR net2373 sky130_fd_sc_hd__dlygate4sd3_1
X_24881_ _10478_ net1933 _10650_ VGND VGND VPWR VPWR _10657_ sky130_fd_sc_hd__mux2_1
Xhold1234 rvcpu.dp.rf.reg_file_arr\[25\]\[28\] VGND VGND VPWR VPWR net2384 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1245 rvcpu.dp.rf.reg_file_arr\[3\]\[25\] VGND VGND VPWR VPWR net2395 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1256 datamem.data_ram\[18\]\[14\] VGND VGND VPWR VPWR net2406 sky130_fd_sc_hd__dlygate4sd3_1
X_26620_ _10826_ net2029 _11650_ VGND VGND VPWR VPWR _11658_ sky130_fd_sc_hd__mux2_1
X_23879__440 clknet_1_0__leaf__10221_ VGND VGND VPWR VPWR net566 sky130_fd_sc_hd__inv_2
Xhold1267 rvcpu.dp.rf.reg_file_arr\[3\]\[16\] VGND VGND VPWR VPWR net2417 sky130_fd_sc_hd__dlygate4sd3_1
X_23832_ _10212_ VGND VGND VPWR VPWR _01909_ sky130_fd_sc_hd__clkbuf_1
Xhold1278 rvcpu.dp.rf.reg_file_arr\[0\]\[20\] VGND VGND VPWR VPWR net2428 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1289 datamem.data_ram\[30\]\[23\] VGND VGND VPWR VPWR net2439 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__10220_ _10220_ VGND VGND VPWR VPWR clknet_0__10220_ sky130_fd_sc_hd__clkbuf_16
XANTENNA_407 _06645_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_212_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_418 _06751_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_603 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26551_ _10570_ _11123_ _10998_ VGND VGND VPWR VPWR _11620_ sky130_fd_sc_hd__a21oi_4
X_20975_ _08262_ _08263_ _07819_ VGND VGND VPWR VPWR _08264_ sky130_fd_sc_hd__mux2_1
XANTENNA_429 _06790_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25502_ _10824_ net3620 _10999_ VGND VGND VPWR VPWR _11006_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22714_ rvcpu.dp.rf.reg_file_arr\[12\]\[21\] rvcpu.dp.rf.reg_file_arr\[13\]\[21\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[21\] rvcpu.dp.rf.reg_file_arr\[15\]\[21\] _09386_
+ _09419_ VGND VGND VPWR VPWR _09859_ sky130_fd_sc_hd__mux4_1
XFILLER_0_71_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29270_ _09284_ net3700 _13150_ VGND VGND VPWR VPWR _13156_ sky130_fd_sc_hd__mux2_1
X_26482_ _11252_ _11153_ _11599_ _11600_ _10780_ VGND VGND VPWR VPWR _03171_ sky130_fd_sc_hd__a221oi_1
XTAP_TAPCELL_ROW_157_4261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_157_4272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28221_ _12579_ VGND VGND VPWR VPWR _03931_ sky130_fd_sc_hd__clkbuf_1
X_25433_ _10756_ net4008 _10970_ VGND VGND VPWR VPWR _10973_ sky130_fd_sc_hd__mux2_1
X_22645_ _09534_ _09793_ VGND VGND VPWR VPWR _09794_ sky130_fd_sc_hd__and2_1
Xclkbuf_0__10082_ _10082_ VGND VGND VPWR VPWR clknet_0__10082_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_165_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_153_4158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25364_ _10076_ _10923_ VGND VGND VPWR VPWR _10931_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_153_4169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28152_ _12542_ VGND VGND VPWR VPWR _03899_ sky130_fd_sc_hd__clkbuf_1
X_22576_ _09726_ _09727_ _09449_ VGND VGND VPWR VPWR _09728_ sky130_fd_sc_hd__mux2_1
XFILLER_0_192_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27103_ _11938_ net1885 _11940_ _11948_ VGND VGND VPWR VPWR _03444_ sky130_fd_sc_hd__a31o_1
XFILLER_0_8_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24315_ _09318_ net2644 _10328_ VGND VGND VPWR VPWR _10333_ sky130_fd_sc_hd__mux2_1
X_21527_ rvcpu.dp.rf.reg_file_arr\[28\]\[8\] rvcpu.dp.rf.reg_file_arr\[30\]\[8\] rvcpu.dp.rf.reg_file_arr\[29\]\[8\]
+ rvcpu.dp.rf.reg_file_arr\[31\]\[8\] _08635_ _08637_ VGND VGND VPWR VPWR _08781_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25295_ _10890_ VGND VGND VPWR VPWR _02694_ sky130_fd_sc_hd__clkbuf_1
X_28083_ _12439_ net3261 _12501_ VGND VGND VPWR VPWR _12506_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_1221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27034_ _11833_ _11899_ VGND VGND VPWR VPWR _11906_ sky130_fd_sc_hd__and2_1
X_23470__118 clknet_1_0__leaf__10158_ VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__inv_2
X_24246_ _10294_ VGND VGND VPWR VPWR _02241_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_3290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21458_ _08663_ _08713_ _08715_ _08575_ VGND VGND VPWR VPWR _08716_ sky130_fd_sc_hd__o211a_1
XFILLER_0_161_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_189_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20409_ _06601_ _07698_ _07700_ VGND VGND VPWR VPWR _07701_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_187_4980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput8 net8 VGND VGND VPWR VPWR Instr[15] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_187_4991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput10 net10 VGND VGND VPWR VPWR Instr[17] sky130_fd_sc_hd__buf_2
X_21389_ rvcpu.dp.rf.reg_file_arr\[8\]\[1\] rvcpu.dp.rf.reg_file_arr\[10\]\[1\] rvcpu.dp.rf.reg_file_arr\[9\]\[1\]
+ rvcpu.dp.rf.reg_file_arr\[11\]\[1\] _08649_ _08537_ VGND VGND VPWR VPWR _08650_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_222_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput21 net21 VGND VGND VPWR VPWR Instr[27] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_112_3187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput32 net32 VGND VGND VPWR VPWR Instr[8] sky130_fd_sc_hd__buf_2
XFILLER_0_222_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23128_ clknet_1_0__leaf__10087_ VGND VGND VPWR VPWR _10106_ sky130_fd_sc_hd__buf_1
XFILLER_0_208_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28985_ _12692_ net3182 _12999_ VGND VGND VPWR VPWR _13002_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_183_4877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_4888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23092__772 clknet_1_0__leaf__10102_ VGND VGND VPWR VPWR net898 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_183_4899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27936_ _12140_ net4380 _12412_ VGND VGND VPWR VPWR _12420_ sky130_fd_sc_hd__mux2_1
X_15950_ rvcpu.dp.rf.reg_file_arr\[5\]\[31\] _13173_ _14311_ VGND VGND VPWR VPWR _14312_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_125_3504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23014__718 clknet_1_1__leaf__10086_ VGND VGND VPWR VPWR net844 sky130_fd_sc_hd__inv_2
Xhold3170 rvcpu.dp.rf.reg_file_arr\[23\]\[11\] VGND VGND VPWR VPWR net4320 sky130_fd_sc_hd__dlygate4sd3_1
X_14901_ _13448_ _13450_ _13451_ _13333_ VGND VGND VPWR VPWR _13452_ sky130_fd_sc_hd__a31o_1
Xhold3181 rvcpu.dp.rf.reg_file_arr\[2\]\[7\] VGND VGND VPWR VPWR net4331 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3192 datamem.data_ram\[35\]\[7\] VGND VGND VPWR VPWR net4342 sky130_fd_sc_hd__dlygate4sd3_1
X_27867_ _10668_ _12345_ _12356_ VGND VGND VPWR VPWR _12382_ sky130_fd_sc_hd__a21oi_2
X_15881_ _14274_ VGND VGND VPWR VPWR _14275_ sky130_fd_sc_hd__clkbuf_4
X_29606_ net960 _01341_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[25\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_17620_ _05081_ VGND VGND VPWR VPWR _05082_ sky130_fd_sc_hd__buf_4
Xhold2480 datamem.data_ram\[40\]\[13\] VGND VGND VPWR VPWR net3630 sky130_fd_sc_hd__dlygate4sd3_1
X_26818_ _11676_ _11774_ VGND VGND VPWR VPWR _11775_ sky130_fd_sc_hd__and2_1
X_14832_ _13314_ VGND VGND VPWR VPWR _13385_ sky130_fd_sc_hd__clkbuf_4
Xhold2491 datamem.data_ram\[21\]\[30\] VGND VGND VPWR VPWR net3641 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27798_ _12134_ net2502 _12336_ VGND VGND VPWR VPWR _12341_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_86_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23129__805 clknet_1_0__leaf__10106_ VGND VGND VPWR VPWR net931 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_86_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_3895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29537_ net891 _01272_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[27\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_17551_ _14129_ _04464_ VGND VGND VPWR VPWR _05045_ sky130_fd_sc_hd__nand2_2
Xhold1790 datamem.data_ram\[51\]\[11\] VGND VGND VPWR VPWR net2940 sky130_fd_sc_hd__dlygate4sd3_1
X_26749_ _11700_ net1709 _11724_ _11732_ VGND VGND VPWR VPWR _03306_ sky130_fd_sc_hd__a31o_1
X_14763_ _13290_ _13310_ _13315_ VGND VGND VPWR VPWR _13316_ sky130_fd_sc_hd__a21oi_1
X_16502_ _04488_ VGND VGND VPWR VPWR _01792_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_224_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17482_ _05008_ VGND VGND VPWR VPWR _01300_ sky130_fd_sc_hd__clkbuf_1
X_29468_ net830 _01203_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[2\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14694_ _13255_ VGND VGND VPWR VPWR _03180_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_224_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19221_ rvcpu.dp.plde.ImmExtE\[26\] rvcpu.dp.plde.PCE\[26\] VGND VGND VPWR VPWR _06528_
+ sky130_fd_sc_hd__or2_1
X_16433_ _14560_ VGND VGND VPWR VPWR _04451_ sky130_fd_sc_hd__clkbuf_4
X_28419_ _12686_ VGND VGND VPWR VPWR _04022_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_15_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29399_ clknet_leaf_0_clk _01134_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD2E\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_15_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19152_ _06465_ _06467_ VGND VGND VPWR VPWR _06468_ sky130_fd_sc_hd__xnor2_1
X_31430_ clknet_leaf_61_clk _03133_ VGND VGND VPWR VPWR datamem.data_ram\[44\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16364_ _14546_ VGND VGND VPWR VPWR _01856_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23934__489 clknet_1_1__leaf__10227_ VGND VGND VPWR VPWR net615 sky130_fd_sc_hd__inv_2
XFILLER_0_229_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18103_ _05469_ _05470_ VGND VGND VPWR VPWR _05471_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15315_ _13542_ _13851_ VGND VGND VPWR VPWR _13852_ sky130_fd_sc_hd__nor2_1
X_19083_ rvcpu.dp.plde.ImmExtE\[9\] rvcpu.dp.plde.PCE\[9\] VGND VGND VPWR VPWR _06407_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_186_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31361_ clknet_leaf_22_clk _03064_ VGND VGND VPWR VPWR rvcpu.dp.plde.ImmExtE\[10\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_14_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16295_ net2835 _14461_ _14500_ VGND VGND VPWR VPWR _14510_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18034_ _05368_ _05401_ _05403_ _05366_ VGND VGND VPWR VPWR _05404_ sky130_fd_sc_hd__a211o_1
X_30312_ net658 _02047_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[5\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_15246_ _13358_ _13432_ _13488_ _13685_ _13598_ VGND VGND VPWR VPWR _13786_ sky130_fd_sc_hd__o32a_1
X_31292_ clknet_leaf_22_clk _02995_ VGND VGND VPWR VPWR rvcpu.dp.plde.JalrE sky130_fd_sc_hd__dfxtp_2
XFILLER_0_164_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__10140_ clknet_0__10140_ VGND VGND VPWR VPWR clknet_1_0__leaf__10140_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_152_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30243_ net597 _01978_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[7\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_15177_ _13346_ _13391_ _13483_ _13298_ VGND VGND VPWR VPWR _13720_ sky130_fd_sc_hd__a211o_1
XFILLER_0_2_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19985_ datamem.data_ram\[10\]\[2\] _06930_ _06946_ datamem.data_ram\[9\]\[2\] VGND
+ VGND VPWR VPWR _07279_ sky130_fd_sc_hd__a22o_1
X_30174_ clknet_leaf_207_clk _01909_ VGND VGND VPWR VPWR datamem.data_ram\[58\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23216__866 clknet_1_1__leaf__10124_ VGND VGND VPWR VPWR net992 sky130_fd_sc_hd__inv_2
XFILLER_0_10_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18936_ _05661_ _06027_ _06273_ _05703_ _06274_ VGND VGND VPWR VPWR _06275_ sky130_fd_sc_hd__a221o_1
XFILLER_0_123_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_105_Left_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18867_ _05481_ _06194_ _05479_ VGND VGND VPWR VPWR _06210_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_222_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17818_ _05206_ VGND VGND VPWR VPWR rvcpu.dp.SrcBFW_Mux.y\[27\] sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_27_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18798_ _05511_ _05784_ _05974_ _05510_ VGND VGND VPWR VPWR _06146_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_55_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32815_ clknet_leaf_282_clk _04237_ VGND VGND VPWR VPWR datamem.data_ram\[13\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_17749_ _13272_ net3575 _05140_ VGND VGND VPWR VPWR _05150_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20760_ datamem.data_ram\[2\]\[6\] _07837_ _08049_ _07636_ VGND VGND VPWR VPWR _08050_
+ sky130_fd_sc_hd__o211a_1
X_32746_ clknet_leaf_184_clk _04168_ VGND VGND VPWR VPWR datamem.data_ram\[15\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19419_ _06714_ VGND VGND VPWR VPWR _06715_ sky130_fd_sc_hd__buf_8
XFILLER_0_134_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23794__379 clknet_1_1__leaf__10205_ VGND VGND VPWR VPWR net505 sky130_fd_sc_hd__inv_2
XFILLER_0_147_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20691_ datamem.data_ram\[61\]\[5\] _06969_ _06955_ datamem.data_ram\[60\]\[5\] VGND
+ VGND VPWR VPWR _07982_ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32677_ clknet_leaf_240_clk _04099_ VGND VGND VPWR VPWR datamem.data_ram\[18\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_114_Left_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_77_Right_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22430_ rvcpu.dp.rf.reg_file_arr\[8\]\[6\] rvcpu.dp.rf.reg_file_arr\[10\]\[6\] rvcpu.dp.rf.reg_file_arr\[9\]\[6\]
+ rvcpu.dp.rf.reg_file_arr\[11\]\[6\] _09431_ _09532_ VGND VGND VPWR VPWR _09590_
+ sky130_fd_sc_hd__mux4_1
X_31628_ clknet_leaf_48_clk net1238 VGND VGND VPWR VPWR rvcpu.dp.plmw.lAuiPCW\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22361_ _09451_ _09520_ _09522_ _09523_ VGND VGND VPWR VPWR _09524_ sky130_fd_sc_hd__o211a_1
XFILLER_0_190_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31559_ clknet_leaf_71_clk datamem.rd_data_mem\[9\] VGND VGND VPWR VPWR rvcpu.dp.plmw.ReadDataW\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23449__99 clknet_1_1__leaf__10156_ VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__inv_2
XFILLER_0_142_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21312_ _08572_ _08573_ VGND VGND VPWR VPWR _08574_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25080_ _10771_ VGND VGND VPWR VPWR _02598_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22292_ _09404_ VGND VGND VPWR VPWR _09457_ sky130_fd_sc_hd__buf_4
XFILLER_0_5_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold320 datamem.data_ram\[20\]\[5\] VGND VGND VPWR VPWR net1470 sky130_fd_sc_hd__dlygate4sd3_1
X_21243_ datamem.data_ram\[53\]\[2\] datamem.data_ram\[52\]\[26\] datamem.data_ram\[52\]\[18\]
+ datamem.data_ram\[52\]\[2\] VGND VGND VPWR VPWR _08506_ sky130_fd_sc_hd__and4b_1
Xhold331 datamem.data_ram\[60\]\[1\] VGND VGND VPWR VPWR net1481 sky130_fd_sc_hd__dlygate4sd3_1
Xhold342 datamem.data_ram\[23\]\[7\] VGND VGND VPWR VPWR net1492 sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 datamem.data_ram\[59\]\[0\] VGND VGND VPWR VPWR net1503 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold364 datamem.data_ram\[28\]\[4\] VGND VGND VPWR VPWR net1514 sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 datamem.data_ram\[34\]\[4\] VGND VGND VPWR VPWR net1525 sky130_fd_sc_hd__dlygate4sd3_1
X_21174_ _06714_ _08447_ _08462_ _07177_ VGND VGND VPWR VPWR _08463_ sky130_fd_sc_hd__a22o_1
X_23688__284 clknet_1_1__leaf__10194_ VGND VGND VPWR VPWR net410 sky130_fd_sc_hd__inv_2
XFILLER_0_111_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold386 datamem.data_ram\[12\]\[1\] VGND VGND VPWR VPWR net1536 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold397 datamem.data_ram\[28\]\[2\] VGND VGND VPWR VPWR net1547 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_123_Left_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_86_Right_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_229_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_225_5884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_280_clk clknet_5_24__leaf_clk VGND VGND VPWR VPWR clknet_leaf_280_clk
+ sky130_fd_sc_hd__clkbuf_8
X_20125_ datamem.data_ram\[5\]\[27\] _06664_ _06648_ datamem.data_ram\[0\]\[27\] _07417_
+ VGND VGND VPWR VPWR _07418_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_225_5895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28770_ _12885_ VGND VGND VPWR VPWR _04174_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_176_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25982_ rvcpu.dp.plfd.InstrD\[12\] _11302_ _11312_ _11314_ VGND VGND VPWR VPWR _02957_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27721_ _12299_ VGND VGND VPWR VPWR _03711_ sky130_fd_sc_hd__clkbuf_1
X_24933_ _10478_ net2560 _10678_ VGND VGND VPWR VPWR _10685_ sky130_fd_sc_hd__mux2_1
X_20056_ datamem.data_ram\[42\]\[26\] _06609_ _06704_ datamem.data_ram\[47\]\[26\]
+ _07349_ VGND VGND VPWR VPWR _07350_ sky130_fd_sc_hd__o221a_1
XFILLER_0_77_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1020 rvcpu.dp.rf.reg_file_arr\[12\]\[31\] VGND VGND VPWR VPWR net2170 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1031 rvcpu.dp.rf.reg_file_arr\[9\]\[5\] VGND VGND VPWR VPWR net2181 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_175_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1042 datamem.data_ram\[49\]\[15\] VGND VGND VPWR VPWR net2192 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27652_ _12262_ VGND VGND VPWR VPWR _03679_ sky130_fd_sc_hd__clkbuf_1
Xhold1053 datamem.data_ram\[19\]\[30\] VGND VGND VPWR VPWR net2203 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_159_4301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24864_ _10398_ net2217 _10641_ VGND VGND VPWR VPWR _10648_ sky130_fd_sc_hd__mux2_1
XFILLER_0_217_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_159_4312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1064 datamem.data_ram\[1\]\[31\] VGND VGND VPWR VPWR net2214 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1075 rvcpu.dp.rf.reg_file_arr\[10\]\[13\] VGND VGND VPWR VPWR net2225 sky130_fd_sc_hd__dlygate4sd3_1
X_26603_ _11064_ _11640_ VGND VGND VPWR VPWR _11649_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_159_4323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1086 rvcpu.dp.rf.reg_file_arr\[17\]\[30\] VGND VGND VPWR VPWR net2236 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1097 rvcpu.dp.rf.reg_file_arr\[8\]\[10\] VGND VGND VPWR VPWR net2247 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_204 _09526_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27583_ _12225_ VGND VGND VPWR VPWR _03647_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_215 _09750_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_23__f_clk clknet_2_2_0_clk VGND VGND VPWR VPWR clknet_5_23__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_24795_ _10480_ net2901 net94 VGND VGND VPWR VPWR _10610_ sky130_fd_sc_hd__mux2_1
XANTENNA_226 _10066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_0__10203_ _10203_ VGND VGND VPWR VPWR clknet_0__10203_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_96_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29322_ clknet_leaf_12_clk _01057_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD1E\[29\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_237 _10388_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_1_1__f__10103_ clknet_0__10103_ VGND VGND VPWR VPWR clknet_1_1__leaf__10103_
+ sky130_fd_sc_hd__clkbuf_16
X_26534_ _11078_ _11610_ VGND VGND VPWR VPWR _11611_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_155_4209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_248 _13176_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20958_ datamem.data_ram\[53\]\[15\] _06660_ _06616_ datamem.data_ram\[52\]\[15\]
+ _08246_ VGND VGND VPWR VPWR _08247_ sky130_fd_sc_hd__o221a_1
XANTENNA_259 _13207_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_132_Left_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_191_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0__10134_ _10134_ VGND VGND VPWR VPWR clknet_0__10134_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_95_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_95_Right_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29253_ _09251_ net3765 _13141_ VGND VGND VPWR VPWR _13147_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26465_ rvcpu.dp.pcreg.q\[26\] _11573_ _11588_ _11570_ VGND VGND VPWR VPWR _03166_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_166_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20889_ _08173_ _08178_ _08124_ VGND VGND VPWR VPWR _08179_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_193_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28204_ _12458_ net3718 net46 VGND VGND VPWR VPWR _12570_ sky130_fd_sc_hd__mux2_1
X_25416_ _10756_ net3874 _10961_ VGND VGND VPWR VPWR _10964_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_118_3330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_187_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29184_ _13109_ VGND VGND VPWR VPWR _04364_ sky130_fd_sc_hd__clkbuf_1
X_22628_ _09777_ VGND VGND VPWR VPWR _01140_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23321__961 clknet_1_0__leaf__10134_ VGND VGND VPWR VPWR net1087 sky130_fd_sc_hd__inv_2
X_26396_ _11539_ VGND VGND VPWR VPWR _11540_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_64_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28135_ _12533_ VGND VGND VPWR VPWR _03891_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25347_ _10051_ VGND VGND VPWR VPWR _10921_ sky130_fd_sc_hd__buf_2
X_22559_ _09399_ _09711_ _09472_ VGND VGND VPWR VPWR _09712_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_114_3227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15100_ _13393_ _13523_ _13470_ VGND VGND VPWR VPWR _13645_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_114_3238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28066_ _12365_ net3466 _12492_ VGND VGND VPWR VPWR _12497_ sky130_fd_sc_hd__mux2_1
X_16080_ net2154 _13272_ _14371_ VGND VGND VPWR VPWR _14381_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25278_ _10881_ VGND VGND VPWR VPWR _02686_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_79_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_185_4928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15031_ _13424_ _13577_ VGND VGND VPWR VPWR _13578_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_185_4939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27017_ _11837_ _11886_ VGND VGND VPWR VPWR _11895_ sky130_fd_sc_hd__and2_1
X_24229_ _10285_ VGND VGND VPWR VPWR _02233_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_224_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_141_Left_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_271_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_271_clk
+ sky130_fd_sc_hd__clkbuf_8
X_19770_ datamem.data_ram\[29\]\[25\] _06768_ _06760_ datamem.data_ram\[31\]\[25\]
+ VGND VGND VPWR VPWR _07065_ sky130_fd_sc_hd__o22a_1
X_28968_ _12727_ net1495 _12988_ _12992_ VGND VGND VPWR VPWR _04265_ sky130_fd_sc_hd__a31o_1
X_16982_ _04743_ VGND VGND VPWR VPWR _01551_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_88_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18721_ _05436_ _05727_ _05730_ _05434_ VGND VGND VPWR VPWR _06073_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27919_ _12157_ net2183 net47 VGND VGND VPWR VPWR _12411_ sky130_fd_sc_hd__mux2_1
X_15933_ _14302_ VGND VGND VPWR VPWR _02059_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_144_3946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28899_ _12954_ VGND VGND VPWR VPWR _04234_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_204_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30930_ clknet_leaf_137_clk _02665_ VGND VGND VPWR VPWR datamem.data_ram\[40\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_18652_ _05696_ _06007_ VGND VGND VPWR VPWR _06008_ sky130_fd_sc_hd__nand2_1
X_15864_ _14264_ VGND VGND VPWR VPWR _02090_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_204_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_192_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17603_ _13257_ net3189 _05068_ VGND VGND VPWR VPWR _05073_ sky130_fd_sc_hd__mux2_1
X_14815_ _13312_ VGND VGND VPWR VPWR _13368_ sky130_fd_sc_hd__buf_4
X_18583_ _05360_ _05784_ _05732_ _05402_ VGND VGND VPWR VPWR _05942_ sky130_fd_sc_hd__o22a_1
X_30861_ clknet_leaf_264_clk _02596_ VGND VGND VPWR VPWR datamem.data_ram\[43\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15795_ _14227_ VGND VGND VPWR VPWR _02130_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_192_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_150_Left_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32600_ clknet_leaf_274_clk _04022_ VGND VGND VPWR VPWR datamem.data_ram\[21\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_17534_ _05036_ VGND VGND VPWR VPWR _01276_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_47_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14746_ _13286_ rvcpu.dp.pcreg.q\[3\] VGND VGND VPWR VPWR _13299_ sky130_fd_sc_hd__and2_1
XFILLER_0_114_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30792_ clknet_leaf_260_clk _02527_ VGND VGND VPWR VPWR datamem.data_ram\[46\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_103_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_1107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32531_ clknet_leaf_240_clk _03953_ VGND VGND VPWR VPWR datamem.data_ram\[23\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_103_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17465_ _14179_ net3105 _04996_ VGND VGND VPWR VPWR _05000_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14677_ _13242_ VGND VGND VPWR VPWR _03184_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19204_ _06513_ VGND VGND VPWR VPWR rvcpu.dp.lAuiPCE\[23\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16416_ _14574_ VGND VGND VPWR VPWR _01832_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_184_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32462_ clknet_leaf_246_clk _03884_ VGND VGND VPWR VPWR datamem.data_ram\[26\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_17396_ _04963_ VGND VGND VPWR VPWR _01341_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19135_ _06451_ _06452_ VGND VGND VPWR VPWR _06453_ sky130_fd_sc_hd__xnor2_1
X_31413_ clknet_leaf_23_clk _03116_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCE\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16347_ net1985 _14445_ _14536_ VGND VGND VPWR VPWR _14538_ sky130_fd_sc_hd__mux2_1
X_32393_ clknet_leaf_76_clk _03815_ VGND VGND VPWR VPWR datamem.data_ram\[29\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19066_ _06392_ rvcpu.dp.plde.ImmExtE\[6\] _06355_ VGND VGND VPWR VPWR _06393_ sky130_fd_sc_hd__mux2_1
X_31344_ clknet_leaf_19_clk _03047_ VGND VGND VPWR VPWR rvcpu.dp.plde.ALUControlE\[0\]
+ sky130_fd_sc_hd__dfxtp_2
X_23099__778 clknet_1_0__leaf__10103_ VGND VGND VPWR VPWR net904 sky130_fd_sc_hd__inv_2
XFILLER_0_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16278_ _14501_ VGND VGND VPWR VPWR _01897_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18017_ _05386_ _05293_ VGND VGND VPWR VPWR _05387_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15229_ _13439_ _13581_ _13766_ _13769_ VGND VGND VPWR VPWR _13770_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_112_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31275_ clknet_leaf_126_clk _02978_ VGND VGND VPWR VPWR datamem.data_ram\[24\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30226_ net580 _01961_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[7\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_262_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_262_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_61_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout118 _00000_ VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__buf_2
XFILLER_0_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30157_ net519 _01892_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[0\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_19968_ _06602_ _07259_ _07261_ VGND VGND VPWR VPWR _07262_ sky130_fd_sc_hd__and3_1
X_18919_ _05866_ _06031_ _06138_ _06137_ VGND VGND VPWR VPWR _06259_ sky130_fd_sc_hd__o31a_1
XFILLER_0_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30088_ net450 _01823_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[11\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_19899_ datamem.data_ram\[2\]\[17\] _06612_ _06863_ datamem.data_ram\[3\]\[17\] _06776_
+ VGND VGND VPWR VPWR _07194_ sky130_fd_sc_hd__o221a_1
XFILLER_0_207_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_220_5770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_220_5781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21930_ _09161_ _09162_ _08673_ VGND VGND VPWR VPWR _09163_ sky130_fd_sc_hd__mux2_1
X_24174__15 clknet_1_1__leaf__10265_ VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__inv_2
XFILLER_0_59_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21861_ _08523_ _09097_ _08748_ VGND VGND VPWR VPWR _09098_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23802__386 clknet_1_1__leaf__10206_ VGND VGND VPWR VPWR net512 sky130_fd_sc_hd__inv_2
XFILLER_0_136_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20812_ datamem.data_ram\[59\]\[30\] _06940_ _06934_ datamem.data_ram\[57\]\[30\]
+ VGND VGND VPWR VPWR _08102_ sky130_fd_sc_hd__o22a_1
XFILLER_0_136_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24580_ _10490_ VGND VGND VPWR VPWR _02379_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21792_ _08835_ _09032_ VGND VGND VPWR VPWR _09033_ sky130_fd_sc_hd__or2_1
XFILLER_0_65_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20743_ rvcpu.dp.plem.ALUResultM\[4\] datamem.data_ram\[46\]\[6\] _07821_ _07836_
+ VGND VGND VPWR VPWR _08033_ sky130_fd_sc_hd__a31o_1
XFILLER_0_147_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32729_ clknet_leaf_79_clk _04151_ VGND VGND VPWR VPWR datamem.data_ram\[16\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26250_ _11438_ _11458_ _11459_ net1315 VGND VGND VPWR VPWR _03080_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_135_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20674_ _07920_ net36 _06911_ VGND VGND VPWR VPWR _07965_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_150_4106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_189_5028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23043__744 clknet_1_0__leaf__10089_ VGND VGND VPWR VPWR net870 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_189_5039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25201_ _10838_ _10601_ _10828_ VGND VGND VPWR VPWR _10839_ sky130_fd_sc_hd__a21oi_1
X_22413_ _09476_ _09571_ _09573_ _09489_ VGND VGND VPWR VPWR _09574_ sky130_fd_sc_hd__o211a_1
XFILLER_0_174_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26181_ _11427_ VGND VGND VPWR VPWR _03043_ sky130_fd_sc_hd__clkbuf_1
X_23393_ _10147_ VGND VGND VPWR VPWR _01535_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25132_ _10474_ net4212 net87 VGND VGND VPWR VPWR _10798_ sky130_fd_sc_hd__mux2_1
X_22344_ _09482_ _09507_ VGND VGND VPWR VPWR _09508_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23158__831 clknet_1_0__leaf__10109_ VGND VGND VPWR VPWR net957 sky130_fd_sc_hd__inv_2
XFILLER_0_27_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25063_ _10760_ net3786 _10752_ VGND VGND VPWR VPWR _10761_ sky130_fd_sc_hd__mux2_1
X_29940_ net310 _01675_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[16\]\[31\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_227_5935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22275_ _09440_ VGND VGND VPWR VPWR _01124_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_227_5946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_148_4046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold150 rvcpu.dp.plfd.InstrD\[29\] VGND VGND VPWR VPWR net1300 sky130_fd_sc_hd__dlygate4sd3_1
X_21226_ _08468_ _08123_ _08489_ VGND VGND VPWR VPWR _04438_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_148_4057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29871_ net249 _01606_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[17\]\[2\] sky130_fd_sc_hd__dfxtp_1
Xhold161 datamem.data_ram\[41\]\[1\] VGND VGND VPWR VPWR net1311 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold172 datamem.data_ram\[43\]\[7\] VGND VGND VPWR VPWR net1322 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold183 datamem.data_ram\[45\]\[0\] VGND VGND VPWR VPWR net1333 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_180_4814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold194 datamem.data_ram\[44\]\[2\] VGND VGND VPWR VPWR net1344 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_180_4825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_253_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_253_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_40_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28822_ _12913_ VGND VGND VPWR VPWR _04198_ sky130_fd_sc_hd__clkbuf_1
X_21157_ _07862_ _08442_ _08445_ _06598_ VGND VGND VPWR VPWR _08446_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_6_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20108_ datamem.data_ram\[22\]\[10\] _06717_ _06669_ datamem.data_ram\[23\]\[10\]
+ VGND VGND VPWR VPWR _07402_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_70_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28753_ _12876_ VGND VGND VPWR VPWR _04166_ sky130_fd_sc_hd__clkbuf_1
X_21088_ datamem.data_ram\[53\]\[7\] _06918_ _06923_ datamem.data_ram\[55\]\[7\] _08376_
+ VGND VGND VPWR VPWR _08377_ sky130_fd_sc_hd__a221o_1
X_25965_ net28 _11153_ _11300_ _11305_ VGND VGND VPWR VPWR _02949_ sky130_fd_sc_hd__o211a_1
XFILLER_0_176_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27704_ _12290_ VGND VGND VPWR VPWR _03703_ sky130_fd_sc_hd__clkbuf_1
X_24916_ _10398_ net1903 _10669_ VGND VGND VPWR VPWR _10676_ sky130_fd_sc_hd__mux2_1
X_20039_ datamem.data_ram\[19\]\[26\] _06635_ _07329_ _07332_ VGND VGND VPWR VPWR
+ _07333_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_107_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28684_ _12766_ net2561 _12832_ VGND VGND VPWR VPWR _12840_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25896_ net1854 _11263_ VGND VGND VPWR VPWR _11266_ sky130_fd_sc_hd__or2_1
XFILLER_0_198_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27635_ _12128_ net3043 _12251_ VGND VGND VPWR VPWR _12253_ sky130_fd_sc_hd__mux2_1
X_24847_ _10638_ VGND VGND VPWR VPWR _02498_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_178_4765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_4776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14600_ _13183_ VGND VGND VPWR VPWR _13184_ sky130_fd_sc_hd__buf_4
X_27566_ _12216_ VGND VGND VPWR VPWR _03639_ sky130_fd_sc_hd__clkbuf_1
X_15580_ _14097_ VGND VGND VPWR VPWR _02215_ sky130_fd_sc_hd__clkbuf_1
X_24778_ _10599_ VGND VGND VPWR VPWR _10600_ sky130_fd_sc_hd__buf_8
XFILLER_0_29_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29305_ clknet_leaf_0_clk _01040_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD1E\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_185_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26517_ _07132_ _10050_ VGND VGND VPWR VPWR _11603_ sky130_fd_sc_hd__nand2_4
XFILLER_0_200_269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27497_ _12142_ net3371 _12179_ VGND VGND VPWR VPWR _12180_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17250_ _04885_ VGND VGND VPWR VPWR _01417_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_42_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29236_ _09321_ net2368 _13132_ VGND VGND VPWR VPWR _13138_ sky130_fd_sc_hd__mux2_1
X_26448_ _11524_ rvcpu.ALUResultE\[21\] _11288_ VGND VGND VPWR VPWR _11577_ sky130_fd_sc_hd__a21o_1
XFILLER_0_154_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23476__124 clknet_1_1__leaf__10158_ VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__inv_2
XFILLER_0_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_3772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16201_ _14452_ VGND VGND VPWR VPWR _01933_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_181_655 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29167_ _13100_ VGND VGND VPWR VPWR _04356_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_3783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17181_ _14168_ net3028 _04840_ VGND VGND VPWR VPWR _04849_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26379_ _11524_ rvcpu.ALUResultE\[2\] _11148_ _11526_ VGND VGND VPWR VPWR _11527_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_137_3794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28118_ _12524_ VGND VGND VPWR VPWR _03883_ sky130_fd_sc_hd__clkbuf_1
X_16132_ net2317 _13248_ _14407_ VGND VGND VPWR VPWR _14409_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29098_ _09321_ net3572 net40 VGND VGND VPWR VPWR _13064_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28049_ _12456_ net4224 net96 VGND VGND VPWR VPWR _12488_ sky130_fd_sc_hd__mux2_1
X_16063_ _14372_ VGND VGND VPWR VPWR _01991_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_219_Left_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15014_ rvcpu.dp.pcreg.q\[5\] _13281_ VGND VGND VPWR VPWR _13562_ sky130_fd_sc_hd__nor2_2
X_31060_ clknet_leaf_90_clk _02795_ VGND VGND VPWR VPWR datamem.data_ram\[38\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_184_Right_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_244_clk clknet_5_17__leaf_clk VGND VGND VPWR VPWR clknet_leaf_244_clk
+ sky130_fd_sc_hd__clkbuf_8
X_30011_ clknet_leaf_174_clk _01746_ VGND VGND VPWR VPWR datamem.data_ram\[59\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_19822_ _07107_ _07108_ _07111_ _07116_ VGND VGND VPWR VPWR _07117_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_36_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16965_ _04734_ VGND VGND VPWR VPWR _01559_ sky130_fd_sc_hd__clkbuf_1
X_19753_ datamem.data_ram\[61\]\[25\] _07037_ _06657_ datamem.data_ram\[57\]\[25\]
+ VGND VGND VPWR VPWR _07048_ sky130_fd_sc_hd__o22a_1
XFILLER_0_223_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18704_ _05607_ _06041_ _05410_ VGND VGND VPWR VPWR _06057_ sky130_fd_sc_hd__a21o_1
X_15916_ _14293_ VGND VGND VPWR VPWR _02067_ sky130_fd_sc_hd__clkbuf_1
X_19684_ datamem.data_ram\[56\]\[0\] _06936_ _06947_ datamem.data_ram\[57\]\[0\] VGND
+ VGND VPWR VPWR _06980_ sky130_fd_sc_hd__a22o_1
X_31962_ clknet_leaf_122_clk _03384_ VGND VGND VPWR VPWR datamem.data_ram\[28\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_1166 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16896_ net2378 _14447_ _04695_ VGND VGND VPWR VPWR _04698_ sky130_fd_sc_hd__mux2_1
X_18635_ _05985_ _05991_ _05805_ VGND VGND VPWR VPWR _05992_ sky130_fd_sc_hd__a21oi_1
X_30913_ clknet_leaf_261_clk _02648_ VGND VGND VPWR VPWR datamem.data_ram\[41\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15847_ _14255_ VGND VGND VPWR VPWR _02098_ sky130_fd_sc_hd__clkbuf_1
X_31893_ clknet_leaf_113_clk _03347_ VGND VGND VPWR VPWR datamem.data_ram\[36\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_228_Left_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23328__967 clknet_1_1__leaf__10135_ VGND VGND VPWR VPWR net1093 sky130_fd_sc_hd__inv_2
XFILLER_0_91_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18566_ _05752_ _05762_ _05674_ VGND VGND VPWR VPWR _05926_ sky130_fd_sc_hd__mux2_1
X_30844_ clknet_leaf_172_clk _02579_ VGND VGND VPWR VPWR datamem.data_ram\[44\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_15778_ _14218_ VGND VGND VPWR VPWR _02138_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17517_ _05027_ VGND VGND VPWR VPWR _01284_ sky130_fd_sc_hd__clkbuf_1
X_14729_ _13281_ VGND VGND VPWR VPWR _13282_ sky130_fd_sc_hd__buf_2
XFILLER_0_47_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18497_ _05776_ _05854_ _05857_ _05858_ VGND VGND VPWR VPWR _05859_ sky130_fd_sc_hd__a2bb2o_1
X_30775_ clknet_leaf_202_clk _02510_ VGND VGND VPWR VPWR datamem.data_ram\[46\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32514_ clknet_leaf_81_clk _03936_ VGND VGND VPWR VPWR datamem.data_ram\[24\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17448_ _14162_ net3912 _04985_ VGND VGND VPWR VPWR _04991_ sky130_fd_sc_hd__mux2_1
X_23107__785 clknet_1_1__leaf__10104_ VGND VGND VPWR VPWR net911 sky130_fd_sc_hd__inv_2
XFILLER_0_55_650 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32445_ clknet_leaf_78_clk _03867_ VGND VGND VPWR VPWR datamem.data_ram\[27\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17379_ _04954_ VGND VGND VPWR VPWR _01349_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19118_ _06436_ _06437_ VGND VGND VPWR VPWR _06438_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20390_ datamem.data_ram\[16\]\[28\] _06646_ _06705_ datamem.data_ram\[23\]\[28\]
+ VGND VGND VPWR VPWR _07682_ sky130_fd_sc_hd__o22a_1
XFILLER_0_67_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32376_ clknet_leaf_279_clk _03798_ VGND VGND VPWR VPWR datamem.data_ram\[2\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_19049_ _06377_ rvcpu.dp.plde.ImmExtE\[4\] _06355_ VGND VGND VPWR VPWR _06378_ sky130_fd_sc_hd__mux2_1
X_31327_ clknet_leaf_24_clk _03030_ VGND VGND VPWR VPWR rvcpu.dp.plde.funct3E\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_30_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22060_ _09278_ VGND VGND VPWR VPWR _09279_ sky130_fd_sc_hd__buf_2
X_31258_ clknet_leaf_15_clk _02961_ VGND VGND VPWR VPWR rvcpu.dp.plfd.InstrD\[16\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_140_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__10106_ clknet_0__10106_ VGND VGND VPWR VPWR clknet_1_0__leaf__10106_
+ sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_151_Right_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_235_clk clknet_5_20__leaf_clk VGND VGND VPWR VPWR clknet_leaf_235_clk
+ sky130_fd_sc_hd__clkbuf_8
X_21011_ datamem.data_ram\[62\]\[31\] datamem.data_ram\[63\]\[31\] _07912_ VGND VGND
+ VPWR VPWR _08300_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30209_ net563 _01944_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[8\]\[28\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_222_5821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_222_5832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31189_ clknet_leaf_38_clk _02892_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCPlus4D\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25750_ _13335_ _13717_ VGND VGND VPWR VPWR _11154_ sky130_fd_sc_hd__nand2_1
XFILLER_0_173_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24701_ _10450_ net4321 _10552_ VGND VGND VPWR VPWR _10558_ sky130_fd_sc_hd__mux2_1
X_21913_ rvcpu.dp.rf.reg_file_arr\[24\]\[28\] rvcpu.dp.rf.reg_file_arr\[25\]\[28\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[28\] rvcpu.dp.rf.reg_file_arr\[27\]\[28\] _08549_
+ _08553_ VGND VGND VPWR VPWR _09147_ sky130_fd_sc_hd__mux4_1
X_25681_ _11110_ VGND VGND VPWR VPWR _11111_ sky130_fd_sc_hd__clkbuf_2
X_22893_ rvcpu.dp.rf.reg_file_arr\[24\]\[31\] rvcpu.dp.rf.reg_file_arr\[25\]\[31\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[31\] rvcpu.dp.rf.reg_file_arr\[27\]\[31\] _08592_
+ _08595_ VGND VGND VPWR VPWR _10028_ sky130_fd_sc_hd__mux4_1
XFILLER_0_223_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27420_ _09243_ VGND VGND VPWR VPWR _12132_ sky130_fd_sc_hd__clkbuf_2
X_24632_ _10454_ net2173 _10511_ VGND VGND VPWR VPWR _10519_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21844_ _08513_ _09075_ _09077_ _09079_ _09081_ VGND VGND VPWR VPWR _09082_ sky130_fd_sc_hd__o32a_1
XFILLER_0_210_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_194_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27351_ _12092_ VGND VGND VPWR VPWR _03548_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_176_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21775_ rvcpu.dp.rf.reg_file_arr\[8\]\[20\] rvcpu.dp.rf.reg_file_arr\[10\]\[20\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[20\] rvcpu.dp.rf.reg_file_arr\[11\]\[20\] _08534_
+ _08818_ VGND VGND VPWR VPWR _09017_ sky130_fd_sc_hd__mux4_1
XFILLER_0_93_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24563_ _10481_ VGND VGND VPWR VPWR _02371_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_216_5669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_4640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_4651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26302_ net1692 _11478_ VGND VGND VPWR VPWR _11484_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20726_ datamem.data_ram\[22\]\[6\] _07159_ _06927_ datamem.data_ram\[23\]\[6\] _07081_
+ VGND VGND VPWR VPWR _08016_ sky130_fd_sc_hd__a221o_1
X_23514_ _10165_ VGND VGND VPWR VPWR _01638_ sky130_fd_sc_hd__clkbuf_1
X_27282_ _12052_ VGND VGND VPWR VPWR _12053_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_175_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24494_ _10437_ VGND VGND VPWR VPWR _02346_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1088 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29021_ _13022_ VGND VGND VPWR VPWR _04288_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26233_ _03029_ _11379_ _11454_ VGND VGND VPWR VPWR _03066_ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20657_ datamem.data_ram\[46\]\[29\] _06627_ _06805_ datamem.data_ram\[44\]\[29\]
+ VGND VGND VPWR VPWR _07948_ sky130_fd_sc_hd__o22a_1
XFILLER_0_123_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_208_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26164_ net4447 _11408_ VGND VGND VPWR VPWR _11419_ sky130_fd_sc_hd__and2_1
XFILLER_0_150_327 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20588_ datamem.data_ram\[53\]\[13\] _06703_ _06620_ datamem.data_ram\[52\]\[13\]
+ _07878_ VGND VGND VPWR VPWR _07879_ sky130_fd_sc_hd__o221a_1
XFILLER_0_116_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25115_ _10733_ net3650 net88 VGND VGND VPWR VPWR _10789_ sky130_fd_sc_hd__mux2_1
XFILLER_0_225_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22327_ _09460_ _09475_ _09490_ _09491_ VGND VGND VPWR VPWR _01125_ sky130_fd_sc_hd__o31a_1
X_26095_ _11382_ VGND VGND VPWR VPWR _03001_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_182_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25046_ _10749_ VGND VGND VPWR VPWR _02586_ sky130_fd_sc_hd__clkbuf_1
X_29923_ net293 _01658_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[16\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_22258_ _09400_ VGND VGND VPWR VPWR _09424_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_218_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_4499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21209_ rvcpu.dp.plem.funct3M\[2\] _06580_ VGND VGND VPWR VPWR _08488_ sky130_fd_sc_hd__or2_4
Xclkbuf_leaf_226_clk clknet_5_21__leaf_clk VGND VGND VPWR VPWR clknet_leaf_226_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_143_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29854_ net232 _01589_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[18\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22189_ _09248_ net3965 _09362_ VGND VGND VPWR VPWR _09367_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_109_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28805_ _12904_ VGND VGND VPWR VPWR _04190_ sky130_fd_sc_hd__clkbuf_1
X_29785_ net1131 _01520_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[20\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_26997_ _10766_ net3298 _11875_ VGND VGND VPWR VPWR _11883_ sky130_fd_sc_hd__mux2_1
X_28736_ _12867_ VGND VGND VPWR VPWR _04158_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_31_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16750_ _04620_ VGND VGND VPWR VPWR _01668_ sky130_fd_sc_hd__clkbuf_1
X_25948_ net1588 _11155_ VGND VGND VPWR VPWR _11296_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_31_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_219_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15701_ _14171_ VGND VGND VPWR VPWR _02168_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_220_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16681_ _14145_ net3511 _04576_ VGND VGND VPWR VPWR _04584_ sky130_fd_sc_hd__mux2_1
X_28667_ _12702_ net3944 _12823_ VGND VGND VPWR VPWR _12831_ sky130_fd_sc_hd__mux2_1
X_25879_ _11255_ VGND VGND VPWR VPWR _02913_ sky130_fd_sc_hd__clkbuf_1
X_18420_ _05783_ VGND VGND VPWR VPWR _05784_ sky130_fd_sc_hd__buf_2
XFILLER_0_9_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27618_ _12083_ net3333 net80 VGND VGND VPWR VPWR _12244_ sky130_fd_sc_hd__mux2_1
X_15632_ _14124_ VGND VGND VPWR VPWR _02190_ sky130_fd_sc_hd__clkbuf_1
X_28598_ _12749_ net3571 _12786_ VGND VGND VPWR VPWR _12794_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_100_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18351_ _05677_ _05715_ _05694_ VGND VGND VPWR VPWR _05716_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_139_3823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15563_ _13466_ _14081_ _14086_ _13904_ VGND VGND VPWR VPWR _14087_ sky130_fd_sc_hd__o211a_1
XFILLER_0_186_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_3834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27549_ _12207_ VGND VGND VPWR VPWR _03631_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24072__598 clknet_1_1__leaf__10248_ VGND VGND VPWR VPWR net724 sky130_fd_sc_hd__inv_2
X_17302_ net3005 _13212_ _04913_ VGND VGND VPWR VPWR _04914_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_29_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18282_ _05305_ _05562_ _05641_ _05646_ VGND VGND VPWR VPWR _05647_ sky130_fd_sc_hd__a31o_1
XFILLER_0_126_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30560_ clknet_leaf_219_clk _02295_ VGND VGND VPWR VPWR datamem.data_ram\[54\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_15494_ _13800_ _13893_ _13475_ VGND VGND VPWR VPWR _14022_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29219_ _10069_ _13123_ VGND VGND VPWR VPWR _13129_ sky130_fd_sc_hd__and2_1
XFILLER_0_126_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17233_ _14151_ net2165 _04876_ VGND VGND VPWR VPWR _04877_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30491_ clknet_leaf_195_clk _02226_ VGND VGND VPWR VPWR datamem.data_ram\[57\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_32230_ clknet_leaf_88_clk _03652_ VGND VGND VPWR VPWR datamem.data_ram\[35\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_17164_ _04828_ VGND VGND VPWR VPWR _04840_ sky130_fd_sc_hd__buf_4
XFILLER_0_52_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16115_ net2359 _13223_ _14396_ VGND VGND VPWR VPWR _14400_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32161_ clknet_leaf_241_clk _03583_ VGND VGND VPWR VPWR datamem.data_ram\[38\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold908 datamem.data_ram\[37\]\[31\] VGND VGND VPWR VPWR net2058 sky130_fd_sc_hd__dlygate4sd3_1
Xhold919 rvcpu.dp.rf.reg_file_arr\[14\]\[19\] VGND VGND VPWR VPWR net2069 sky130_fd_sc_hd__dlygate4sd3_1
X_17095_ _04803_ VGND VGND VPWR VPWR _01490_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31112_ clknet_leaf_59_clk _02847_ VGND VGND VPWR VPWR datamem.data_ram\[43\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_16046_ _14363_ VGND VGND VPWR VPWR _01999_ sky130_fd_sc_hd__clkbuf_1
X_32092_ clknet_leaf_234_clk _03514_ VGND VGND VPWR VPWR datamem.data_ram\[8\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_217_clk clknet_5_21__leaf_clk VGND VGND VPWR VPWR clknet_leaf_217_clk
+ sky130_fd_sc_hd__clkbuf_8
X_31043_ clknet_leaf_84_clk _02778_ VGND VGND VPWR VPWR datamem.data_ram\[41\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2309 datamem.data_ram\[9\]\[13\] VGND VGND VPWR VPWR net3459 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19805_ datamem.data_ram\[8\]\[9\] _06698_ _06739_ datamem.data_ram\[11\]\[9\] _07099_
+ VGND VGND VPWR VPWR _07100_ sky130_fd_sc_hd__o221a_1
X_17997_ _05363_ _05365_ VGND VGND VPWR VPWR _05367_ sky130_fd_sc_hd__nand2_1
Xhold1608 rvcpu.dp.rf.reg_file_arr\[31\]\[27\] VGND VGND VPWR VPWR net2758 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_193_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1619 rvcpu.dp.rf.reg_file_arr\[20\]\[8\] VGND VGND VPWR VPWR net2769 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19736_ _06769_ VGND VGND VPWR VPWR _07031_ sky130_fd_sc_hd__buf_8
X_16948_ _04725_ VGND VGND VPWR VPWR _01567_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_223_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32994_ net13 VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_1
XFILLER_0_223_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31945_ clknet_leaf_115_clk _03367_ VGND VGND VPWR VPWR datamem.data_ram\[32\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_19667_ datamem.data_ram\[45\]\[0\] _06920_ _06961_ datamem.data_ram\[43\]\[0\] _06962_
+ VGND VGND VPWR VPWR _06963_ sky130_fd_sc_hd__a221o_1
XFILLER_0_126_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16879_ net3802 _14430_ _04684_ VGND VGND VPWR VPWR _04689_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_205_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18618_ _05782_ _05971_ _05973_ _05975_ VGND VGND VPWR VPWR _05976_ sky130_fd_sc_hd__o211a_1
X_31876_ clknet_leaf_123_clk _03330_ VGND VGND VPWR VPWR datamem.data_ram\[56\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_23261__907 clknet_1_0__leaf__10128_ VGND VGND VPWR VPWR net1033 sky130_fd_sc_hd__inv_2
X_19598_ datamem.data_ram\[50\]\[8\] _06609_ _06780_ datamem.data_ram\[49\]\[8\] _06677_
+ VGND VGND VPWR VPWR _06894_ sky130_fd_sc_hd__o221a_1
XFILLER_0_59_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30827_ clknet_leaf_194_clk _02562_ VGND VGND VPWR VPWR datamem.data_ram\[44\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_18549_ _05909_ VGND VGND VPWR VPWR rvcpu.ALUResultE\[3\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_34_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_191_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21560_ _08540_ VGND VGND VPWR VPWR _08813_ sky130_fd_sc_hd__clkbuf_4
X_30758_ clknet_leaf_156_clk _02493_ VGND VGND VPWR VPWR datamem.data_ram\[47\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20511_ datamem.data_ram\[61\]\[21\] _06665_ _06636_ datamem.data_ram\[59\]\[21\]
+ VGND VGND VPWR VPWR _07802_ sky130_fd_sc_hd__o22a_1
XFILLER_0_142_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_220_Right_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21491_ rvcpu.dp.rf.reg_file_arr\[24\]\[6\] rvcpu.dp.rf.reg_file_arr\[25\]\[6\] rvcpu.dp.rf.reg_file_arr\[26\]\[6\]
+ rvcpu.dp.rf.reg_file_arr\[27\]\[6\] _08517_ _08519_ VGND VGND VPWR VPWR _08747_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_211_5555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30689_ clknet_leaf_261_clk _02424_ VGND VGND VPWR VPWR datamem.data_ram\[4\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_211_5566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32428_ clknet_leaf_253_clk _03850_ VGND VGND VPWR VPWR datamem.data_ram\[28\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_20442_ datamem.data_ram\[27\]\[12\] _06634_ _07730_ _07733_ VGND VGND VPWR VPWR
+ _07734_ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_338 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload340 clknet_1_0__leaf__10128_ VGND VGND VPWR VPWR clkload340/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_15_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20373_ datamem.data_ram\[46\]\[28\] _06625_ _06645_ datamem.data_ram\[40\]\[28\]
+ _07664_ VGND VGND VPWR VPWR _07665_ sky130_fd_sc_hd__o221a_1
X_32359_ clknet_leaf_275_clk _03781_ VGND VGND VPWR VPWR datamem.data_ram\[30\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload351 clknet_1_0__leaf__10090_ VGND VGND VPWR VPWR clkload351/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload70 clknet_leaf_68_clk VGND VGND VPWR VPWR clkload70/X sky130_fd_sc_hd__clkbuf_4
X_22112_ rvcpu.dp.plem.WriteDataM\[29\] _09221_ _09295_ rvcpu.dp.plem.WriteDataM\[13\]
+ _09320_ VGND VGND VPWR VPWR _09321_ sky130_fd_sc_hd__a221o_4
Xclkload81 clknet_leaf_39_clk VGND VGND VPWR VPWR clkload81/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_3_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload92 clknet_leaf_73_clk VGND VGND VPWR VPWR clkload92/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_100_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_208_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_208_clk
+ sky130_fd_sc_hd__clkbuf_8
X_26920_ _11837_ _11823_ VGND VGND VPWR VPWR _11838_ sky130_fd_sc_hd__and2_1
X_22043_ _09216_ _09262_ _09220_ VGND VGND VPWR VPWR _09265_ sky130_fd_sc_hd__a21o_4
Xhold2810 datamem.data_ram\[9\]\[27\] VGND VGND VPWR VPWR net3960 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26851_ _11781_ net1866 _11785_ _11793_ VGND VGND VPWR VPWR _03347_ sky130_fd_sc_hd__a31o_1
Xhold2821 datamem.data_ram\[5\]\[9\] VGND VGND VPWR VPWR net3971 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2832 datamem.data_ram\[56\]\[31\] VGND VGND VPWR VPWR net3982 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2843 datamem.data_ram\[20\]\[30\] VGND VGND VPWR VPWR net3993 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_162_4374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25802_ net1671 _11181_ _11177_ _11193_ VGND VGND VPWR VPWR _02898_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_162_4385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2854 datamem.data_ram\[42\]\[19\] VGND VGND VPWR VPWR net4004 sky130_fd_sc_hd__dlygate4sd3_1
X_23808__392 clknet_1_0__leaf__10206_ VGND VGND VPWR VPWR net518 sky130_fd_sc_hd__inv_2
XFILLER_0_227_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29570_ net924 _01305_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[26\]\[5\] sky130_fd_sc_hd__dfxtp_1
Xhold2865 rvcpu.dp.rf.reg_file_arr\[29\]\[2\] VGND VGND VPWR VPWR net4015 sky130_fd_sc_hd__dlygate4sd3_1
X_26782_ _11752_ VGND VGND VPWR VPWR _11753_ sky130_fd_sc_hd__clkbuf_4
Xhold2876 datamem.data_ram\[32\]\[24\] VGND VGND VPWR VPWR net4026 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2887 rvcpu.dp.rf.reg_file_arr\[22\]\[10\] VGND VGND VPWR VPWR net4037 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2898 rvcpu.dp.rf.reg_file_arr\[27\]\[26\] VGND VGND VPWR VPWR net4048 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_214_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28521_ _09290_ VGND VGND VPWR VPWR _12749_ sky130_fd_sc_hd__clkbuf_2
X_25733_ _11140_ VGND VGND VPWR VPWR _02882_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22945_ _10072_ VGND VGND VPWR VPWR _10073_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_74_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_175_4702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28452_ _12437_ net3142 _12704_ VGND VGND VPWR VPWR _12708_ sky130_fd_sc_hd__mux2_1
X_25664_ _11085_ net1928 _11097_ _11100_ VGND VGND VPWR VPWR _02853_ sky130_fd_sc_hd__a31o_1
X_22876_ _09516_ _10009_ _10011_ _09523_ VGND VGND VPWR VPWR _10012_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_65_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27403_ _12121_ VGND VGND VPWR VPWR _03571_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_121_3392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24615_ _10480_ net1970 _10502_ VGND VGND VPWR VPWR _10510_ sky130_fd_sc_hd__mux2_1
X_21827_ rvcpu.dp.rf.reg_file_arr\[12\]\[23\] rvcpu.dp.rf.reg_file_arr\[13\]\[23\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[23\] rvcpu.dp.rf.reg_file_arr\[15\]\[23\] _08578_
+ _08684_ VGND VGND VPWR VPWR _09066_ sky130_fd_sc_hd__mux4_1
X_28383_ _12371_ net3584 _12659_ VGND VGND VPWR VPWR _12667_ sky130_fd_sc_hd__mux2_1
X_25595_ _11047_ _11055_ VGND VGND VPWR VPWR _11061_ sky130_fd_sc_hd__and2_1
XFILLER_0_195_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27334_ _10598_ _11123_ _11713_ VGND VGND VPWR VPWR _12081_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_164_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24546_ _09309_ VGND VGND VPWR VPWR _10470_ sky130_fd_sc_hd__buf_2
XFILLER_0_109_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21758_ _08695_ _09000_ VGND VGND VPWR VPWR _09001_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20709_ datamem.data_ram\[26\]\[5\] _06932_ _06969_ datamem.data_ram\[29\]\[5\] VGND
+ VGND VPWR VPWR _08000_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_134_3720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27265_ _10811_ net3671 _12043_ VGND VGND VPWR VPWR _12044_ sky130_fd_sc_hd__mux2_1
X_24477_ _10428_ VGND VGND VPWR VPWR _02338_ sky130_fd_sc_hd__clkbuf_1
Xwire113 net34 VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__buf_1
X_21689_ rvcpu.dp.rf.reg_file_arr\[16\]\[16\] rvcpu.dp.rf.reg_file_arr\[17\]\[16\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[16\] rvcpu.dp.rf.reg_file_arr\[19\]\[16\] _08703_
+ _08721_ VGND VGND VPWR VPWR _08935_ sky130_fd_sc_hd__mux4_1
XFILLER_0_80_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29004_ _10060_ _13010_ VGND VGND VPWR VPWR _13013_ sky130_fd_sc_hd__and2_1
XFILLER_0_163_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_202_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26216_ net1315 _11436_ _11444_ VGND VGND VPWR VPWR _11446_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_24_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27196_ _12006_ VGND VGND VPWR VPWR _12007_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_130_3606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_3617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26147_ net1849 _11408_ VGND VGND VPWR VPWR _11410_ sky130_fd_sc_hd__and2_1
XFILLER_0_132_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26078_ _11370_ VGND VGND VPWR VPWR _02996_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_91_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29906_ clknet_leaf_142_clk _01641_ VGND VGND VPWR VPWR datamem.data_ram\[59\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_17920_ _05252_ VGND VGND VPWR VPWR _05293_ sky130_fd_sc_hd__clkbuf_4
X_25029_ _10739_ net1969 _10725_ VGND VGND VPWR VPWR _10740_ sky130_fd_sc_hd__mux2_1
X_17851_ rvcpu.dp.plem.ALUResultM\[11\] _05228_ _05176_ VGND VGND VPWR VPWR _05229_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_3557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29837_ net215 _01572_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[18\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_128_3568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_218_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_3579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16802_ _04647_ VGND VGND VPWR VPWR _04648_ sky130_fd_sc_hd__buf_4
XFILLER_0_218_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17782_ _05154_ VGND VGND VPWR VPWR _05179_ sky130_fd_sc_hd__buf_2
XFILLER_0_205_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14994_ _13358_ VGND VGND VPWR VPWR _13542_ sky130_fd_sc_hd__clkbuf_4
X_29768_ net1114 _01503_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[20\]\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_50_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16733_ _14089_ _14273_ VGND VGND VPWR VPWR _04611_ sky130_fd_sc_hd__nor2_2
X_19521_ datamem.data_ram\[58\]\[24\] _06803_ _06815_ datamem.data_ram\[61\]\[24\]
+ _06816_ VGND VGND VPWR VPWR _06817_ sky130_fd_sc_hd__o221a_1
X_26505__57 clknet_1_1__leaf__11602_ VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__inv_2
X_28719_ _12858_ VGND VGND VPWR VPWR _04150_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_50_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29699_ net1045 _01434_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[23\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19452_ datamem.data_ram\[43\]\[16\] _06739_ _06740_ _06747_ VGND VGND VPWR VPWR
+ _06748_ sky130_fd_sc_hd__o211a_1
X_31730_ net179 _03188_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[9\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_199_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16664_ _04574_ VGND VGND VPWR VPWR _01708_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_186_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18403_ _05766_ VGND VGND VPWR VPWR _05767_ sky130_fd_sc_hd__inv_2
X_15615_ net2273 _13248_ _14114_ VGND VGND VPWR VPWR _14116_ sky130_fd_sc_hd__mux2_1
X_31661_ clknet_leaf_71_clk net1257 VGND VGND VPWR VPWR rvcpu.dp.plmw.ALUResultW\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19383_ _06678_ VGND VGND VPWR VPWR _06679_ sky130_fd_sc_hd__buf_8
XFILLER_0_158_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16595_ _04537_ VGND VGND VPWR VPWR _01748_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18334_ _05456_ _05463_ _05469_ _05475_ _05666_ _05671_ VGND VGND VPWR VPWR _05699_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30612_ clknet_leaf_199_clk _02347_ VGND VGND VPWR VPWR datamem.data_ram\[52\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_15546_ _13638_ _14063_ _14069_ _14071_ VGND VGND VPWR VPWR _14072_ sky130_fd_sc_hd__and4_1
X_31592_ clknet_leaf_51_clk net1249 VGND VGND VPWR VPWR rvcpu.dp.plmw.PCPlus4W\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_189_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18265_ _05619_ _05620_ _05629_ VGND VGND VPWR VPWR _05630_ sky130_fd_sc_hd__a21o_1
X_30543_ clknet_leaf_147_clk _02278_ VGND VGND VPWR VPWR datamem.data_ram\[55\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15477_ _13308_ _13598_ _13600_ VGND VGND VPWR VPWR _14006_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_115_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17216_ _14135_ net2260 _04865_ VGND VGND VPWR VPWR _04868_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18196_ _05298_ _05556_ VGND VGND VPWR VPWR _05561_ sky130_fd_sc_hd__nor2_2
XFILLER_0_126_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30474_ net152 _02209_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[19\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32213_ clknet_leaf_250_clk _03635_ VGND VGND VPWR VPWR datamem.data_ram\[36\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17147_ _04831_ VGND VGND VPWR VPWR _01466_ sky130_fd_sc_hd__clkbuf_1
Xhold705 datamem.data_ram\[9\]\[7\] VGND VGND VPWR VPWR net1855 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold716 datamem.data_ram\[36\]\[6\] VGND VGND VPWR VPWR net1866 sky130_fd_sc_hd__dlygate4sd3_1
Xhold727 rvcpu.dp.pcreg.q\[23\] VGND VGND VPWR VPWR net1877 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold738 rvcpu.dp.rf.reg_file_arr\[6\]\[18\] VGND VGND VPWR VPWR net1888 sky130_fd_sc_hd__dlygate4sd3_1
X_32144_ clknet_leaf_278_clk _03566_ VGND VGND VPWR VPWR datamem.data_ram\[39\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_17078_ _14133_ net2875 _04793_ VGND VGND VPWR VPWR _04795_ sky130_fd_sc_hd__mux2_1
Xhold749 datamem.data_ram\[34\]\[30\] VGND VGND VPWR VPWR net1899 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16029_ _14354_ VGND VGND VPWR VPWR _02007_ sky130_fd_sc_hd__clkbuf_1
X_32075_ clknet_leaf_93_clk _03497_ VGND VGND VPWR VPWR datamem.data_ram\[33\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_24122__628 clknet_1_1__leaf__10260_ VGND VGND VPWR VPWR net754 sky130_fd_sc_hd__inv_2
Xhold2106 datamem.data_ram\[15\]\[17\] VGND VGND VPWR VPWR net3256 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31026_ clknet_leaf_58_clk _02761_ VGND VGND VPWR VPWR datamem.data_ram\[40\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2117 datamem.data_ram\[40\]\[30\] VGND VGND VPWR VPWR net3267 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2128 datamem.data_ram\[41\]\[21\] VGND VGND VPWR VPWR net3278 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2139 datamem.data_ram\[26\]\[25\] VGND VGND VPWR VPWR net3289 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1405 datamem.data_ram\[60\]\[14\] VGND VGND VPWR VPWR net2555 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_204_5381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1416 datamem.data_ram\[48\]\[14\] VGND VGND VPWR VPWR net2566 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1427 datamem.data_ram\[58\]\[27\] VGND VGND VPWR VPWR net2577 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_204_5392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1438 rvcpu.dp.rf.reg_file_arr\[11\]\[24\] VGND VGND VPWR VPWR net2588 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1449 rvcpu.dp.rf.reg_file_arr\[0\]\[8\] VGND VGND VPWR VPWR net2599 sky130_fd_sc_hd__dlygate4sd3_1
X_19719_ _06916_ _06996_ _07003_ _07014_ VGND VGND VPWR VPWR _07015_ sky130_fd_sc_hd__a31o_1
Xclkbuf_5_4__f_clk clknet_2_0_0_clk VGND VGND VPWR VPWR clknet_5_4__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_20991_ _08278_ _08279_ _06640_ VGND VGND VPWR VPWR _08280_ sky130_fd_sc_hd__mux2_1
XFILLER_0_224_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32977_ clknet_leaf_268_clk _04399_ VGND VGND VPWR VPWR datamem.data_ram\[63\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_200_5289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_196_5193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22730_ _09452_ _09871_ _09873_ _09457_ VGND VGND VPWR VPWR _09874_ sky130_fd_sc_hd__o211a_1
X_31928_ clknet_leaf_123_clk _03350_ VGND VGND VPWR VPWR datamem.data_ram\[60\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22661_ _09622_ _09806_ _09808_ VGND VGND VPWR VPWR _09809_ sky130_fd_sc_hd__a21o_1
X_31859_ clknet_leaf_124_clk _03313_ VGND VGND VPWR VPWR datamem.data_ram\[62\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_213_5606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_213_5617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24400_ _10379_ VGND VGND VPWR VPWR _02310_ sky130_fd_sc_hd__clkbuf_1
X_21612_ _08817_ _08860_ _08862_ _08700_ VGND VGND VPWR VPWR _08863_ sky130_fd_sc_hd__a211o_1
X_25380_ _10067_ _10936_ VGND VGND VPWR VPWR _10942_ sky130_fd_sc_hd__and2_1
X_22592_ rvcpu.dp.rf.reg_file_arr\[16\]\[15\] rvcpu.dp.rf.reg_file_arr\[17\]\[15\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[15\] rvcpu.dp.rf.reg_file_arr\[19\]\[15\] _09384_
+ _09430_ VGND VGND VPWR VPWR _09743_ sky130_fd_sc_hd__mux4_1
XFILLER_0_63_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24331_ _09244_ net4406 _10338_ VGND VGND VPWR VPWR _10342_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21543_ rvcpu.dp.rf.reg_file_arr\[16\]\[9\] rvcpu.dp.rf.reg_file_arr\[17\]\[9\] rvcpu.dp.rf.reg_file_arr\[18\]\[9\]
+ rvcpu.dp.rf.reg_file_arr\[19\]\[9\] _08524_ _08527_ VGND VGND VPWR VPWR _08796_
+ sky130_fd_sc_hd__mux4_2
X_22983__690 clknet_1_0__leaf__10083_ VGND VGND VPWR VPWR net816 sky130_fd_sc_hd__inv_2
XFILLER_0_30_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_209_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27050_ _11904_ net4368 _11910_ _11915_ VGND VGND VPWR VPWR _03424_ sky130_fd_sc_hd__a31o_1
XFILLER_0_145_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24262_ _10303_ VGND VGND VPWR VPWR _02248_ sky130_fd_sc_hd__clkbuf_1
X_21474_ _08511_ _08730_ VGND VGND VPWR VPWR _08731_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26001_ _11146_ VGND VGND VPWR VPWR _11325_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_105_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20425_ datamem.data_ram\[3\]\[12\] _06633_ _07243_ datamem.data_ram\[1\]\[12\] _06678_
+ VGND VGND VPWR VPWR _07717_ sky130_fd_sc_hd__o221a_1
XFILLER_0_15_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20356_ datamem.data_ram\[14\]\[28\] _06764_ _06700_ datamem.data_ram\[9\]\[28\]
+ VGND VGND VPWR VPWR _07648_ sky130_fd_sc_hd__o22a_1
Xclkload170 clknet_leaf_213_clk VGND VGND VPWR VPWR clkload170/X sky130_fd_sc_hd__clkbuf_4
Xclkload181 clknet_leaf_237_clk VGND VGND VPWR VPWR clkload181/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_144_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_164_4425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload192 clknet_leaf_226_clk VGND VGND VPWR VPWR clkload192/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_164_4436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27952_ _12428_ VGND VGND VPWR VPWR _03813_ sky130_fd_sc_hd__clkbuf_1
X_23075_ _10099_ VGND VGND VPWR VPWR _01265_ sky130_fd_sc_hd__clkbuf_1
X_20287_ datamem.data_ram\[21\]\[19\] _06865_ _06672_ datamem.data_ram\[23\]\[19\]
+ VGND VGND VPWR VPWR _07580_ sky130_fd_sc_hd__o22a_1
XFILLER_0_140_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26903_ _11813_ net1396 _11821_ _11826_ VGND VGND VPWR VPWR _03366_ sky130_fd_sc_hd__a31o_1
X_22026_ rvcpu.dp.plem.WriteDataM\[5\] _09215_ _09219_ _09250_ VGND VGND VPWR VPWR
+ _09251_ sky130_fd_sc_hd__a31o_4
X_24097__605 clknet_1_1__leaf__10258_ VGND VGND VPWR VPWR net731 sky130_fd_sc_hd__inv_2
XFILLER_0_101_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27883_ _12390_ VGND VGND VPWR VPWR _03782_ sky130_fd_sc_hd__clkbuf_1
Xhold10 rvcpu.dp.plde.PCPlus4E\[13\] VGND VGND VPWR VPWR net1160 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold21 rvcpu.dp.plem.PCPlus4M\[30\] VGND VGND VPWR VPWR net1171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 rvcpu.dp.plem.PCPlus4M\[14\] VGND VGND VPWR VPWR net1182 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2640 rvcpu.dp.rf.reg_file_arr\[14\]\[24\] VGND VGND VPWR VPWR net3790 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26834_ _11781_ net1656 _11773_ _11783_ VGND VGND VPWR VPWR _03340_ sky130_fd_sc_hd__a31o_1
XFILLER_0_179_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29622_ net976 _01357_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[25\]\[25\] sky130_fd_sc_hd__dfxtp_1
Xhold2651 datamem.data_ram\[27\]\[11\] VGND VGND VPWR VPWR net3801 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 rvcpu.dp.plde.PCPlus4E\[21\] VGND VGND VPWR VPWR net1193 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2662 datamem.data_ram\[31\]\[26\] VGND VGND VPWR VPWR net3812 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 rvcpu.dp.plde.PCPlus4E\[4\] VGND VGND VPWR VPWR net1204 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 rvcpu.dp.plem.lAuiPCM\[5\] VGND VGND VPWR VPWR net1215 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2673 datamem.data_ram\[4\]\[10\] VGND VGND VPWR VPWR net3823 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_67_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold76 rvcpu.dp.plde.PCPlus4E\[8\] VGND VGND VPWR VPWR net1226 sky130_fd_sc_hd__dlygate4sd3_1
X_23741__332 clknet_1_0__leaf__10199_ VGND VGND VPWR VPWR net458 sky130_fd_sc_hd__inv_2
Xhold2684 rvcpu.dp.rf.reg_file_arr\[23\]\[13\] VGND VGND VPWR VPWR net3834 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_67_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold87 rvcpu.dp.plde.PCPlus4E\[10\] VGND VGND VPWR VPWR net1237 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1950 datamem.data_ram\[30\]\[13\] VGND VGND VPWR VPWR net3100 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2695 datamem.data_ram\[19\]\[28\] VGND VGND VPWR VPWR net3845 sky130_fd_sc_hd__dlygate4sd3_1
X_29553_ net907 _01288_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[27\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_26765_ _11735_ net1779 _11737_ _11742_ VGND VGND VPWR VPWR _03312_ sky130_fd_sc_hd__a31o_1
Xhold1961 datamem.data_ram\[14\]\[18\] VGND VGND VPWR VPWR net3111 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_123_3443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold98 rvcpu.dp.plem.PCPlus4M\[11\] VGND VGND VPWR VPWR net1248 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_3454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1972 rvcpu.dp.rf.reg_file_arr\[11\]\[17\] VGND VGND VPWR VPWR net3122 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1983 datamem.data_ram\[7\]\[9\] VGND VGND VPWR VPWR net3133 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28504_ _12737_ net4365 net43 VGND VGND VPWR VPWR _12738_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1994 datamem.data_ram\[44\]\[17\] VGND VGND VPWR VPWR net3144 sky130_fd_sc_hd__dlygate4sd3_1
X_25716_ _11131_ VGND VGND VPWR VPWR _02874_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22928_ rvcpu.dp.plem.WriteDataM\[2\] VGND VGND VPWR VPWR _10060_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_1__f__10265_ clknet_0__10265_ VGND VGND VPWR VPWR clknet_1_1__leaf__10265_
+ sky130_fd_sc_hd__clkbuf_16
X_29484_ net846 _01219_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[2\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_26696_ _11700_ net1645 _11693_ _11702_ VGND VGND VPWR VPWR _03283_ sky130_fd_sc_hd__a31o_1
XFILLER_0_168_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28435_ _12697_ VGND VGND VPWR VPWR _04027_ sky130_fd_sc_hd__clkbuf_1
X_25647_ _11085_ net1387 _11077_ _11093_ VGND VGND VPWR VPWR _02843_ sky130_fd_sc_hd__a31o_1
XFILLER_0_39_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_211_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__10196_ clknet_0__10196_ VGND VGND VPWR VPWR clknet_1_1__leaf__10196_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_38_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22859_ rvcpu.dp.rf.reg_file_arr\[0\]\[29\] rvcpu.dp.rf.reg_file_arr\[1\]\[29\] rvcpu.dp.rf.reg_file_arr\[2\]\[29\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[29\] _09477_ _09383_ VGND VGND VPWR VPWR _09996_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_183_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15400_ _13932_ VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__inv_2
XFILLER_0_13_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16380_ net2108 _14478_ _14547_ VGND VGND VPWR VPWR _14555_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28366_ _12462_ net2742 net95 VGND VGND VPWR VPWR _12658_ sky130_fd_sc_hd__mux2_1
X_25578_ _10418_ _11042_ VGND VGND VPWR VPWR _11050_ sky130_fd_sc_hd__and2_1
XFILLER_0_186_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_183_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15331_ _13867_ _13639_ _13514_ VGND VGND VPWR VPWR _13868_ sky130_fd_sc_hd__o21ai_1
X_27317_ _12061_ net1465 _12065_ _12073_ VGND VGND VPWR VPWR _03533_ sky130_fd_sc_hd__a31o_1
XFILLER_0_171_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_183_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24529_ _10392_ net4300 _10456_ VGND VGND VPWR VPWR _10460_ sky130_fd_sc_hd__mux2_1
X_28297_ _12445_ net4001 _12613_ VGND VGND VPWR VPWR _12621_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_97_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18050_ _05418_ VGND VGND VPWR VPWR _05419_ sky130_fd_sc_hd__buf_2
X_15262_ _13420_ _13514_ _13800_ _13801_ _13503_ VGND VGND VPWR VPWR _13802_ sky130_fd_sc_hd__a32oi_2
X_27248_ _11976_ _12031_ VGND VGND VPWR VPWR _12038_ sky130_fd_sc_hd__and2_1
XFILLER_0_87_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17001_ net2138 _14484_ _04719_ VGND VGND VPWR VPWR _04753_ sky130_fd_sc_hd__mux2_1
XFILLER_0_227_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15193_ _13655_ _13733_ _13734_ _13735_ _13638_ VGND VGND VPWR VPWR _13736_ sky130_fd_sc_hd__o41a_1
X_27179_ _11991_ net1760 _11995_ _11997_ VGND VGND VPWR VPWR _03471_ sky130_fd_sc_hd__a31o_1
XFILLER_0_152_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_7 _05729_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23290__933 clknet_1_0__leaf__10131_ VGND VGND VPWR VPWR net1059 sky130_fd_sc_hd__inv_2
X_30190_ net544 _01925_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[8\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18952_ _05703_ _06284_ _06289_ VGND VGND VPWR VPWR _06290_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17903_ rvcpu.dp.plde.ALUSrcE VGND VGND VPWR VPWR _05276_ sky130_fd_sc_hd__inv_2
XFILLER_0_197_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18883_ _05473_ _05481_ _06194_ _05521_ VGND VGND VPWR VPWR _06225_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_52_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_206_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32900_ clknet_leaf_213_clk _04322_ VGND VGND VPWR VPWR datamem.data_ram\[0\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_283 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17834_ _13212_ rvcpu.dp.plde.RD2E\[21\] _05195_ VGND VGND VPWR VPWR _05217_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32831_ clknet_leaf_157_clk _04253_ VGND VGND VPWR VPWR datamem.data_ram\[12\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_14977_ _13446_ _13524_ VGND VGND VPWR VPWR _13525_ sky130_fd_sc_hd__or2_1
X_17765_ rvcpu.dp.plem.RdM\[4\] rvcpu.dp.plde.Rs2E\[4\] VGND VGND VPWR VPWR _05163_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_206_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19504_ datamem.data_ram\[53\]\[24\] _06723_ _06731_ datamem.data_ram\[51\]\[24\]
+ VGND VGND VPWR VPWR _06800_ sky130_fd_sc_hd__o22a_1
X_16716_ _04602_ VGND VGND VPWR VPWR _01684_ sky130_fd_sc_hd__clkbuf_1
X_32762_ clknet_leaf_274_clk _04184_ VGND VGND VPWR VPWR datamem.data_ram\[15\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_17696_ _05122_ VGND VGND VPWR VPWR _01192_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_198_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_190_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31713_ clknet_leaf_34_clk _03171_ VGND VGND VPWR VPWR rvcpu.dp.pcreg.q\[31\] sky130_fd_sc_hd__dfxtp_1
X_19435_ _06730_ VGND VGND VPWR VPWR _06731_ sky130_fd_sc_hd__buf_6
X_16647_ _14179_ net4322 _04562_ VGND VGND VPWR VPWR _04566_ sky130_fd_sc_hd__mux2_1
XFILLER_0_190_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32693_ clknet_leaf_287_clk _04115_ VGND VGND VPWR VPWR datamem.data_ram\[18\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_186_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31644_ clknet_leaf_28_clk net1156 VGND VGND VPWR VPWR rvcpu.dp.plmw.lAuiPCW\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_191_5090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16578_ _14179_ net4246 _04525_ VGND VGND VPWR VPWR _04529_ sky130_fd_sc_hd__mux2_1
X_19366_ _06661_ VGND VGND VPWR VPWR _06662_ sky130_fd_sc_hd__buf_6
XFILLER_0_45_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15529_ _13664_ _14054_ VGND VGND VPWR VPWR _14055_ sky130_fd_sc_hd__or2_1
X_18317_ _05681_ VGND VGND VPWR VPWR _05682_ sky130_fd_sc_hd__buf_2
XFILLER_0_57_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19297_ _06585_ rvcpu.dp.plem.ALUResultM\[7\] VGND VGND VPWR VPWR _06593_ sky130_fd_sc_hd__and2_1
X_31575_ clknet_leaf_71_clk datamem.rd_data_mem\[25\] VGND VGND VPWR VPWR rvcpu.dp.plmw.ReadDataW\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_178_Left_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18248_ _05311_ _05611_ _05612_ VGND VGND VPWR VPWR _05613_ sky130_fd_sc_hd__o21a_1
X_30526_ clknet_leaf_176_clk _02261_ VGND VGND VPWR VPWR datamem.data_ram\[56\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23911__468 clknet_1_1__leaf__10225_ VGND VGND VPWR VPWR net594 sky130_fd_sc_hd__inv_2
XFILLER_0_53_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18179_ rvcpu.dp.plem.ALUResultM\[26\] _05293_ _05294_ _13197_ VGND VGND VPWR VPWR
+ _05544_ sky130_fd_sc_hd__o22a_1
XFILLER_0_29_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30457_ net135 _02192_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[19\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold502 rvcpu.dp.plfd.InstrD\[8\] VGND VGND VPWR VPWR net1652 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold513 datamem.data_ram\[11\]\[3\] VGND VGND VPWR VPWR net1663 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20210_ _06752_ _07497_ _07502_ _06712_ VGND VGND VPWR VPWR _07503_ sky130_fd_sc_hd__o31a_1
Xhold524 datamem.data_ram\[49\]\[3\] VGND VGND VPWR VPWR net1674 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21190_ _08475_ VGND VGND VPWR VPWR _04446_ sky130_fd_sc_hd__clkbuf_1
Xhold535 datamem.data_ram\[1\]\[0\] VGND VGND VPWR VPWR net1685 sky130_fd_sc_hd__dlygate4sd3_1
X_30388_ clknet_leaf_175_clk _02123_ VGND VGND VPWR VPWR datamem.data_ram\[58\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_23610__229 clknet_1_0__leaf__10179_ VGND VGND VPWR VPWR net355 sky130_fd_sc_hd__inv_2
Xhold546 datamem.data_ram\[35\]\[4\] VGND VGND VPWR VPWR net1696 sky130_fd_sc_hd__dlygate4sd3_1
Xhold557 datamem.data_ram\[36\]\[0\] VGND VGND VPWR VPWR net1707 sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 datamem.data_ram\[15\]\[2\] VGND VGND VPWR VPWR net1718 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20141_ datamem.data_ram\[47\]\[27\] _06704_ _06617_ datamem.data_ram\[44\]\[27\]
+ _07433_ VGND VGND VPWR VPWR _07434_ sky130_fd_sc_hd__o221a_1
X_32127_ clknet_leaf_193_clk _03549_ VGND VGND VPWR VPWR datamem.data_ram\[7\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_206_5432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold579 datamem.data_ram\[49\]\[5\] VGND VGND VPWR VPWR net1729 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_206_5443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32058_ clknet_leaf_118_clk _03480_ VGND VGND VPWR VPWR datamem.data_ram\[48\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_20072_ _07154_ _07338_ _07343_ _07365_ _06860_ VGND VGND VPWR VPWR _07366_ sky130_fd_sc_hd__o32a_1
XPHY_EDGE_ROW_187_Left_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31009_ clknet_leaf_164_clk _02744_ VGND VGND VPWR VPWR datamem.data_ram\[11\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1202 datamem.data_ram\[2\]\[25\] VGND VGND VPWR VPWR net2352 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_198_5244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1213 rvcpu.dp.rf.reg_file_arr\[10\]\[1\] VGND VGND VPWR VPWR net2363 sky130_fd_sc_hd__dlygate4sd3_1
X_24880_ _10656_ VGND VGND VPWR VPWR _02513_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_198_5255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1224 rvcpu.dp.rf.reg_file_arr\[12\]\[9\] VGND VGND VPWR VPWR net2374 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1235 datamem.data_ram\[30\]\[16\] VGND VGND VPWR VPWR net2385 sky130_fd_sc_hd__dlygate4sd3_1
X_23267__913 clknet_1_1__leaf__10128_ VGND VGND VPWR VPWR net1039 sky130_fd_sc_hd__inv_2
Xhold1246 rvcpu.dp.rf.reg_file_arr\[23\]\[23\] VGND VGND VPWR VPWR net2396 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1257 datamem.data_ram\[35\]\[17\] VGND VGND VPWR VPWR net2407 sky130_fd_sc_hd__dlygate4sd3_1
X_23831_ _09306_ net2584 _10210_ VGND VGND VPWR VPWR _10212_ sky130_fd_sc_hd__mux2_1
XFILLER_0_212_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1268 datamem.data_ram\[31\]\[15\] VGND VGND VPWR VPWR net2418 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1279 rvcpu.dp.rf.reg_file_arr\[5\]\[0\] VGND VGND VPWR VPWR net2429 sky130_fd_sc_hd__dlygate4sd3_1
X_26550_ _11618_ net1352 _11608_ _11619_ VGND VGND VPWR VPWR _03220_ sky130_fd_sc_hd__a31o_1
XFILLER_0_68_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_408 _06645_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_196_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_419 _06754_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20974_ datamem.data_ram\[42\]\[15\] datamem.data_ram\[43\]\[15\] _06652_ VGND VGND
+ VPWR VPWR _08263_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25501_ _11005_ VGND VGND VPWR VPWR _02785_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_177_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22713_ _09441_ _09857_ VGND VGND VPWR VPWR _09858_ sky130_fd_sc_hd__nor2_1
X_26481_ _11524_ rvcpu.ALUResultE\[31\] _11289_ VGND VGND VPWR VPWR _11600_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_193_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_4262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_4273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28220_ _12365_ net3052 net45 VGND VGND VPWR VPWR _12579_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25432_ _10972_ VGND VGND VPWR VPWR _02749_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__10081_ _10081_ VGND VGND VPWR VPWR clknet_0__10081_ sky130_fd_sc_hd__clkbuf_16
X_22644_ rvcpu.dp.rf.reg_file_arr\[12\]\[17\] rvcpu.dp.rf.reg_file_arr\[13\]\[17\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[17\] rvcpu.dp.rf.reg_file_arr\[15\]\[17\] _09552_
+ _09721_ VGND VGND VPWR VPWR _09793_ sky130_fd_sc_hd__mux4_1
XFILLER_0_94_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_196_Left_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_153_4159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28151_ _12456_ net2638 net73 VGND VGND VPWR VPWR _12542_ sky130_fd_sc_hd__mux2_1
X_25363_ _10876_ net1389 _10920_ _10930_ VGND VGND VPWR VPWR _02722_ sky130_fd_sc_hd__a31o_1
X_22575_ rvcpu.dp.rf.reg_file_arr\[20\]\[14\] rvcpu.dp.rf.reg_file_arr\[21\]\[14\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[14\] rvcpu.dp.rf.reg_file_arr\[23\]\[14\] _09434_
+ _09558_ VGND VGND VPWR VPWR _09727_ sky130_fd_sc_hd__mux4_1
XFILLER_0_35_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27102_ _11833_ _11941_ VGND VGND VPWR VPWR _11948_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24314_ _10332_ VGND VGND VPWR VPWR _02271_ sky130_fd_sc_hd__clkbuf_1
X_28082_ _12505_ VGND VGND VPWR VPWR _03866_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21526_ _08777_ _08779_ _08743_ VGND VGND VPWR VPWR _08780_ sky130_fd_sc_hd__mux2_2
X_25294_ _10756_ net2748 _10887_ VGND VGND VPWR VPWR _10890_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27033_ _11904_ net1614 _11897_ _11905_ VGND VGND VPWR VPWR _03417_ sky130_fd_sc_hd__a31o_1
XFILLER_0_146_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_116_3280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24245_ _09285_ net3360 _10288_ VGND VGND VPWR VPWR _10294_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_116_3291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21457_ _08542_ _08714_ VGND VGND VPWR VPWR _08715_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20408_ datamem.data_ram\[45\]\[12\] _06662_ _06633_ datamem.data_ram\[43\]\[12\]
+ _07699_ VGND VGND VPWR VPWR _07700_ sky130_fd_sc_hd__o221a_1
X_21388_ _08533_ VGND VGND VPWR VPWR _08649_ sky130_fd_sc_hd__buf_6
Xoutput11 net11 VGND VGND VPWR VPWR Instr[18] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_187_4981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput9 net9 VGND VGND VPWR VPWR Instr[16] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_187_4992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput22 net22 VGND VGND VPWR VPWR Instr[28] sky130_fd_sc_hd__buf_2
Xoutput33 net33 VGND VGND VPWR VPWR Instr[9] sky130_fd_sc_hd__buf_2
XFILLER_0_82_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20339_ _07131_ _07623_ _07625_ _07630_ VGND VGND VPWR VPWR _07631_ sky130_fd_sc_hd__o31a_1
X_23585__206 clknet_1_0__leaf__10177_ VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__inv_2
X_28984_ _13001_ VGND VGND VPWR VPWR _04272_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_222_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_183_4878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_4889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27935_ _12419_ VGND VGND VPWR VPWR _03805_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_125_3505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3160 rvcpu.dp.rf.reg_file_arr\[30\]\[11\] VGND VGND VPWR VPWR net4310 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14900_ _13430_ _13323_ VGND VGND VPWR VPWR _13451_ sky130_fd_sc_hd__nand2_4
Xhold3171 datamem.data_ram\[4\]\[21\] VGND VGND VPWR VPWR net4321 sky130_fd_sc_hd__dlygate4sd3_1
X_22009_ _09237_ VGND VGND VPWR VPWR _01061_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_216_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold3182 datamem.data_ram\[2\]\[19\] VGND VGND VPWR VPWR net4332 sky130_fd_sc_hd__dlygate4sd3_1
X_27866_ _12381_ VGND VGND VPWR VPWR _03774_ sky130_fd_sc_hd__clkbuf_1
X_15880_ _14271_ _14273_ VGND VGND VPWR VPWR _14274_ sky130_fd_sc_hd__nor2_2
XFILLER_0_216_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold3193 datamem.data_ram\[59\]\[17\] VGND VGND VPWR VPWR net4343 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2470 datamem.data_ram\[9\]\[30\] VGND VGND VPWR VPWR net3620 sky130_fd_sc_hd__dlygate4sd3_1
X_14831_ _13382_ _13383_ VGND VGND VPWR VPWR _13384_ sky130_fd_sc_hd__or2_1
X_29605_ net959 _01340_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[25\]\[8\] sky130_fd_sc_hd__dfxtp_1
Xhold2481 datamem.data_ram\[32\]\[25\] VGND VGND VPWR VPWR net3631 sky130_fd_sc_hd__dlygate4sd3_1
X_26817_ _10268_ _08066_ _11609_ VGND VGND VPWR VPWR _11774_ sky130_fd_sc_hd__and3_2
XFILLER_0_204_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27797_ _12340_ VGND VGND VPWR VPWR _03746_ sky130_fd_sc_hd__clkbuf_1
Xhold2492 datamem.data_ram\[15\]\[12\] VGND VGND VPWR VPWR net3642 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_153_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17550_ _05044_ VGND VGND VPWR VPWR _01268_ sky130_fd_sc_hd__clkbuf_1
Xhold1780 rvcpu.dp.rf.reg_file_arr\[25\]\[23\] VGND VGND VPWR VPWR net2930 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_86_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26748_ _11687_ _11726_ VGND VGND VPWR VPWR _11732_ sky130_fd_sc_hd__and2_1
X_14762_ _13312_ _13314_ VGND VGND VPWR VPWR _13315_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_142_3896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29536_ net890 _01271_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[27\]\[3\] sky130_fd_sc_hd__dfxtp_1
Xhold1791 datamem.data_ram\[56\]\[29\] VGND VGND VPWR VPWR net2941 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16501_ net2987 _14461_ _04478_ VGND VGND VPWR VPWR _04488_ sky130_fd_sc_hd__mux2_1
X_17481_ _14195_ net2398 _04973_ VGND VGND VPWR VPWR _05008_ sky130_fd_sc_hd__mux2_1
X_29467_ net829 _01202_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[2\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26679_ _07191_ _10946_ _11494_ VGND VGND VPWR VPWR _11692_ sky130_fd_sc_hd__or3_1
XFILLER_0_196_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14693_ net3815 _13254_ _13245_ VGND VGND VPWR VPWR _13255_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1__f__10248_ clknet_0__10248_ VGND VGND VPWR VPWR clknet_1_1__leaf__10248_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_168_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19220_ rvcpu.dp.plde.ImmExtE\[26\] rvcpu.dp.plde.PCE\[26\] VGND VGND VPWR VPWR _06527_
+ sky130_fd_sc_hd__nand2_1
X_16432_ _14582_ VGND VGND VPWR VPWR _01824_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_183_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28418_ _12462_ net3643 _12678_ VGND VGND VPWR VPWR _12686_ sky130_fd_sc_hd__mux2_1
XFILLER_0_224_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29398_ clknet_leaf_1_clk _01133_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD2E\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_15_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__10179_ clknet_0__10179_ VGND VGND VPWR VPWR clknet_1_1__leaf__10179_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_39_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_184_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19151_ _06466_ _06460_ _06456_ VGND VGND VPWR VPWR _06467_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28349_ _12445_ net4392 _12641_ VGND VGND VPWR VPWR _12649_ sky130_fd_sc_hd__mux2_1
X_16363_ net4067 _14461_ _14536_ VGND VGND VPWR VPWR _14546_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18102_ rvcpu.dp.plde.ImmExtE\[21\] rvcpu.dp.SrcBFW_Mux.y\[21\] _05278_ VGND VGND
+ VPWR VPWR _05470_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15314_ _13850_ _13447_ _13309_ _13598_ _13509_ VGND VGND VPWR VPWR _13851_ sky130_fd_sc_hd__o32a_1
XFILLER_0_137_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19082_ rvcpu.dp.plde.ImmExtE\[9\] rvcpu.dp.plde.PCE\[9\] VGND VGND VPWR VPWR _06406_
+ sky130_fd_sc_hd__and2_1
X_31360_ clknet_leaf_22_clk _03063_ VGND VGND VPWR VPWR rvcpu.dp.plde.ImmExtE\[9\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_171_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16294_ _14509_ VGND VGND VPWR VPWR _01889_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_204_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18033_ _05402_ VGND VGND VPWR VPWR _05403_ sky130_fd_sc_hd__inv_2
X_30311_ net657 _02046_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[5\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_15245_ _13599_ _13379_ VGND VGND VPWR VPWR _13785_ sky130_fd_sc_hd__nand2_1
XFILLER_0_124_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31291_ clknet_leaf_18_clk _02994_ VGND VGND VPWR VPWR rvcpu.dp.plde.unsignE sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30242_ net596 _01977_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[7\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_15176_ _13717_ _13718_ _13374_ _13416_ VGND VGND VPWR VPWR _13719_ sky130_fd_sc_hd__a211o_1
XFILLER_0_22_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23748__338 clknet_1_0__leaf__10200_ VGND VGND VPWR VPWR net464 sky130_fd_sc_hd__inv_2
X_30173_ clknet_leaf_205_clk _01908_ VGND VGND VPWR VPWR datamem.data_ram\[58\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_19984_ datamem.data_ram\[11\]\[2\] _06942_ _06925_ datamem.data_ram\[15\]\[2\] VGND
+ VGND VPWR VPWR _07278_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18935_ _05776_ _05829_ _05531_ _05727_ VGND VGND VPWR VPWR _06274_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_197_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18866_ _05240_ _06195_ _06209_ VGND VGND VPWR VPWR rvcpu.ALUResultE\[20\] sky130_fd_sc_hd__a21o_1
XFILLER_0_20_1046 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17817_ rvcpu.dp.plem.ALUResultM\[27\] _05205_ _05178_ VGND VGND VPWR VPWR _05206_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18797_ _05781_ _06007_ _05819_ VGND VGND VPWR VPWR _06145_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_222_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32814_ clknet_leaf_283_clk _04236_ VGND VGND VPWR VPWR datamem.data_ram\[13\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_193_5130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17748_ _05149_ VGND VGND VPWR VPWR _01167_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_221_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32745_ clknet_leaf_234_clk _04167_ VGND VGND VPWR VPWR datamem.data_ram\[15\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17679_ net3242 _13268_ _05104_ VGND VGND VPWR VPWR _05113_ sky130_fd_sc_hd__mux2_1
XFILLER_0_193_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19418_ _06592_ VGND VGND VPWR VPWR _06714_ sky130_fd_sc_hd__buf_8
X_20690_ datamem.data_ram\[58\]\[5\] _07000_ _07138_ datamem.data_ram\[56\]\[5\] VGND
+ VGND VPWR VPWR _07981_ sky130_fd_sc_hd__a22o_1
XFILLER_0_186_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32676_ clknet_leaf_244_clk _04098_ VGND VGND VPWR VPWR datamem.data_ram\[18\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31627_ clknet_leaf_64_clk net1170 VGND VGND VPWR VPWR rvcpu.dp.plmw.lAuiPCW\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_19349_ _06644_ VGND VGND VPWR VPWR _06645_ sky130_fd_sc_hd__buf_8
XFILLER_0_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23297__939 clknet_1_0__leaf__10132_ VGND VGND VPWR VPWR net1065 sky130_fd_sc_hd__inv_2
XFILLER_0_150_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22360_ _09404_ VGND VGND VPWR VPWR _09523_ sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_198_Right_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31558_ clknet_leaf_71_clk datamem.rd_data_mem\[8\] VGND VGND VPWR VPWR rvcpu.dp.plmw.ReadDataW\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21311_ rvcpu.dp.rf.reg_file_arr\[0\]\[0\] rvcpu.dp.rf.reg_file_arr\[1\]\[0\] rvcpu.dp.rf.reg_file_arr\[2\]\[0\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[0\] _08566_ _08569_ VGND VGND VPWR VPWR _08573_ sky130_fd_sc_hd__mux4_1
X_30509_ clknet_leaf_218_clk _02244_ VGND VGND VPWR VPWR datamem.data_ram\[56\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22291_ rvcpu.dp.rf.reg_file_arr\[24\]\[1\] rvcpu.dp.rf.reg_file_arr\[25\]\[1\] rvcpu.dp.rf.reg_file_arr\[26\]\[1\]
+ rvcpu.dp.rf.reg_file_arr\[27\]\[1\] _09385_ _09431_ VGND VGND VPWR VPWR _09456_
+ sky130_fd_sc_hd__mux4_1
X_31489_ clknet_leaf_48_clk rvcpu.dp.lAuiPCE\[15\] VGND VGND VPWR VPWR rvcpu.dp.plem.lAuiPCM\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_24128__634 clknet_1_1__leaf__10260_ VGND VGND VPWR VPWR net760 sky130_fd_sc_hd__inv_2
XFILLER_0_103_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21242_ datamem.data_ram\[52\]\[17\] datamem.data_ram\[52\]\[9\] VGND VGND VPWR VPWR
+ _08505_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold310 datamem.data_ram\[21\]\[1\] VGND VGND VPWR VPWR net1460 sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 datamem.data_ram\[60\]\[5\] VGND VGND VPWR VPWR net1471 sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 datamem.data_ram\[58\]\[7\] VGND VGND VPWR VPWR net1482 sky130_fd_sc_hd__dlygate4sd3_1
Xhold343 datamem.data_ram\[37\]\[4\] VGND VGND VPWR VPWR net1493 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold354 datamem.data_ram\[59\]\[2\] VGND VGND VPWR VPWR net1504 sky130_fd_sc_hd__dlygate4sd3_1
X_21173_ _08449_ _08453_ _08461_ _06594_ VGND VGND VPWR VPWR _08462_ sky130_fd_sc_hd__a211o_1
Xhold365 datamem.data_ram\[12\]\[0\] VGND VGND VPWR VPWR net1515 sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 datamem.data_ram\[24\]\[3\] VGND VGND VPWR VPWR net1526 sky130_fd_sc_hd__dlygate4sd3_1
Xhold387 datamem.data_ram\[0\]\[1\] VGND VGND VPWR VPWR net1537 sky130_fd_sc_hd__dlygate4sd3_1
Xhold398 datamem.data_ram\[18\]\[4\] VGND VGND VPWR VPWR net1548 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__10199_ clknet_0__10199_ VGND VGND VPWR VPWR clknet_1_0__leaf__10199_
+ sky130_fd_sc_hd__clkbuf_16
X_20124_ datamem.data_ram\[6\]\[27\] _06719_ _06754_ datamem.data_ram\[2\]\[27\] VGND
+ VGND VPWR VPWR _07417_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_225_5885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25981_ net5 _11289_ VGND VGND VPWR VPWR _11314_ sky130_fd_sc_hd__or2_1
XFILLER_0_229_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_225_5896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27720_ _12080_ net4026 net49 VGND VGND VPWR VPWR _12299_ sky130_fd_sc_hd__mux2_1
X_24932_ _10684_ VGND VGND VPWR VPWR _02537_ sky130_fd_sc_hd__clkbuf_1
X_20055_ datamem.data_ram\[43\]\[26\] _06631_ _06684_ datamem.data_ram\[44\]\[26\]
+ VGND VGND VPWR VPWR _07349_ sky130_fd_sc_hd__o22a_1
Xhold1010 rvcpu.dp.rf.reg_file_arr\[7\]\[19\] VGND VGND VPWR VPWR net2160 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1021 rvcpu.dp.pcreg.q\[12\] VGND VGND VPWR VPWR net2171 sky130_fd_sc_hd__dlygate4sd3_1
X_27651_ _12142_ net3697 net79 VGND VGND VPWR VPWR _12262_ sky130_fd_sc_hd__mux2_1
Xhold1032 rvcpu.dp.rf.reg_file_arr\[10\]\[22\] VGND VGND VPWR VPWR net2182 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1043 rvcpu.dp.rf.reg_file_arr\[11\]\[31\] VGND VGND VPWR VPWR net2193 sky130_fd_sc_hd__dlygate4sd3_1
X_24863_ _10647_ VGND VGND VPWR VPWR _02505_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_175_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1054 datamem.data_ram\[1\]\[15\] VGND VGND VPWR VPWR net2204 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_159_4302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1065 datamem.data_ram\[61\]\[9\] VGND VGND VPWR VPWR net2215 sky130_fd_sc_hd__dlygate4sd3_1
X_26602_ _11618_ net1820 _11639_ _11648_ VGND VGND VPWR VPWR _03243_ sky130_fd_sc_hd__a31o_1
XFILLER_0_169_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_159_4313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1076 rvcpu.dp.rf.reg_file_arr\[19\]\[26\] VGND VGND VPWR VPWR net2226 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27582_ _12125_ net3740 _12224_ VGND VGND VPWR VPWR _12225_ sky130_fd_sc_hd__mux2_1
Xhold1087 datamem.data_ram\[23\]\[18\] VGND VGND VPWR VPWR net2237 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1098 datamem.data_ram\[28\]\[23\] VGND VGND VPWR VPWR net2248 sky130_fd_sc_hd__dlygate4sd3_1
X_24794_ _10609_ VGND VGND VPWR VPWR _02474_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_205 _09560_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_216 _09777_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_0__10202_ _10202_ VGND VGND VPWR VPWR clknet_0__10202_ sky130_fd_sc_hd__clkbuf_16
XANTENNA_227 _10072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29321_ clknet_leaf_12_clk _01056_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD1E\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26533_ _10209_ _11054_ _11609_ VGND VGND VPWR VPWR _11610_ sky130_fd_sc_hd__and3_1
Xclkbuf_1_1__f__10102_ clknet_0__10102_ VGND VGND VPWR VPWR clknet_1_1__leaf__10102_
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_238 _10780_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_212_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20957_ _08243_ _08244_ _08245_ _07819_ _06641_ VGND VGND VPWR VPWR _08246_ sky130_fd_sc_hd__a221o_1
XANTENNA_249 _13190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0__10133_ _10133_ VGND VGND VPWR VPWR clknet_0__10133_ sky130_fd_sc_hd__clkbuf_16
X_29252_ _13146_ VGND VGND VPWR VPWR _04395_ sky130_fd_sc_hd__clkbuf_1
X_26464_ _11576_ _11231_ _11540_ _06531_ _11587_ VGND VGND VPWR VPWR _11588_ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20888_ datamem.data_ram\[58\]\[14\] _06804_ _06790_ datamem.data_ram\[57\]\[14\]
+ _08177_ VGND VGND VPWR VPWR _08178_ sky130_fd_sc_hd__o221a_1
X_28203_ _12569_ VGND VGND VPWR VPWR _03923_ sky130_fd_sc_hd__clkbuf_1
X_25415_ _10963_ VGND VGND VPWR VPWR _02741_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29183_ _09251_ net3500 net63 VGND VGND VPWR VPWR _13109_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_118_3320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22627_ _09705_ _09768_ _09772_ _09776_ VGND VGND VPWR VPWR _09777_ sky130_fd_sc_hd__and4_1
X_26395_ _11521_ VGND VGND VPWR VPWR _11539_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_118_3331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28134_ _12439_ net3254 _12528_ VGND VGND VPWR VPWR _12533_ sky130_fd_sc_hd__mux2_1
X_25346_ _10919_ VGND VGND VPWR VPWR _10920_ sky130_fd_sc_hd__buf_2
XFILLER_0_180_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22558_ rvcpu.dp.rf.reg_file_arr\[28\]\[13\] rvcpu.dp.rf.reg_file_arr\[30\]\[13\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[13\] rvcpu.dp.rf.reg_file_arr\[31\]\[13\] _09400_
+ _09484_ VGND VGND VPWR VPWR _09711_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_165_Right_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28065_ _12496_ VGND VGND VPWR VPWR _03858_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_40_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21509_ _08725_ _08763_ VGND VGND VPWR VPWR _08764_ sky130_fd_sc_hd__nor2_1
XFILLER_0_224_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25277_ _10729_ net2521 _10878_ VGND VGND VPWR VPWR _10881_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_79_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22489_ _09469_ _09645_ VGND VGND VPWR VPWR _09646_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_79_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15030_ _13322_ _13492_ VGND VGND VPWR VPWR _13577_ sky130_fd_sc_hd__or2_1
X_27016_ _11889_ net1596 _11885_ _11894_ VGND VGND VPWR VPWR _03411_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_185_4929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24228_ _09252_ net3269 _10279_ VGND VGND VPWR VPWR _10285_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28967_ _10060_ _12989_ VGND VGND VPWR VPWR _12992_ sky130_fd_sc_hd__and2_1
X_16981_ net1926 _14463_ _04742_ VGND VGND VPWR VPWR _04743_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_88_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18720_ _05925_ _05697_ _05837_ VGND VGND VPWR VPWR _06072_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_88_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27918_ _12410_ VGND VGND VPWR VPWR _03797_ sky130_fd_sc_hd__clkbuf_1
X_15932_ net2052 _13257_ _14297_ VGND VGND VPWR VPWR _14302_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_144_3947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28898_ _12741_ net2974 net68 VGND VGND VPWR VPWR _12954_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_144_3958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18651_ _05915_ _06006_ _05705_ VGND VGND VPWR VPWR _06007_ sky130_fd_sc_hd__mux2_1
X_15863_ net2093 _13260_ _14258_ VGND VGND VPWR VPWR _14264_ sky130_fd_sc_hd__mux2_1
X_27849_ _12372_ VGND VGND VPWR VPWR _03766_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_189_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14814_ _13363_ _13364_ _13366_ VGND VGND VPWR VPWR _13367_ sky130_fd_sc_hd__a21oi_1
X_17602_ _05072_ VGND VGND VPWR VPWR _01236_ sky130_fd_sc_hd__clkbuf_1
X_30860_ clknet_leaf_154_clk _02595_ VGND VGND VPWR VPWR datamem.data_ram\[43\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18582_ _05705_ _05939_ _05940_ VGND VGND VPWR VPWR _05941_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_8_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15794_ _14183_ net3608 _14221_ VGND VGND VPWR VPWR _14227_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14745_ _13297_ VGND VGND VPWR VPWR _13298_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_203_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17533_ _13254_ net2370 _05032_ VGND VGND VPWR VPWR _05036_ sky130_fd_sc_hd__mux2_1
X_29519_ net881 _01254_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[28\]\[26\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_47_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30791_ clknet_leaf_264_clk _02526_ VGND VGND VPWR VPWR datamem.data_ram\[46\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_103_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17464_ _04999_ VGND VGND VPWR VPWR _01309_ sky130_fd_sc_hd__clkbuf_1
X_32530_ clknet_leaf_265_clk _03952_ VGND VGND VPWR VPWR datamem.data_ram\[23\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23181__852 clknet_1_1__leaf__10111_ VGND VGND VPWR VPWR net978 sky130_fd_sc_hd__inv_2
X_14676_ net2216 _13241_ _13214_ VGND VGND VPWR VPWR _13242_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19203_ _06512_ rvcpu.dp.plde.ImmExtE\[23\] _06493_ VGND VGND VPWR VPWR _06513_ sky130_fd_sc_hd__mux2_1
X_16415_ net2785 _14445_ _14572_ VGND VGND VPWR VPWR _14574_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_200_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17395_ _14177_ net3007 _04960_ VGND VGND VPWR VPWR _04963_ sky130_fd_sc_hd__mux2_1
X_32461_ clknet_leaf_231_clk _03883_ VGND VGND VPWR VPWR datamem.data_ram\[26\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19134_ _06441_ _06445_ VGND VGND VPWR VPWR _06452_ sky130_fd_sc_hd__nand2_1
X_31412_ clknet_leaf_22_clk _03115_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCE\[29\] sky130_fd_sc_hd__dfxtp_1
X_16346_ _14537_ VGND VGND VPWR VPWR _01865_ sky130_fd_sc_hd__clkbuf_1
X_32392_ clknet_leaf_182_clk _03814_ VGND VGND VPWR VPWR datamem.data_ram\[29\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_132_Right_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19065_ _06388_ _06391_ VGND VGND VPWR VPWR _06392_ sky130_fd_sc_hd__xnor2_2
X_31343_ clknet_leaf_17_clk _03046_ VGND VGND VPWR VPWR rvcpu.dp.plde.Rs1E\[4\] sky130_fd_sc_hd__dfxtp_1
X_23453__103 clknet_1_0__leaf__10156_ VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__inv_2
X_16277_ net2042 _14442_ _14500_ VGND VGND VPWR VPWR _14501_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15228_ _13682_ _13366_ _13526_ _13768_ _13521_ VGND VGND VPWR VPWR _13769_ sky130_fd_sc_hd__o311a_1
X_18016_ rvcpu.dp.plem.ALUResultM\[1\] VGND VGND VPWR VPWR _05386_ sky130_fd_sc_hd__inv_2
X_31274_ clknet_leaf_126_clk _02977_ VGND VGND VPWR VPWR datamem.data_ram\[24\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23982__517 clknet_1_0__leaf__10239_ VGND VGND VPWR VPWR net643 sky130_fd_sc_hd__inv_2
X_23533__160 clknet_1_0__leaf__10171_ VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__inv_2
XFILLER_0_140_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30225_ net579 _01960_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[7\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_15159_ _13305_ _13526_ VGND VGND VPWR VPWR _13703_ sky130_fd_sc_hd__or2_2
XFILLER_0_121_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_205_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30156_ net518 _01891_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[0\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_1035 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout119 _00000_ VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__dlymetal6s2s_1
X_19967_ datamem.data_ram\[11\]\[18\] _06737_ _06619_ datamem.data_ram\[12\]\[18\]
+ _07260_ VGND VGND VPWR VPWR _07261_ sky130_fd_sc_hd__o221a_1
XFILLER_0_201_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18918_ _05702_ _06010_ _06143_ _05990_ _06257_ VGND VGND VPWR VPWR _06258_ sky130_fd_sc_hd__o221a_1
X_30087_ net449 _01822_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[11\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19898_ datamem.data_ram\[7\]\[17\] _07020_ _06658_ datamem.data_ram\[1\]\[17\] VGND
+ VGND VPWR VPWR _07193_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_220_5771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18849_ _05655_ _06184_ _06190_ _06193_ VGND VGND VPWR VPWR rvcpu.ALUResultE\[19\]
+ sky130_fd_sc_hd__o211ai_2
XTAP_TAPCELL_ROW_220_5782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21860_ rvcpu.dp.rf.reg_file_arr\[28\]\[25\] rvcpu.dp.rf.reg_file_arr\[30\]\[25\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[25\] rvcpu.dp.rf.reg_file_arr\[31\]\[25\] _08568_
+ _08683_ VGND VGND VPWR VPWR _09097_ sky130_fd_sc_hd__mux4_1
XFILLER_0_77_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20811_ datamem.data_ram\[40\]\[30\] _06973_ _08096_ _07636_ _08100_ VGND VGND VPWR
+ VPWR _08101_ sky130_fd_sc_hd__a221o_1
XFILLER_0_222_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21791_ rvcpu.dp.rf.reg_file_arr\[8\]\[21\] rvcpu.dp.rf.reg_file_arr\[10\]\[21\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[21\] rvcpu.dp.rf.reg_file_arr\[11\]\[21\] _08560_
+ _08561_ VGND VGND VPWR VPWR _09032_ sky130_fd_sc_hd__mux4_1
X_30989_ clknet_leaf_59_clk _02724_ VGND VGND VPWR VPWR datamem.data_ram\[13\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20742_ datamem.data_ram\[47\]\[6\] _06623_ _06615_ datamem.data_ram\[45\]\[6\] _08031_
+ VGND VGND VPWR VPWR _08032_ sky130_fd_sc_hd__a221o_1
X_23305__946 clknet_1_0__leaf__10133_ VGND VGND VPWR VPWR net1072 sky130_fd_sc_hd__inv_2
X_32728_ clknet_leaf_181_clk _04150_ VGND VGND VPWR VPWR datamem.data_ram\[16\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_174_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23917__474 clknet_1_1__leaf__10225_ VGND VGND VPWR VPWR net600 sky130_fd_sc_hd__inv_2
XFILLER_0_190_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_150_4107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32659_ clknet_leaf_171_clk _04081_ VGND VGND VPWR VPWR datamem.data_ram\[19\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_20673_ _06596_ _07930_ _07941_ _07963_ VGND VGND VPWR VPWR _07964_ sky130_fd_sc_hd__a211oi_2
XTAP_TAPCELL_ROW_189_5029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25200_ _07122_ VGND VGND VPWR VPWR _10838_ sky130_fd_sc_hd__buf_8
XFILLER_0_163_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22412_ _09482_ _09572_ VGND VGND VPWR VPWR _09573_ sky130_fd_sc_hd__or2_1
X_26180_ _08570_ _11413_ VGND VGND VPWR VPWR _11427_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_171_4590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23392_ _09314_ net2401 _10143_ VGND VGND VPWR VPWR _10147_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25131_ _10797_ VGND VGND VPWR VPWR _02623_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22343_ rvcpu.dp.rf.reg_file_arr\[8\]\[2\] rvcpu.dp.rf.reg_file_arr\[10\]\[2\] rvcpu.dp.rf.reg_file_arr\[9\]\[2\]
+ rvcpu.dp.rf.reg_file_arr\[11\]\[2\] _09483_ _09485_ VGND VGND VPWR VPWR _09507_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_66_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25062_ _09247_ VGND VGND VPWR VPWR _10760_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_227_5936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22274_ _09389_ _09414_ _09428_ _09439_ VGND VGND VPWR VPWR _09440_ sky130_fd_sc_hd__and4_1
XFILLER_0_182_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_227_5947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_4036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold140 rvcpu.dp.plem.ALUResultM\[19\] VGND VGND VPWR VPWR net1290 sky130_fd_sc_hd__dlygate4sd3_1
X_21225_ _08468_ net36 _08489_ VGND VGND VPWR VPWR _04436_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_148_4047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold151 datamem.data_ram\[41\]\[7\] VGND VGND VPWR VPWR net1301 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_4058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29870_ net248 _01605_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[17\]\[1\] sky130_fd_sc_hd__dfxtp_1
Xhold162 datamem.data_ram\[43\]\[5\] VGND VGND VPWR VPWR net1312 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold173 datamem.data_ram\[42\]\[0\] VGND VGND VPWR VPWR net1323 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_180_4804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold184 datamem.data_ram\[41\]\[2\] VGND VGND VPWR VPWR net1334 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_180_4815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28821_ _12702_ net4304 _12905_ VGND VGND VPWR VPWR _12913_ sky130_fd_sc_hd__mux2_1
Xhold195 datamem.data_ram\[44\]\[4\] VGND VGND VPWR VPWR net1345 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_180_4826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21156_ _06922_ _08443_ _08444_ _07866_ VGND VGND VPWR VPWR _08445_ sky130_fd_sc_hd__o22a_1
X_23351__988 clknet_1_1__leaf__10137_ VGND VGND VPWR VPWR net1114 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_70_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20107_ datamem.data_ram\[16\]\[10\] _06696_ _06656_ datamem.data_ram\[17\]\[10\]
+ VGND VGND VPWR VPWR _07401_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_6_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21087_ _06605_ datamem.data_ram\[51\]\[7\] _07911_ datamem.data_ram\[50\]\[7\] _07636_
+ VGND VGND VPWR VPWR _08376_ sky130_fd_sc_hd__o221a_1
XFILLER_0_176_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25964_ rvcpu.dp.plfd.InstrD\[4\] _11155_ VGND VGND VPWR VPWR _11305_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_70_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28752_ _12749_ net4407 net41 VGND VGND VPWR VPWR _12876_ sky130_fd_sc_hd__mux2_1
XFILLER_0_176_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27703_ _12142_ net3635 _12289_ VGND VGND VPWR VPWR _12290_ sky130_fd_sc_hd__mux2_1
X_20038_ datamem.data_ram\[20\]\[26\] _06619_ _07330_ _07331_ VGND VGND VPWR VPWR
+ _07332_ sky130_fd_sc_hd__o211a_1
X_24915_ _10675_ VGND VGND VPWR VPWR _02529_ sky130_fd_sc_hd__clkbuf_1
X_25895_ _13682_ _11256_ _11258_ _11265_ VGND VGND VPWR VPWR _02919_ sky130_fd_sc_hd__o211a_1
X_28683_ _12839_ VGND VGND VPWR VPWR _04133_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_107_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24846_ _10452_ net2957 _10631_ VGND VGND VPWR VPWR _10638_ sky130_fd_sc_hd__mux2_1
X_27634_ _12252_ VGND VGND VPWR VPWR _03671_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_178_4766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_178_4777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27565_ _12080_ net3905 net82 VGND VGND VPWR VPWR _12216_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24777_ _08124_ _07858_ VGND VGND VPWR VPWR _10599_ sky130_fd_sc_hd__nand2_2
XFILLER_0_205_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21989_ _09218_ VGND VGND VPWR VPWR _09219_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_200_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29304_ clknet_leaf_0_clk _01039_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD1E\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27496_ _12178_ _12106_ _12168_ VGND VGND VPWR VPWR _12179_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_194_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23245__893 clknet_1_0__leaf__10126_ VGND VGND VPWR VPWR net1019 sky130_fd_sc_hd__inv_2
XFILLER_0_3_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26447_ _11145_ VGND VGND VPWR VPWR _11576_ sky130_fd_sc_hd__buf_2
XFILLER_0_139_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29235_ _13137_ VGND VGND VPWR VPWR _04387_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_42_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16200_ net3895 _14451_ _14443_ VGND VGND VPWR VPWR _14452_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_193_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29166_ _09251_ net3566 _13094_ VGND VGND VPWR VPWR _13100_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_3773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17180_ _04848_ VGND VGND VPWR VPWR _01450_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26378_ _11525_ VGND VGND VPWR VPWR _11526_ sky130_fd_sc_hd__buf_2
XFILLER_0_187_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_3784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_3795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28117_ _12365_ net3468 net74 VGND VGND VPWR VPWR _12524_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16131_ _14408_ VGND VGND VPWR VPWR _01959_ sky130_fd_sc_hd__clkbuf_1
X_25329_ _10910_ VGND VGND VPWR VPWR _02708_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29097_ _13063_ VGND VGND VPWR VPWR _04323_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28048_ _12487_ VGND VGND VPWR VPWR _03850_ sky130_fd_sc_hd__clkbuf_1
X_16062_ net2554 _13244_ _14371_ VGND VGND VPWR VPWR _14372_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_224_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15013_ _13303_ _13560_ VGND VGND VPWR VPWR _13561_ sky130_fd_sc_hd__and2_2
X_30010_ clknet_leaf_268_clk _01745_ VGND VGND VPWR VPWR datamem.data_ram\[59\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_19821_ datamem.data_ram\[31\]\[9\] _06672_ _07112_ _07115_ VGND VGND VPWR VPWR _07116_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_209_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29999_ net369 _01734_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[14\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_19752_ _06715_ _07041_ _07046_ VGND VGND VPWR VPWR _07047_ sky130_fd_sc_hd__or3_1
X_16964_ net2551 _14447_ _04731_ VGND VGND VPWR VPWR _04734_ sky130_fd_sc_hd__mux2_1
X_18703_ _05410_ _05607_ _06041_ VGND VGND VPWR VPWR _06056_ sky130_fd_sc_hd__nand3_1
X_15915_ net2430 _13232_ _14286_ VGND VGND VPWR VPWR _14293_ sky130_fd_sc_hd__mux2_1
XFILLER_0_223_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19683_ datamem.data_ram\[62\]\[0\] _06978_ _06926_ datamem.data_ram\[63\]\[0\] VGND
+ VGND VPWR VPWR _06979_ sky130_fd_sc_hd__a22o_1
X_31961_ clknet_leaf_122_clk _03383_ VGND VGND VPWR VPWR datamem.data_ram\[28\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16895_ _04697_ VGND VGND VPWR VPWR _01592_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_194_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18634_ _05363_ _05988_ _05989_ _05990_ VGND VGND VPWR VPWR _05991_ sky130_fd_sc_hd__o22a_1
X_30912_ clknet_leaf_260_clk _02647_ VGND VGND VPWR VPWR datamem.data_ram\[41\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_24157__660 clknet_1_0__leaf__10263_ VGND VGND VPWR VPWR net786 sky130_fd_sc_hd__inv_2
X_15846_ net1977 _13235_ _14247_ VGND VGND VPWR VPWR _14255_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31892_ clknet_leaf_108_clk _03346_ VGND VGND VPWR VPWR datamem.data_ram\[36\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23563__186 clknet_1_1__leaf__10175_ VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__inv_2
XFILLER_0_189_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_201_Right_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18565_ _05675_ _05759_ VGND VGND VPWR VPWR _05925_ sky130_fd_sc_hd__or2_2
X_30843_ clknet_leaf_173_clk _02578_ VGND VGND VPWR VPWR datamem.data_ram\[44\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15777_ _14166_ net3381 _14210_ VGND VGND VPWR VPWR _14218_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17516_ _13229_ net3879 _05021_ VGND VGND VPWR VPWR _05027_ sky130_fd_sc_hd__mux2_1
X_14728_ _13280_ VGND VGND VPWR VPWR _13281_ sky130_fd_sc_hd__buf_4
XFILLER_0_185_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18496_ _05782_ VGND VGND VPWR VPWR _05858_ sky130_fd_sc_hd__inv_2
X_30774_ clknet_leaf_221_clk _02509_ VGND VGND VPWR VPWR datamem.data_ram\[46\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_23027__729 clknet_1_1__leaf__10088_ VGND VGND VPWR VPWR net855 sky130_fd_sc_hd__inv_2
XFILLER_0_28_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32513_ clknet_leaf_77_clk _03935_ VGND VGND VPWR VPWR datamem.data_ram\[24\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_17447_ _04990_ VGND VGND VPWR VPWR _01317_ sky130_fd_sc_hd__clkbuf_1
X_14659_ _13228_ VGND VGND VPWR VPWR _13229_ sky130_fd_sc_hd__clkbuf_8
Xclkbuf_leaf_180_clk clknet_5_19__leaf_clk VGND VGND VPWR VPWR clknet_leaf_180_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_184_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32444_ clknet_leaf_80_clk _03866_ VGND VGND VPWR VPWR datamem.data_ram\[27\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17378_ _14160_ net4218 _04949_ VGND VGND VPWR VPWR _04954_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19117_ _06421_ _06429_ _06430_ _06427_ VGND VGND VPWR VPWR _06437_ sky130_fd_sc_hd__a31o_1
X_16329_ _14528_ VGND VGND VPWR VPWR _01873_ sky130_fd_sc_hd__clkbuf_1
X_32375_ clknet_leaf_277_clk _03797_ VGND VGND VPWR VPWR datamem.data_ram\[2\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19048_ _06375_ _06376_ VGND VGND VPWR VPWR _06377_ sky130_fd_sc_hd__xnor2_2
X_31326_ clknet_leaf_24_clk _03029_ VGND VGND VPWR VPWR rvcpu.dp.plde.funct3E\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_140_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31257_ clknet_leaf_15_clk _02960_ VGND VGND VPWR VPWR rvcpu.dp.plfd.InstrD\[15\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_26_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_929 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__10105_ clknet_0__10105_ VGND VGND VPWR VPWR clknet_1_0__leaf__10105_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21010_ _08298_ VGND VGND VPWR VPWR _08299_ sky130_fd_sc_hd__inv_2
X_30208_ net562 _01943_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[8\]\[27\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_222_5822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31188_ clknet_leaf_40_clk _02891_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCPlus4D\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_222_5833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30139_ net501 _01874_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[10\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_1006 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_214_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24700_ _10557_ VGND VGND VPWR VPWR _02432_ sky130_fd_sc_hd__clkbuf_1
X_21912_ _09144_ _09145_ _08540_ VGND VGND VPWR VPWR _09146_ sky130_fd_sc_hd__mux2_1
XFILLER_0_223_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25680_ _07808_ _11109_ _10044_ VGND VGND VPWR VPWR _11110_ sky130_fd_sc_hd__or3_1
X_22892_ rvcpu.dp.rf.reg_file_arr\[28\]\[31\] rvcpu.dp.rf.reg_file_arr\[30\]\[31\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[31\] rvcpu.dp.rf.reg_file_arr\[31\]\[31\] _09381_
+ _09423_ VGND VGND VPWR VPWR _10027_ sky130_fd_sc_hd__mux4_1
XFILLER_0_179_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24631_ _10518_ VGND VGND VPWR VPWR _02402_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21843_ _08542_ _09080_ _08513_ VGND VGND VPWR VPWR _09081_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_214_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27350_ _12091_ net4075 _12081_ VGND VGND VPWR VPWR _12092_ sky130_fd_sc_hd__mux2_1
X_24562_ _10480_ net3624 _10466_ VGND VGND VPWR VPWR _10481_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21774_ _08692_ _09013_ _09015_ VGND VGND VPWR VPWR _09016_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_173_4641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26301_ _11483_ VGND VGND VPWR VPWR _03107_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_173_4652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23513_ _09240_ net4337 _10162_ VGND VGND VPWR VPWR _10165_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20725_ _07822_ _08013_ _08014_ _07845_ VGND VGND VPWR VPWR _08015_ sky130_fd_sc_hd__o211a_1
X_27281_ _07791_ _08133_ _11839_ VGND VGND VPWR VPWR _12052_ sky130_fd_sc_hd__or3_1
XFILLER_0_148_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_171_clk clknet_5_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_171_clk
+ sky130_fd_sc_hd__clkbuf_8
X_24493_ _09326_ datamem.data_ram\[52\]\[30\] _10430_ VGND VGND VPWR VPWR _10437_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_191_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29020_ _12737_ net3458 net66 VGND VGND VPWR VPWR _13022_ sky130_fd_sc_hd__mux2_1
X_26232_ _11451_ _11454_ _11455_ _11456_ VGND VGND VPWR VPWR _03065_ sky130_fd_sc_hd__a211o_1
X_23850__414 clknet_1_1__leaf__10208_ VGND VGND VPWR VPWR net540 sky130_fd_sc_hd__inv_2
X_23444_ clknet_1_0__leaf__10152_ VGND VGND VPWR VPWR _10156_ sky130_fd_sc_hd__buf_1
XFILLER_0_11_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20656_ datamem.data_ram\[42\]\[29\] _06804_ _06837_ datamem.data_ram\[40\]\[29\]
+ VGND VGND VPWR VPWR _07947_ sky130_fd_sc_hd__o22a_1
XFILLER_0_68_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26163_ _11418_ VGND VGND VPWR VPWR _03034_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20587_ datamem.data_ram\[54\]\[13\] _06628_ _06706_ datamem.data_ram\[55\]\[13\]
+ _07877_ VGND VGND VPWR VPWR _07878_ sky130_fd_sc_hd__o221a_1
XFILLER_0_6_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25114_ _10788_ VGND VGND VPWR VPWR _02615_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22326_ _09389_ VGND VGND VPWR VPWR _09491_ sky130_fd_sc_hd__clkbuf_4
X_26094_ net2400 _11372_ VGND VGND VPWR VPWR _11382_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_132_3670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_72_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29922_ net292 _01657_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[16\]\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_72_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25045_ _10478_ net2377 _10742_ VGND VGND VPWR VPWR _10749_ sky130_fd_sc_hd__mux2_1
X_22257_ _09401_ VGND VGND VPWR VPWR _09423_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_197_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24026__557 clknet_1_1__leaf__10243_ VGND VGND VPWR VPWR net683 sky130_fd_sc_hd__inv_2
X_21208_ _08468_ VGND VGND VPWR VPWR _08487_ sky130_fd_sc_hd__buf_2
XFILLER_0_218_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29853_ net231 _01588_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[18\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22188_ _09366_ VGND VGND VPWR VPWR _01111_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_109_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_109_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28804_ _12749_ net2361 _12896_ VGND VGND VPWR VPWR _12904_ sky130_fd_sc_hd__mux2_1
XFILLER_0_218_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21139_ datamem.data_ram\[53\]\[23\] _06722_ _06765_ datamem.data_ram\[52\]\[23\]
+ _08427_ VGND VGND VPWR VPWR _08428_ sky130_fd_sc_hd__o221a_1
X_29784_ net1130 _01519_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[20\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26996_ _11882_ VGND VGND VPWR VPWR _03403_ sky130_fd_sc_hd__clkbuf_1
X_28735_ _12766_ net4152 _12859_ VGND VGND VPWR VPWR _12867_ sky130_fd_sc_hd__mux2_1
XFILLER_0_219_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25947_ net1929 _11290_ _11286_ _11295_ VGND VGND VPWR VPWR _02941_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_31_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15700_ _14170_ net2553 _14152_ VGND VGND VPWR VPWR _14171_ sky130_fd_sc_hd__mux2_1
X_16680_ _04583_ VGND VGND VPWR VPWR _01701_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_198_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25878_ _08620_ _08621_ _11254_ VGND VGND VPWR VPWR _11255_ sky130_fd_sc_hd__and3_1
X_28666_ _12830_ VGND VGND VPWR VPWR _04125_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24829_ _10628_ VGND VGND VPWR VPWR _02490_ sky130_fd_sc_hd__clkbuf_1
X_27617_ _12243_ VGND VGND VPWR VPWR _03663_ sky130_fd_sc_hd__clkbuf_1
X_15631_ net1966 _13272_ _14114_ VGND VGND VPWR VPWR _14124_ sky130_fd_sc_hd__mux2_1
X_28597_ _12793_ VGND VGND VPWR VPWR _04093_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_198_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_201_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15562_ _13441_ _14083_ _14084_ _13366_ _14085_ VGND VGND VPWR VPWR _14086_ sky130_fd_sc_hd__o221a_1
XFILLER_0_150_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18350_ _05713_ _05714_ _05671_ VGND VGND VPWR VPWR _05715_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_3824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27548_ _12142_ net3587 net98 VGND VGND VPWR VPWR _12207_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_139_3835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17301_ _04901_ VGND VGND VPWR VPWR _04913_ sky130_fd_sc_hd__buf_4
XFILLER_0_138_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_29_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15493_ _13682_ _14020_ _13599_ VGND VGND VPWR VPWR _14021_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_154_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27479_ _12125_ net2967 _12169_ VGND VGND VPWR VPWR _12170_ sky130_fd_sc_hd__mux2_1
X_18281_ _05642_ _05297_ _05645_ VGND VGND VPWR VPWR _05646_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_84_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_182_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_162_clk clknet_5_25__leaf_clk VGND VGND VPWR VPWR clknet_leaf_162_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_29_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29218_ _11533_ net1607 _13122_ _13128_ VGND VGND VPWR VPWR _04379_ sky130_fd_sc_hd__a31o_1
XFILLER_0_182_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17232_ _04864_ VGND VGND VPWR VPWR _04876_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_61_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30490_ clknet_leaf_205_clk _02225_ VGND VGND VPWR VPWR datamem.data_ram\[57\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17163_ _04839_ VGND VGND VPWR VPWR _01458_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29149_ _09284_ net4239 _13085_ VGND VGND VPWR VPWR _13091_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16114_ _14399_ VGND VGND VPWR VPWR _01967_ sky130_fd_sc_hd__clkbuf_1
X_32160_ clknet_leaf_162_clk _03582_ VGND VGND VPWR VPWR datamem.data_ram\[38\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17094_ _14149_ net4428 _04793_ VGND VGND VPWR VPWR _04803_ sky130_fd_sc_hd__mux2_1
Xhold909 rvcpu.dp.rf.reg_file_arr\[9\]\[9\] VGND VGND VPWR VPWR net2059 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31111_ clknet_leaf_61_clk _02846_ VGND VGND VPWR VPWR datamem.data_ram\[43\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_16045_ net1974 _13220_ _14360_ VGND VGND VPWR VPWR _14363_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32091_ clknet_leaf_213_clk _03513_ VGND VGND VPWR VPWR datamem.data_ram\[8\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31042_ clknet_leaf_98_clk _02777_ VGND VGND VPWR VPWR datamem.data_ram\[41\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19804_ datamem.data_ram\[14\]\[9\] _06764_ _06692_ datamem.data_ram\[10\]\[9\] VGND
+ VGND VPWR VPWR _07099_ sky130_fd_sc_hd__o22a_1
XFILLER_0_23_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17996_ _05363_ _05365_ VGND VGND VPWR VPWR _05366_ sky130_fd_sc_hd__nor2_1
XFILLER_0_208_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1609 datamem.data_ram\[61\]\[15\] VGND VGND VPWR VPWR net2759 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_193_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19735_ datamem.data_ram\[5\]\[25\] _06703_ _06707_ datamem.data_ram\[7\]\[25\] VGND
+ VGND VPWR VPWR _07030_ sky130_fd_sc_hd__o22a_1
XFILLER_0_193_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16947_ net2122 _14430_ _04720_ VGND VGND VPWR VPWR _04725_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_223_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31944_ clknet_leaf_115_clk _03366_ VGND VGND VPWR VPWR datamem.data_ram\[32\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_19666_ datamem.data_ram\[40\]\[0\] _06936_ _06954_ datamem.data_ram\[44\]\[0\] VGND
+ VGND VPWR VPWR _06962_ sky130_fd_sc_hd__a22o_1
X_16878_ _04688_ VGND VGND VPWR VPWR _01600_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18617_ _05354_ _05974_ _05784_ _05355_ VGND VGND VPWR VPWR _05975_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_17_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15829_ net2413 _13210_ _14236_ VGND VGND VPWR VPWR _14246_ sky130_fd_sc_hd__mux2_1
X_31875_ clknet_leaf_122_clk _03329_ VGND VGND VPWR VPWR datamem.data_ram\[56\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_19597_ datamem.data_ram\[54\]\[8\] _06626_ _06811_ datamem.data_ram\[48\]\[8\] VGND
+ VGND VPWR VPWR _06893_ sky130_fd_sc_hd__o22a_1
XFILLER_0_177_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_1295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18548_ _05883_ _05885_ _05888_ _05908_ VGND VGND VPWR VPWR _05909_ sky130_fd_sc_hd__or4_1
X_30826_ clknet_leaf_221_clk _02561_ VGND VGND VPWR VPWR datamem.data_ram\[44\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30757_ clknet_leaf_154_clk _02492_ VGND VGND VPWR VPWR datamem.data_ram\[47\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_153_clk clknet_5_28__leaf_clk VGND VGND VPWR VPWR clknet_leaf_153_clk
+ sky130_fd_sc_hd__clkbuf_8
X_18479_ _05838_ _05840_ _05676_ VGND VGND VPWR VPWR _05841_ sky130_fd_sc_hd__mux2_1
XFILLER_0_185_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20510_ _07131_ _07798_ _07800_ VGND VGND VPWR VPWR _07801_ sky130_fd_sc_hd__and3_1
XFILLER_0_145_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21490_ _08725_ _08745_ VGND VGND VPWR VPWR _08746_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_211_5556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30688_ clknet_leaf_258_clk _02423_ VGND VGND VPWR VPWR datamem.data_ram\[4\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_23988__523 clknet_1_1__leaf__10239_ VGND VGND VPWR VPWR net649 sky130_fd_sc_hd__inv_2
XFILLER_0_28_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_211_5567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32427_ clknet_leaf_247_clk _03849_ VGND VGND VPWR VPWR datamem.data_ram\[28\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_20441_ datamem.data_ram\[31\]\[12\] _06705_ _07732_ _06600_ VGND VGND VPWR VPWR
+ _07733_ sky130_fd_sc_hd__o211a_1
XFILLER_0_166_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload330 clknet_1_1__leaf__10130_ VGND VGND VPWR VPWR clkload330/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_207_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32358_ clknet_leaf_250_clk _03780_ VGND VGND VPWR VPWR datamem.data_ram\[30\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_20372_ datamem.data_ram\[42\]\[28\] _06608_ _06667_ datamem.data_ram\[47\]\[28\]
+ VGND VGND VPWR VPWR _07664_ sky130_fd_sc_hd__o22a_1
Xclkload341 clknet_1_0__leaf__10127_ VGND VGND VPWR VPWR clkload341/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload352 clknet_1_0__leaf__10089_ VGND VGND VPWR VPWR clkload352/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload60 clknet_leaf_7_clk VGND VGND VPWR VPWR clkload60/Y sky130_fd_sc_hd__inv_6
X_22111_ rvcpu.dp.plem.WriteDataM\[5\] _08488_ _09293_ VGND VGND VPWR VPWR _09320_
+ sky130_fd_sc_hd__and3_1
X_31309_ clknet_leaf_48_clk _03012_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCPlus4E\[15\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload71 clknet_leaf_70_clk VGND VGND VPWR VPWR clkload71/Y sky130_fd_sc_hd__inv_8
Xclkload82 clknet_leaf_43_clk VGND VGND VPWR VPWR clkload82/Y sky130_fd_sc_hd__clkinv_8
X_32289_ clknet_leaf_226_clk _03711_ VGND VGND VPWR VPWR datamem.data_ram\[32\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload93 clknet_leaf_74_clk VGND VGND VPWR VPWR clkload93/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_228_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22042_ _09263_ VGND VGND VPWR VPWR _09264_ sky130_fd_sc_hd__buf_4
Xhold2800 datamem.data_ram\[61\]\[10\] VGND VGND VPWR VPWR net3950 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2811 datamem.data_ram\[11\]\[11\] VGND VGND VPWR VPWR net3961 sky130_fd_sc_hd__dlygate4sd3_1
X_26850_ _11689_ _11786_ VGND VGND VPWR VPWR _11793_ sky130_fd_sc_hd__and2_1
XFILLER_0_220_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2822 datamem.data_ram\[22\]\[14\] VGND VGND VPWR VPWR net3972 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2833 datamem.data_ram\[26\]\[15\] VGND VGND VPWR VPWR net3983 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_162_4375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2844 datamem.data_ram\[46\]\[10\] VGND VGND VPWR VPWR net3994 sky130_fd_sc_hd__dlygate4sd3_1
X_25801_ _11191_ _11192_ _11149_ VGND VGND VPWR VPWR _11193_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_162_4386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2855 rvcpu.dp.rf.reg_file_arr\[27\]\[29\] VGND VGND VPWR VPWR net4005 sky130_fd_sc_hd__dlygate4sd3_1
X_26781_ _06587_ VGND VGND VPWR VPWR _11752_ sky130_fd_sc_hd__buf_2
Xhold2866 rvcpu.dp.rf.reg_file_arr\[31\]\[5\] VGND VGND VPWR VPWR net4016 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2877 datamem.data_ram\[58\]\[8\] VGND VGND VPWR VPWR net4027 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_173_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2888 datamem.data_ram\[39\]\[27\] VGND VGND VPWR VPWR net4038 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_104_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2899 datamem.data_ram\[29\]\[30\] VGND VGND VPWR VPWR net4049 sky130_fd_sc_hd__dlygate4sd3_1
X_25732_ _10824_ net1998 _11133_ VGND VGND VPWR VPWR _11140_ sky130_fd_sc_hd__mux2_1
X_28520_ _12748_ VGND VGND VPWR VPWR _04061_ sky130_fd_sc_hd__clkbuf_1
X_22944_ rvcpu.dp.plem.WriteDataM\[6\] VGND VGND VPWR VPWR _10072_ sky130_fd_sc_hd__buf_4
XFILLER_0_39_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_175_4703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25663_ _11081_ _11098_ VGND VGND VPWR VPWR _11100_ sky130_fd_sc_hd__and2_1
XFILLER_0_195_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28451_ _12707_ VGND VGND VPWR VPWR _04033_ sky130_fd_sc_hd__clkbuf_1
X_22875_ _09390_ _10010_ VGND VGND VPWR VPWR _10011_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27402_ _12089_ net2938 net85 VGND VGND VPWR VPWR _12121_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24614_ _10509_ VGND VGND VPWR VPWR _02394_ sky130_fd_sc_hd__clkbuf_1
X_28382_ _12666_ VGND VGND VPWR VPWR _04005_ sky130_fd_sc_hd__clkbuf_1
X_21826_ _08510_ _09064_ VGND VGND VPWR VPWR _09065_ sky130_fd_sc_hd__nor2_1
X_25594_ _11057_ net1420 _11053_ _11060_ VGND VGND VPWR VPWR _02823_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_121_3393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27333_ _09297_ VGND VGND VPWR VPWR _12080_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_93_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_183_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24545_ _10469_ VGND VGND VPWR VPWR _02365_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_144_clk clknet_5_29__leaf_clk VGND VGND VPWR VPWR clknet_leaf_144_clk
+ sky130_fd_sc_hd__clkbuf_8
X_21757_ rvcpu.dp.rf.reg_file_arr\[12\]\[19\] rvcpu.dp.rf.reg_file_arr\[13\]\[19\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[19\] rvcpu.dp.rf.reg_file_arr\[15\]\[19\] _08696_
+ _08553_ VGND VGND VPWR VPWR _09000_ sky130_fd_sc_hd__mux4_1
XFILLER_0_66_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_182_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20708_ datamem.data_ram\[24\]\[5\] _07138_ _06949_ datamem.data_ram\[25\]\[5\] VGND
+ VGND VPWR VPWR _07999_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27264_ _10838_ _10997_ _11713_ VGND VGND VPWR VPWR _12043_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_134_3710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24476_ _09326_ net4180 _10421_ VGND VGND VPWR VPWR _10428_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_3721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21688_ _08934_ VGND VGND VPWR VPWR _01043_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29003_ _12995_ net1780 _13009_ _13012_ VGND VGND VPWR VPWR _04280_ sky130_fd_sc_hd__a31o_1
X_26215_ _11445_ VGND VGND VPWR VPWR _03059_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_184_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27195_ _10402_ _10980_ VGND VGND VPWR VPWR _12006_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_24_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20639_ _06777_ _07922_ _07924_ _07929_ VGND VGND VPWR VPWR _07930_ sky130_fd_sc_hd__a31o_1
XFILLER_0_202_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_130_3607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_3618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26146_ _11409_ VGND VGND VPWR VPWR _03025_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23358_ clknet_1_0__leaf__10130_ VGND VGND VPWR VPWR _10138_ sky130_fd_sc_hd__buf_1
XFILLER_0_62_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23357__994 clknet_1_0__leaf__10137_ VGND VGND VPWR VPWR net1120 sky130_fd_sc_hd__inv_2
XFILLER_0_61_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22309_ _09473_ VGND VGND VPWR VPWR _09474_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_221_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26077_ _08622_ _11369_ VGND VGND VPWR VPWR _11370_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_219_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29905_ clknet_leaf_145_clk _01640_ VGND VGND VPWR VPWR datamem.data_ram\[59\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_25028_ _09290_ VGND VGND VPWR VPWR _10739_ sky130_fd_sc_hd__buf_2
X_23056__755 clknet_1_0__leaf__10091_ VGND VGND VPWR VPWR net881 sky130_fd_sc_hd__inv_2
XFILLER_0_219_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17850_ _13243_ rvcpu.dp.plde.RD2E\[11\] _05194_ VGND VGND VPWR VPWR _05228_ sky130_fd_sc_hd__mux2_1
X_29836_ net214 _01571_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[1\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_3558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_3569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16801_ _13179_ _14089_ VGND VGND VPWR VPWR _04647_ sky130_fd_sc_hd__nor2_2
XFILLER_0_79_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17781_ _05172_ _05173_ _05178_ net1293 VGND VGND VPWR VPWR rvcpu.dp.SrcBFW_Mux.y\[0\]
+ sky130_fd_sc_hd__o2bb2a_1
X_29767_ net1113 _01502_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[20\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_14993_ _13397_ _13371_ VGND VGND VPWR VPWR _13541_ sky130_fd_sc_hd__nor2_2
X_26979_ _11863_ net1711 _11865_ _11873_ VGND VGND VPWR VPWR _03395_ sky130_fd_sc_hd__a31o_1
X_19520_ datamem.data_ram\[62\]\[24\] _06626_ _06685_ datamem.data_ram\[60\]\[24\]
+ VGND VGND VPWR VPWR _06816_ sky130_fd_sc_hd__o22a_1
X_16732_ _04610_ VGND VGND VPWR VPWR _01676_ sky130_fd_sc_hd__clkbuf_1
X_28718_ _12702_ net2356 _12850_ VGND VGND VPWR VPWR _12858_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29698_ net1044 _01433_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[23\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19451_ datamem.data_ram\[45\]\[16\] _06724_ _06742_ _06746_ VGND VGND VPWR VPWR
+ _06747_ sky130_fd_sc_hd__o211a_1
X_16663_ _14195_ net4176 _04539_ VGND VGND VPWR VPWR _04574_ sky130_fd_sc_hd__mux2_1
X_28649_ _12821_ VGND VGND VPWR VPWR _04117_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18402_ _05342_ _05349_ _05358_ _05679_ _05683_ _05688_ VGND VGND VPWR VPWR _05766_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_202_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15614_ _14115_ VGND VGND VPWR VPWR _02199_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31660_ clknet_leaf_63_clk net1280 VGND VGND VPWR VPWR rvcpu.dp.plmw.ALUResultW\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_19382_ _06677_ VGND VGND VPWR VPWR _06678_ sky130_fd_sc_hd__buf_6
X_16594_ _14195_ net2096 _04502_ VGND VGND VPWR VPWR _04537_ sky130_fd_sc_hd__mux2_1
XFILLER_0_174_718 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18333_ _05697_ VGND VGND VPWR VPWR _05698_ sky130_fd_sc_hd__buf_2
X_30611_ clknet_leaf_195_clk _02346_ VGND VGND VPWR VPWR datamem.data_ram\[52\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_201_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15545_ _13649_ _14070_ _13442_ VGND VGND VPWR VPWR _14071_ sky130_fd_sc_hd__a21o_1
XFILLER_0_56_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31591_ clknet_leaf_52_clk net1234 VGND VGND VPWR VPWR rvcpu.dp.plmw.PCPlus4W\[9\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_135_clk clknet_5_30__leaf_clk VGND VGND VPWR VPWR clknet_leaf_135_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_16_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15476_ _13909_ _13811_ _14003_ _14004_ _13319_ VGND VGND VPWR VPWR _14005_ sky130_fd_sc_hd__o221a_1
XFILLER_0_189_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18264_ _05461_ _05467_ _05624_ _05628_ VGND VGND VPWR VPWR _05629_ sky130_fd_sc_hd__o31ai_2
X_30542_ clknet_leaf_148_clk _02277_ VGND VGND VPWR VPWR datamem.data_ram\[55\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17215_ _04867_ VGND VGND VPWR VPWR _01434_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18195_ _05284_ _05559_ VGND VGND VPWR VPWR _05560_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30473_ net151 _02208_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[19\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32212_ clknet_leaf_254_clk _03634_ VGND VGND VPWR VPWR datamem.data_ram\[36\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17146_ _14133_ net3574 _04829_ VGND VGND VPWR VPWR _04831_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold706 datamem.data_ram\[62\]\[6\] VGND VGND VPWR VPWR net1856 sky130_fd_sc_hd__dlygate4sd3_1
Xhold717 rvcpu.dp.pcreg.q\[21\] VGND VGND VPWR VPWR net1867 sky130_fd_sc_hd__dlygate4sd3_1
Xhold728 datamem.data_ram\[34\]\[1\] VGND VGND VPWR VPWR net1878 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17077_ _04794_ VGND VGND VPWR VPWR _01499_ sky130_fd_sc_hd__clkbuf_1
X_32143_ clknet_leaf_276_clk _03565_ VGND VGND VPWR VPWR datamem.data_ram\[39\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold739 rvcpu.dp.rf.reg_file_arr\[17\]\[21\] VGND VGND VPWR VPWR net1889 sky130_fd_sc_hd__dlygate4sd3_1
X_23489__135 clknet_1_0__leaf__10160_ VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__inv_2
X_16028_ net2583 _13195_ _14349_ VGND VGND VPWR VPWR _14354_ sky130_fd_sc_hd__mux2_1
X_32074_ clknet_leaf_94_clk _03496_ VGND VGND VPWR VPWR datamem.data_ram\[33\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31025_ clknet_leaf_58_clk _02760_ VGND VGND VPWR VPWR datamem.data_ram\[40\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2107 rvcpu.dp.rf.reg_file_arr\[6\]\[13\] VGND VGND VPWR VPWR net3257 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_62_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2118 datamem.data_ram\[8\]\[29\] VGND VGND VPWR VPWR net3268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2129 datamem.data_ram\[57\]\[31\] VGND VGND VPWR VPWR net3279 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23569__192 clknet_1_0__leaf__10175_ VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__inv_2
XFILLER_0_100_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1406 rvcpu.dp.rf.reg_file_arr\[8\]\[11\] VGND VGND VPWR VPWR net2556 sky130_fd_sc_hd__dlygate4sd3_1
X_23412__65 clknet_1_1__leaf__10153_ VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__inv_2
XFILLER_0_224_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_204_5382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1417 rvcpu.dp.rf.reg_file_arr\[31\]\[11\] VGND VGND VPWR VPWR net2567 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_204_5393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1428 datamem.data_ram\[32\]\[20\] VGND VGND VPWR VPWR net2578 sky130_fd_sc_hd__dlygate4sd3_1
X_17979_ _13259_ _05179_ _05180_ VGND VGND VPWR VPWR _05350_ sky130_fd_sc_hd__nand3b_1
Xhold1439 rvcpu.dp.rf.reg_file_arr\[19\]\[15\] VGND VGND VPWR VPWR net2589 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19718_ _06716_ _07008_ _07013_ _06713_ VGND VGND VPWR VPWR _07014_ sky130_fd_sc_hd__a31o_1
X_32976_ clknet_leaf_146_clk _04398_ VGND VGND VPWR VPWR datamem.data_ram\[63\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_20990_ datamem.data_ram\[2\]\[15\] datamem.data_ram\[3\]\[15\] _06650_ VGND VGND
+ VPWR VPWR _08279_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31927_ clknet_leaf_123_clk _03349_ VGND VGND VPWR VPWR datamem.data_ram\[60\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_196_5194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19649_ _06944_ _06934_ VGND VGND VPWR VPWR _06945_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_217_5710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22660_ _09433_ _09807_ _09789_ VGND VGND VPWR VPWR _09808_ sky130_fd_sc_hd__a21o_1
X_31858_ clknet_leaf_110_clk _03312_ VGND VGND VPWR VPWR datamem.data_ram\[62\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24055__583 clknet_1_0__leaf__10246_ VGND VGND VPWR VPWR net709 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_213_5607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_213_5618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21611_ _08695_ _08861_ VGND VGND VPWR VPWR _08862_ sky130_fd_sc_hd__and2_1
XFILLER_0_177_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30809_ clknet_leaf_152_clk _02544_ VGND VGND VPWR VPWR datamem.data_ram\[45\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_126_clk clknet_5_30__leaf_clk VGND VGND VPWR VPWR clknet_leaf_126_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_30_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22591_ _09734_ _09738_ _09742_ _09491_ VGND VGND VPWR VPWR _01138_ sky130_fd_sc_hd__o31a_1
X_31789_ clknet_leaf_104_clk _03243_ VGND VGND VPWR VPWR datamem.data_ram\[8\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24330_ _10341_ VGND VGND VPWR VPWR _02278_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21542_ _08557_ VGND VGND VPWR VPWR _08795_ sky130_fd_sc_hd__buf_2
XFILLER_0_63_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24261_ _09318_ net4099 _10298_ VGND VGND VPWR VPWR _10303_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21473_ _08627_ _08724_ _08727_ _08729_ VGND VGND VPWR VPWR _08730_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_161_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26000_ _09478_ _11315_ _11312_ _11324_ VGND VGND VPWR VPWR _02965_ sky130_fd_sc_hd__o211a_1
X_20424_ datamem.data_ram\[2\]\[12\] _06610_ _06815_ datamem.data_ram\[5\]\[12\] VGND
+ VGND VPWR VPWR _07716_ sky130_fd_sc_hd__o22a_1
XFILLER_0_120_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20355_ datamem.data_ram\[11\]\[28\] _06738_ VGND VGND VPWR VPWR _07647_ sky130_fd_sc_hd__or2_1
Xclkload160 clknet_leaf_179_clk VGND VGND VPWR VPWR clkload160/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_31_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload171 clknet_leaf_214_clk VGND VGND VPWR VPWR clkload171/Y sky130_fd_sc_hd__clkinv_4
Xclkload182 clknet_leaf_238_clk VGND VGND VPWR VPWR clkload182/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_219_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload193 clknet_leaf_227_clk VGND VGND VPWR VPWR clkload193/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_164_4426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_164_4437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27951_ _12369_ net4049 _12421_ VGND VGND VPWR VPWR _12428_ sky130_fd_sc_hd__mux2_1
X_23074_ _09285_ net3767 _10093_ VGND VGND VPWR VPWR _10099_ sky130_fd_sc_hd__mux2_1
X_20286_ datamem.data_ram\[26\]\[19\] _06613_ _07575_ _07578_ VGND VGND VPWR VPWR
+ _07579_ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26902_ _11825_ _11823_ VGND VGND VPWR VPWR _11826_ sky130_fd_sc_hd__and2_1
X_22025_ rvcpu.dp.plem.WriteDataM\[21\] _09220_ VGND VGND VPWR VPWR _09250_ sky130_fd_sc_hd__and2_1
X_27882_ _12157_ net2357 _12382_ VGND VGND VPWR VPWR _12390_ sky130_fd_sc_hd__mux2_1
XFILLER_0_216_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold11 rvcpu.dp.plem.PCPlus4M\[16\] VGND VGND VPWR VPWR net1161 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2630 datamem.data_ram\[46\]\[27\] VGND VGND VPWR VPWR net3780 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_216_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold22 rvcpu.dp.plde.PCPlus4E\[29\] VGND VGND VPWR VPWR net1172 sky130_fd_sc_hd__dlygate4sd3_1
X_29621_ net975 _01356_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[25\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold33 rvcpu.dp.plde.PCPlus4E\[5\] VGND VGND VPWR VPWR net1183 sky130_fd_sc_hd__dlygate4sd3_1
X_26833_ _11672_ _11774_ VGND VGND VPWR VPWR _11783_ sky130_fd_sc_hd__and2_1
Xhold2641 datamem.data_ram\[6\]\[17\] VGND VGND VPWR VPWR net3791 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 rvcpu.dp.plem.lAuiPCM\[23\] VGND VGND VPWR VPWR net1194 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2652 rvcpu.dp.rf.reg_file_arr\[18\]\[27\] VGND VGND VPWR VPWR net3802 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 rvcpu.dp.plem.PCPlus4M\[20\] VGND VGND VPWR VPWR net1205 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2663 datamem.data_ram\[55\]\[25\] VGND VGND VPWR VPWR net3813 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2674 rvcpu.dp.rf.reg_file_arr\[1\]\[14\] VGND VGND VPWR VPWR net3824 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 rvcpu.dp.plem.lAuiPCM\[27\] VGND VGND VPWR VPWR net1216 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1940 datamem.data_ram\[41\]\[30\] VGND VGND VPWR VPWR net3090 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2685 datamem.data_ram\[25\]\[26\] VGND VGND VPWR VPWR net3835 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_67_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold77 rvcpu.dp.plem.lAuiPCM\[16\] VGND VGND VPWR VPWR net1227 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1951 rvcpu.dp.rf.reg_file_arr\[12\]\[8\] VGND VGND VPWR VPWR net3101 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_67_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29552_ net906 _01287_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[27\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_26764_ _11684_ _11738_ VGND VGND VPWR VPWR _11742_ sky130_fd_sc_hd__and2_1
Xhold88 rvcpu.dp.plem.lAuiPCM\[8\] VGND VGND VPWR VPWR net1238 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2696 datamem.data_ram\[53\]\[28\] VGND VGND VPWR VPWR net3846 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 rvcpu.dp.plem.PCPlus4M\[10\] VGND VGND VPWR VPWR net1249 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_123_3444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1962 datamem.data_ram\[46\]\[11\] VGND VGND VPWR VPWR net3112 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_123_3455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1973 rvcpu.dp.rf.reg_file_arr\[23\]\[30\] VGND VGND VPWR VPWR net3123 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1984 rvcpu.dp.rf.reg_file_arr\[8\]\[24\] VGND VGND VPWR VPWR net3134 sky130_fd_sc_hd__dlygate4sd3_1
X_28503_ _09272_ VGND VGND VPWR VPWR _12737_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_196_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22927_ _10056_ net1732 _10046_ _10059_ VGND VGND VPWR VPWR _01157_ sky130_fd_sc_hd__a31o_1
Xhold1995 datamem.data_ram\[13\]\[18\] VGND VGND VPWR VPWR net3145 sky130_fd_sc_hd__dlygate4sd3_1
X_25715_ _10824_ net2682 _11124_ VGND VGND VPWR VPWR _11131_ sky130_fd_sc_hd__mux2_1
X_26695_ _11689_ _11694_ VGND VGND VPWR VPWR _11702_ sky130_fd_sc_hd__and2_1
Xclkbuf_1_1__f__10264_ clknet_0__10264_ VGND VGND VPWR VPWR clknet_1_1__leaf__10264_
+ sky130_fd_sc_hd__clkbuf_16
X_29483_ net845 _01218_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[2\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_211_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28434_ _12696_ net3349 _12688_ VGND VGND VPWR VPWR _12697_ sky130_fd_sc_hd__mux2_1
X_25646_ _11064_ _11079_ VGND VGND VPWR VPWR _11093_ sky130_fd_sc_hd__and2_1
XFILLER_0_196_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22858_ _09510_ _09988_ _09990_ _09994_ _09525_ VGND VGND VPWR VPWR _09995_ sky130_fd_sc_hd__a311o_1
XFILLER_0_97_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__10195_ clknet_0__10195_ VGND VGND VPWR VPWR clknet_1_1__leaf__10195_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_168_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21809_ rvcpu.dp.rf.reg_file_arr\[4\]\[22\] rvcpu.dp.rf.reg_file_arr\[5\]\[22\] rvcpu.dp.rf.reg_file_arr\[6\]\[22\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[22\] _08628_ _08856_ VGND VGND VPWR VPWR _09049_
+ sky130_fd_sc_hd__mux4_1
X_25577_ _11018_ net1470 _11041_ _11049_ VGND VGND VPWR VPWR _02817_ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_117_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_117_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_26_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28365_ _12657_ VGND VGND VPWR VPWR _03997_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22789_ _09636_ _09929_ VGND VGND VPWR VPWR _09930_ sky130_fd_sc_hd__or2_1
XFILLER_0_155_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15330_ _13430_ _13399_ VGND VGND VPWR VPWR _13867_ sky130_fd_sc_hd__nor2_1
XFILLER_0_186_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27316_ _11978_ _12066_ VGND VGND VPWR VPWR _12073_ sky130_fd_sc_hd__and2_1
X_24528_ _10459_ VGND VGND VPWR VPWR _02358_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28296_ _12620_ VGND VGND VPWR VPWR _03965_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_97_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15261_ _13430_ _13628_ _13484_ VGND VGND VPWR VPWR _13801_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27247_ _12036_ net1414 _12030_ _12037_ VGND VGND VPWR VPWR _03499_ sky130_fd_sc_hd__a31o_1
X_24459_ _10418_ _10406_ VGND VGND VPWR VPWR _10419_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17000_ _04752_ VGND VGND VPWR VPWR _01542_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_163_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15192_ _13392_ _13434_ _13423_ VGND VGND VPWR VPWR _13735_ sky130_fd_sc_hd__a21oi_1
X_27178_ _11965_ _11996_ VGND VGND VPWR VPWR _11997_ sky130_fd_sc_hd__and2_1
XFILLER_0_152_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_8 _06594_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26129_ _11400_ VGND VGND VPWR VPWR _03017_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18951_ _05806_ _05845_ _06048_ _05661_ _06288_ VGND VGND VPWR VPWR _06289_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_56_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17902_ _05274_ VGND VGND VPWR VPWR _05275_ sky130_fd_sc_hd__buf_2
XFILLER_0_24_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18882_ _05240_ _06211_ _06224_ VGND VGND VPWR VPWR rvcpu.ALUResultE\[21\] sky130_fd_sc_hd__a21o_1
XFILLER_0_197_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17833_ _05216_ VGND VGND VPWR VPWR rvcpu.dp.SrcBFW_Mux.y\[22\] sky130_fd_sc_hd__clkbuf_2
X_29819_ net197 _01554_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[1\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_218_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32830_ clknet_leaf_159_clk _04252_ VGND VGND VPWR VPWR datamem.data_ram\[12\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_17764_ rvcpu.dp.plem.RdM\[0\] VGND VGND VPWR VPWR _05162_ sky130_fd_sc_hd__inv_2
XFILLER_0_221_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14976_ _13335_ _13523_ VGND VGND VPWR VPWR _13524_ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19503_ _06596_ _06711_ _06798_ VGND VGND VPWR VPWR _06799_ sky130_fd_sc_hd__a21oi_4
X_16715_ _14179_ net3750 _04598_ VGND VGND VPWR VPWR _04602_ sky130_fd_sc_hd__mux2_1
X_32761_ clknet_leaf_254_clk _04183_ VGND VGND VPWR VPWR datamem.data_ram\[15\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17695_ _13190_ net3009 _05118_ VGND VGND VPWR VPWR _05122_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31712_ clknet_leaf_34_clk _03170_ VGND VGND VPWR VPWR rvcpu.dp.pcreg.q\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19434_ _06729_ VGND VGND VPWR VPWR _06730_ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_179_Right_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16646_ _04565_ VGND VGND VPWR VPWR _01717_ sky130_fd_sc_hd__clkbuf_1
X_32692_ clknet_leaf_253_clk _04114_ VGND VGND VPWR VPWR datamem.data_ram\[18\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_191_5080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31643_ clknet_leaf_29_clk net1194 VGND VGND VPWR VPWR rvcpu.dp.plmw.lAuiPCW\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_19365_ _06660_ VGND VGND VPWR VPWR _06661_ sky130_fd_sc_hd__buf_8
XFILLER_0_9_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22967__675 clknet_1_1__leaf__10082_ VGND VGND VPWR VPWR net801 sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_108_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_108_clk
+ sky130_fd_sc_hd__clkbuf_8
X_16577_ _04528_ VGND VGND VPWR VPWR _01757_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_191_5091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_225_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18316_ _05390_ _05392_ VGND VGND VPWR VPWR _05681_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15528_ _14009_ _14053_ _13706_ VGND VGND VPWR VPWR _14054_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31574_ clknet_leaf_72_clk datamem.rd_data_mem\[24\] VGND VGND VPWR VPWR rvcpu.dp.plmw.ReadDataW\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_19296_ _06591_ _05347_ VGND VGND VPWR VPWR _06592_ sky130_fd_sc_hd__nor2_8
XFILLER_0_17_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18247_ net105 _05310_ VGND VGND VPWR VPWR _05612_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30525_ clknet_leaf_267_clk _02260_ VGND VGND VPWR VPWR datamem.data_ram\[56\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_15459_ _13665_ _13346_ _13484_ _13639_ _13581_ VGND VGND VPWR VPWR _13989_ sky130_fd_sc_hd__a311o_1
XFILLER_0_143_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18178_ _05541_ _05542_ VGND VGND VPWR VPWR _05543_ sky130_fd_sc_hd__nor2_2
X_30456_ net134 _02191_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[19\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold503 rvcpu.dp.plfd.PCPlus4D\[23\] VGND VGND VPWR VPWR net1653 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold514 datamem.data_ram\[51\]\[2\] VGND VGND VPWR VPWR net1664 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17129_ _04821_ VGND VGND VPWR VPWR _01474_ sky130_fd_sc_hd__clkbuf_1
Xhold525 rvcpu.dp.plfd.PCPlus4D\[14\] VGND VGND VPWR VPWR net1675 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_229_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold536 datamem.data_ram\[2\]\[3\] VGND VGND VPWR VPWR net1686 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30387_ clknet_leaf_174_clk _02122_ VGND VGND VPWR VPWR datamem.data_ram\[58\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold547 datamem.data_ram\[16\]\[1\] VGND VGND VPWR VPWR net1697 sky130_fd_sc_hd__dlygate4sd3_1
Xhold558 datamem.data_ram\[17\]\[2\] VGND VGND VPWR VPWR net1708 sky130_fd_sc_hd__dlygate4sd3_1
X_20140_ datamem.data_ram\[45\]\[27\] _06721_ _06654_ datamem.data_ram\[41\]\[27\]
+ VGND VGND VPWR VPWR _07433_ sky130_fd_sc_hd__o22a_1
X_32126_ clknet_leaf_215_clk _03548_ VGND VGND VPWR VPWR datamem.data_ram\[7\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold569 datamem.data_ram\[63\]\[1\] VGND VGND VPWR VPWR net1719 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_206_5433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_206_5444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32057_ clknet_leaf_119_clk _03479_ VGND VGND VPWR VPWR datamem.data_ram\[48\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_20071_ _07348_ _07353_ _07359_ _07364_ VGND VGND VPWR VPWR _07365_ sky130_fd_sc_hd__o22a_1
X_23725__317 clknet_1_1__leaf__10198_ VGND VGND VPWR VPWR net443 sky130_fd_sc_hd__inv_2
X_31008_ clknet_leaf_163_clk _02743_ VGND VGND VPWR VPWR datamem.data_ram\[11\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1203 datamem.data_ram\[34\]\[21\] VGND VGND VPWR VPWR net2353 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_198_5245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1214 datamem.data_ram\[42\]\[15\] VGND VGND VPWR VPWR net2364 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_198_5256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1225 rvcpu.dp.pcreg.q\[18\] VGND VGND VPWR VPWR net2375 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_1053 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23830_ _10211_ VGND VGND VPWR VPWR _01908_ sky130_fd_sc_hd__clkbuf_1
Xhold1236 datamem.data_ram\[30\]\[31\] VGND VGND VPWR VPWR net2386 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1247 datamem.data_ram\[55\]\[15\] VGND VGND VPWR VPWR net2397 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1258 datamem.data_ram\[14\]\[9\] VGND VGND VPWR VPWR net2408 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1269 rvcpu.dp.rf.reg_file_arr\[16\]\[15\] VGND VGND VPWR VPWR net2419 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_197_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_178_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32959_ clknet_leaf_84_clk _04381_ VGND VGND VPWR VPWR datamem.data_ram\[6\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20973_ datamem.data_ram\[40\]\[15\] datamem.data_ram\[41\]\[15\] _06652_ VGND VGND
+ VPWR VPWR _08262_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_409 _06645_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_221_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25500_ _10822_ net3221 _10999_ VGND VGND VPWR VPWR _11005_ sky130_fd_sc_hd__mux2_1
X_22712_ _09442_ _09852_ _09854_ _09856_ VGND VGND VPWR VPWR _09857_ sky130_fd_sc_hd__o2bb2a_1
X_26480_ _11261_ _11253_ _11597_ _11598_ VGND VGND VPWR VPWR _11599_ sky130_fd_sc_hd__o211ai_1
X_26496__49 clknet_1_0__leaf__11601_ VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__inv_2
XFILLER_0_215_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_146_Right_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_178_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_157_4252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_4263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25431_ _10754_ net3724 _10970_ VGND VGND VPWR VPWR _10972_ sky130_fd_sc_hd__mux2_1
Xclkbuf_0__10080_ _10080_ VGND VGND VPWR VPWR clknet_0__10080_ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_157_4274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22643_ rvcpu.dp.rf.reg_file_arr\[8\]\[17\] rvcpu.dp.rf.reg_file_arr\[10\]\[17\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[17\] rvcpu.dp.rf.reg_file_arr\[11\]\[17\] _09608_
+ _09532_ VGND VGND VPWR VPWR _09792_ sky130_fd_sc_hd__mux4_1
XFILLER_0_137_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_554 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25362_ _10418_ _10923_ VGND VGND VPWR VPWR _10930_ sky130_fd_sc_hd__and2_1
X_28150_ _12541_ VGND VGND VPWR VPWR _03898_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22574_ rvcpu.dp.rf.reg_file_arr\[16\]\[14\] rvcpu.dp.rf.reg_file_arr\[17\]\[14\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[14\] rvcpu.dp.rf.reg_file_arr\[19\]\[14\] _09445_
+ _09447_ VGND VGND VPWR VPWR _09726_ sky130_fd_sc_hd__mux4_1
XFILLER_0_90_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27101_ _11938_ net1693 _11940_ _11947_ VGND VGND VPWR VPWR _03443_ sky130_fd_sc_hd__a31o_1
XFILLER_0_145_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23771__359 clknet_1_1__leaf__10202_ VGND VGND VPWR VPWR net485 sky130_fd_sc_hd__inv_2
X_24313_ _09314_ net2971 _10328_ VGND VGND VPWR VPWR _10332_ sky130_fd_sc_hd__mux2_1
X_28081_ _12437_ net3286 _12501_ VGND VGND VPWR VPWR _12505_ sky130_fd_sc_hd__mux2_1
X_21525_ rvcpu.dp.rf.reg_file_arr\[20\]\[8\] rvcpu.dp.rf.reg_file_arr\[21\]\[8\] rvcpu.dp.rf.reg_file_arr\[22\]\[8\]
+ rvcpu.dp.rf.reg_file_arr\[23\]\[8\] _08778_ _08632_ VGND VGND VPWR VPWR _08779_
+ sky130_fd_sc_hd__mux4_1
X_25293_ _10889_ VGND VGND VPWR VPWR _02693_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_146_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_185_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27032_ _11803_ _11899_ VGND VGND VPWR VPWR _11905_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_116_3270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24244_ _10293_ VGND VGND VPWR VPWR _02240_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21456_ rvcpu.dp.rf.reg_file_arr\[0\]\[4\] rvcpu.dp.rf.reg_file_arr\[1\]\[4\] rvcpu.dp.rf.reg_file_arr\[2\]\[4\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[4\] _08550_ _08554_ VGND VGND VPWR VPWR _08714_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_116_3281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20407_ datamem.data_ram\[47\]\[12\] _06704_ _06780_ datamem.data_ram\[41\]\[12\]
+ VGND VGND VPWR VPWR _07699_ sky130_fd_sc_hd__o22a_1
X_23886__446 clknet_1_1__leaf__10222_ VGND VGND VPWR VPWR net572 sky130_fd_sc_hd__inv_2
X_21387_ rvcpu.dp.rf.reg_file_arr\[12\]\[1\] rvcpu.dp.rf.reg_file_arr\[13\]\[1\] rvcpu.dp.rf.reg_file_arr\[14\]\[1\]
+ rvcpu.dp.rf.reg_file_arr\[15\]\[1\] _08567_ _08570_ VGND VGND VPWR VPWR _08648_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_187_4982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_187_4993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput12 net12 VGND VGND VPWR VPWR Instr[19] sky130_fd_sc_hd__buf_2
XFILLER_0_120_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_3178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput23 net23 VGND VGND VPWR VPWR Instr[29] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_112_3189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24105__613 clknet_1_0__leaf__10258_ VGND VGND VPWR VPWR net739 sky130_fd_sc_hd__inv_2
X_20338_ datamem.data_ram\[33\]\[4\] _07133_ _07626_ _07629_ VGND VGND VPWR VPWR _07630_
+ sky130_fd_sc_hd__a211o_1
Xoutput34 net113 VGND VGND VPWR VPWR correct sky130_fd_sc_hd__buf_2
X_28983_ _12690_ net3720 _12999_ VGND VGND VPWR VPWR _13001_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_183_4879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27934_ _12138_ net4352 _12412_ VGND VGND VPWR VPWR _12419_ sky130_fd_sc_hd__mux2_1
X_20269_ _06681_ _07554_ _07556_ _07561_ VGND VGND VPWR VPWR _07562_ sky130_fd_sc_hd__a31o_1
Xhold3150 datamem.data_ram\[52\]\[11\] VGND VGND VPWR VPWR net4300 sky130_fd_sc_hd__dlygate4sd3_1
X_22008_ _09236_ net4336 _09232_ VGND VGND VPWR VPWR _09237_ sky130_fd_sc_hd__mux2_1
Xhold3161 datamem.data_ram\[62\]\[20\] VGND VGND VPWR VPWR net4311 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_125_3506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3172 rvcpu.dp.rf.reg_file_arr\[14\]\[8\] VGND VGND VPWR VPWR net4322 sky130_fd_sc_hd__dlygate4sd3_1
X_23665__264 clknet_1_0__leaf__10191_ VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__inv_2
X_27865_ _12140_ net2439 _12373_ VGND VGND VPWR VPWR _12381_ sky130_fd_sc_hd__mux2_1
Xhold3183 datamem.data_ram\[4\]\[20\] VGND VGND VPWR VPWR net4333 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3194 datamem.data_ram\[24\]\[14\] VGND VGND VPWR VPWR net4344 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2460 datamem.data_ram\[37\]\[14\] VGND VGND VPWR VPWR net3610 sky130_fd_sc_hd__dlygate4sd3_1
X_29604_ net958 _01339_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[25\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_26816_ _11772_ VGND VGND VPWR VPWR _11773_ sky130_fd_sc_hd__buf_2
X_14830_ _13282_ _13330_ VGND VGND VPWR VPWR _13383_ sky130_fd_sc_hd__nor2_1
Xhold2471 datamem.data_ram\[57\]\[8\] VGND VGND VPWR VPWR net3621 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2482 datamem.data_ram\[14\]\[8\] VGND VGND VPWR VPWR net3632 sky130_fd_sc_hd__dlygate4sd3_1
X_27796_ _12132_ net3140 _12336_ VGND VGND VPWR VPWR _12340_ sky130_fd_sc_hd__mux2_1
Xhold2493 datamem.data_ram\[21\]\[15\] VGND VGND VPWR VPWR net3643 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1770 datamem.data_ram\[33\]\[17\] VGND VGND VPWR VPWR net2920 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_187_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29535_ net889 _01270_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[27\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_4_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26747_ _11700_ net1845 _11724_ _11731_ VGND VGND VPWR VPWR _03305_ sky130_fd_sc_hd__a31o_1
X_14761_ _13313_ VGND VGND VPWR VPWR _13314_ sky130_fd_sc_hd__clkbuf_4
Xhold1781 datamem.data_ram\[42\]\[10\] VGND VGND VPWR VPWR net2931 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1792 datamem.data_ram\[39\]\[22\] VGND VGND VPWR VPWR net2942 sky130_fd_sc_hd__dlygate4sd3_1
X_23959_ _10233_ VGND VGND VPWR VPWR _02015_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_142_3897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16500_ _04487_ VGND VGND VPWR VPWR _01793_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14692_ _13253_ VGND VGND VPWR VPWR _13254_ sky130_fd_sc_hd__clkbuf_8
X_29466_ net828 _01201_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[2\]\[5\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__10247_ clknet_0__10247_ VGND VGND VPWR VPWR clknet_1_1__leaf__10247_
+ sky130_fd_sc_hd__clkbuf_16
X_17480_ _05007_ VGND VGND VPWR VPWR _01301_ sky130_fd_sc_hd__clkbuf_1
X_26678_ _11683_ net1855 _11675_ _11691_ VGND VGND VPWR VPWR _03276_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_113_Right_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_224_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_690 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16431_ net4132 _14461_ _14572_ VGND VGND VPWR VPWR _14582_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28417_ _12685_ VGND VGND VPWR VPWR _04021_ sky130_fd_sc_hd__clkbuf_1
X_25629_ _11081_ _11079_ VGND VGND VPWR VPWR _11082_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29397_ clknet_leaf_1_clk _01132_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD2E\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__10178_ clknet_0__10178_ VGND VGND VPWR VPWR clknet_1_1__leaf__10178_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_39_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19150_ _06457_ VGND VGND VPWR VPWR _06466_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28348_ _12648_ VGND VGND VPWR VPWR _03989_ sky130_fd_sc_hd__clkbuf_1
X_16362_ _14545_ VGND VGND VPWR VPWR _01857_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_45_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18101_ rvcpu.dp.plde.RD1E\[21\] _05292_ _05468_ VGND VGND VPWR VPWR _05469_ sky130_fd_sc_hd__o21a_2
XFILLER_0_13_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15313_ _13392_ VGND VGND VPWR VPWR _13850_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19081_ _06405_ VGND VGND VPWR VPWR rvcpu.dp.lAuiPCE\[8\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16293_ net4073 _14459_ _14500_ VGND VGND VPWR VPWR _14509_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28279_ _12371_ net3729 _12603_ VGND VGND VPWR VPWR _12611_ sky130_fd_sc_hd__mux2_1
X_18032_ _05358_ _05359_ VGND VGND VPWR VPWR _05402_ sky130_fd_sc_hd__nand2_1
X_30310_ net656 _02045_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[5\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_15244_ _13777_ _13778_ _13783_ _13501_ VGND VGND VPWR VPWR _13784_ sky130_fd_sc_hd__o211a_1
XFILLER_0_152_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31290_ clknet_leaf_76_clk _02993_ VGND VGND VPWR VPWR rvcpu.dp.plde.MemWriteE sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15175_ _13320_ _13349_ _13430_ VGND VGND VPWR VPWR _13718_ sky130_fd_sc_hd__o21a_1
X_30241_ net595 _01976_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[7\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30172_ net534 _01907_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[0\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_19983_ _06911_ _06580_ _06582_ VGND VGND VPWR VPWR _07277_ sky130_fd_sc_hd__o21a_2
XFILLER_0_162_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18934_ _06159_ _06272_ _05697_ VGND VGND VPWR VPWR _06273_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_193_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18865_ _06199_ _06206_ _06208_ VGND VGND VPWR VPWR _06209_ sky130_fd_sc_hd__or3b_1
XFILLER_0_206_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_201_5330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17816_ _13194_ rvcpu.dp.plde.RD2E\[27\] _05196_ VGND VGND VPWR VPWR _05205_ sky130_fd_sc_hd__mux2_1
X_18796_ _05658_ _05771_ _05720_ _06143_ _06004_ VGND VGND VPWR VPWR _06144_ sky130_fd_sc_hd__o221a_1
XFILLER_0_27_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_19_Left_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32813_ clknet_leaf_286_clk _04235_ VGND VGND VPWR VPWR datamem.data_ram\[13\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_222_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_193_5120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17747_ _13269_ net3605 _05140_ VGND VGND VPWR VPWR _05149_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_193_5131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14959_ _13307_ _13505_ _13507_ _13402_ VGND VGND VPWR VPWR _13508_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_178_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32744_ clknet_leaf_284_clk _04166_ VGND VGND VPWR VPWR datamem.data_ram\[16\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_17678_ _05112_ VGND VGND VPWR VPWR _01200_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19417_ _06712_ VGND VGND VPWR VPWR _06713_ sky130_fd_sc_hd__buf_6
X_16629_ _04556_ VGND VGND VPWR VPWR _01725_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32675_ clknet_leaf_239_clk _04097_ VGND VGND VPWR VPWR datamem.data_ram\[18\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31626_ clknet_leaf_64_clk net1211 VGND VGND VPWR VPWR rvcpu.dp.plmw.lAuiPCW\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19348_ _06643_ VGND VGND VPWR VPWR _06644_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_190_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31557_ clknet_leaf_64_clk datamem.rd_data_mem\[7\] VGND VGND VPWR VPWR rvcpu.dp.plmw.ReadDataW\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_19279_ _06570_ rvcpu.dp.plfd.InstrD\[12\] rvcpu.dp.plfd.InstrD\[13\] VGND VGND VPWR
+ VPWR _06577_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_150_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_28_Left_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21310_ _08541_ VGND VGND VPWR VPWR _08572_ sky130_fd_sc_hd__clkbuf_8
X_30508_ clknet_leaf_175_clk _02243_ VGND VGND VPWR VPWR datamem.data_ram\[57\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22290_ _09452_ _09454_ VGND VGND VPWR VPWR _09455_ sky130_fd_sc_hd__nor2_1
X_31488_ clknet_leaf_48_clk rvcpu.dp.lAuiPCE\[14\] VGND VGND VPWR VPWR rvcpu.dp.plem.lAuiPCM\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold300 datamem.data_ram\[32\]\[3\] VGND VGND VPWR VPWR net1450 sky130_fd_sc_hd__dlygate4sd3_1
X_21241_ datamem.data_ram\[52\]\[0\] datamem.data_ram\[53\]\[0\] _08502_ _08503_ VGND
+ VGND VPWR VPWR _08504_ sky130_fd_sc_hd__or4_2
Xhold311 datamem.data_ram\[38\]\[1\] VGND VGND VPWR VPWR net1461 sky130_fd_sc_hd__dlygate4sd3_1
X_30439_ net777 _02174_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[29\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold322 datamem.data_ram\[5\]\[3\] VGND VGND VPWR VPWR net1472 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__10267_ clknet_0__10267_ VGND VGND VPWR VPWR clknet_1_0__leaf__10267_
+ sky130_fd_sc_hd__clkbuf_16
Xhold333 datamem.data_ram\[36\]\[4\] VGND VGND VPWR VPWR net1483 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold344 datamem.data_ram\[15\]\[5\] VGND VGND VPWR VPWR net1494 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold355 datamem.data_ram\[38\]\[5\] VGND VGND VPWR VPWR net1505 sky130_fd_sc_hd__dlygate4sd3_1
X_21172_ _07866_ _08456_ _08458_ _08460_ VGND VGND VPWR VPWR _08461_ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold366 datamem.data_ram\[30\]\[1\] VGND VGND VPWR VPWR net1516 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold377 datamem.data_ram\[13\]\[1\] VGND VGND VPWR VPWR net1527 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__10198_ clknet_0__10198_ VGND VGND VPWR VPWR clknet_1_0__leaf__10198_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_111_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold388 datamem.data_ram\[28\]\[5\] VGND VGND VPWR VPWR net1538 sky130_fd_sc_hd__dlygate4sd3_1
X_32109_ clknet_leaf_120_clk _03531_ VGND VGND VPWR VPWR datamem.data_ram\[58\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_20123_ _06915_ _07276_ _07416_ VGND VGND VPWR VPWR _04437_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_111_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold399 datamem.data_ram\[55\]\[4\] VGND VGND VPWR VPWR net1549 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_225_5886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25980_ net1705 _11302_ _11312_ _11313_ VGND VGND VPWR VPWR _02956_ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_225_5897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_215_Right_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_176_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24931_ _10476_ net3888 net91 VGND VGND VPWR VPWR _10684_ sky130_fd_sc_hd__mux2_1
X_20054_ _06678_ _07345_ _07347_ VGND VGND VPWR VPWR _07348_ sky130_fd_sc_hd__and3_1
Xhold1000 rvcpu.dp.rf.reg_file_arr\[6\]\[31\] VGND VGND VPWR VPWR net2150 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_0_Left_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_225_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1011 rvcpu.dp.rf.reg_file_arr\[18\]\[9\] VGND VGND VPWR VPWR net2161 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1022 datamem.data_ram\[51\]\[0\] VGND VGND VPWR VPWR net2172 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_37_Left_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27650_ _10520_ _12106_ _12260_ VGND VGND VPWR VPWR _12261_ sky130_fd_sc_hd__a21oi_1
Xhold1033 datamem.data_ram\[2\]\[15\] VGND VGND VPWR VPWR net2183 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1044 rvcpu.dp.rf.reg_file_arr\[9\]\[11\] VGND VGND VPWR VPWR net2194 sky130_fd_sc_hd__dlygate4sd3_1
X_24862_ _10396_ net3367 net93 VGND VGND VPWR VPWR _10647_ sky130_fd_sc_hd__mux2_1
XFILLER_0_225_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1055 datamem.data_ram\[3\]\[21\] VGND VGND VPWR VPWR net2205 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_159_4303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26601_ _11091_ _11640_ VGND VGND VPWR VPWR _11648_ sky130_fd_sc_hd__and2_1
Xhold1066 rvcpu.dp.rf.reg_file_arr\[9\]\[12\] VGND VGND VPWR VPWR net2216 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_159_4314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1077 rvcpu.dp.rf.reg_file_arr\[20\]\[19\] VGND VGND VPWR VPWR net2227 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_1_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27581_ _10741_ _10908_ _12168_ VGND VGND VPWR VPWR _12224_ sky130_fd_sc_hd__a21oi_4
X_24793_ _10478_ net3609 _10602_ VGND VGND VPWR VPWR _10609_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1088 rvcpu.dp.rf.reg_file_arr\[0\]\[26\] VGND VGND VPWR VPWR net2238 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1099 datamem.data_ram\[19\]\[22\] VGND VGND VPWR VPWR net2249 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_206 _09560_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0__10201_ _10201_ VGND VGND VPWR VPWR clknet_0__10201_ sky130_fd_sc_hd__clkbuf_16
X_29320_ clknet_leaf_12_clk _01055_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD1E\[27\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_217 _09786_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_228 _10072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26532_ _10051_ VGND VGND VPWR VPWR _11609_ sky130_fd_sc_hd__clkbuf_4
X_23744_ clknet_1_0__leaf__10192_ VGND VGND VPWR VPWR _10200_ sky130_fd_sc_hd__buf_1
XANTENNA_239 _10783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20956_ datamem.data_ram\[50\]\[15\] datamem.data_ram\[51\]\[15\] _06652_ VGND VGND
+ VPWR VPWR _08245_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0__10132_ _10132_ VGND VGND VPWR VPWR clknet_0__10132_ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_81_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29251_ _09247_ net3989 _13141_ VGND VGND VPWR VPWR _13146_ sky130_fd_sc_hd__mux2_1
X_26463_ _11535_ rvcpu.ALUResultE\[26\] _11288_ VGND VGND VPWR VPWR _11587_ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20887_ _07839_ _08174_ _08176_ _07844_ VGND VGND VPWR VPWR _08177_ sky130_fd_sc_hd__a211o_1
XFILLER_0_49_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_187_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28202_ _12456_ net4228 net46 VGND VGND VPWR VPWR _12569_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25414_ _10754_ net3995 _10961_ VGND VGND VPWR VPWR _10963_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22626_ _09627_ _09773_ _09775_ _09438_ VGND VGND VPWR VPWR _09776_ sky130_fd_sc_hd__a211o_1
X_26394_ _11161_ _11526_ VGND VGND VPWR VPWR _11538_ sky130_fd_sc_hd__nand2_1
X_29182_ _13108_ VGND VGND VPWR VPWR _04363_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_118_3321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25345_ _07791_ _10918_ _10897_ VGND VGND VPWR VPWR _10919_ sky130_fd_sc_hd__or3_1
X_28133_ _12532_ VGND VGND VPWR VPWR _03890_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_46_Left_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22557_ _09391_ _09709_ VGND VGND VPWR VPWR _09710_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_114_3229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21508_ rvcpu.dp.rf.reg_file_arr\[28\]\[7\] rvcpu.dp.rf.reg_file_arr\[30\]\[7\] rvcpu.dp.rf.reg_file_arr\[29\]\[7\]
+ rvcpu.dp.rf.reg_file_arr\[31\]\[7\] _08635_ _08637_ VGND VGND VPWR VPWR _08763_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_228_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_540 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28064_ _12363_ net4271 _12492_ VGND VGND VPWR VPWR _12496_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25276_ _10880_ VGND VGND VPWR VPWR _02685_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22488_ rvcpu.dp.rf.reg_file_arr\[8\]\[9\] rvcpu.dp.rf.reg_file_arr\[10\]\[9\] rvcpu.dp.rf.reg_file_arr\[9\]\[9\]
+ rvcpu.dp.rf.reg_file_arr\[11\]\[9\] _09418_ _09485_ VGND VGND VPWR VPWR _09645_
+ sky130_fd_sc_hd__mux4_1
X_23020__724 clknet_1_0__leaf__10086_ VGND VGND VPWR VPWR net850 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_79_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27015_ _11835_ _11886_ VGND VGND VPWR VPWR _11894_ sky130_fd_sc_hd__and2_1
XFILLER_0_134_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24227_ _10284_ VGND VGND VPWR VPWR _02232_ sky130_fd_sc_hd__clkbuf_1
X_21439_ _08695_ _08697_ VGND VGND VPWR VPWR _08698_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23135__811 clknet_1_1__leaf__10106_ VGND VGND VPWR VPWR net937 sky130_fd_sc_hd__inv_2
X_28966_ _12727_ net1519 _12988_ _12991_ VGND VGND VPWR VPWR _04264_ sky130_fd_sc_hd__a31o_1
XFILLER_0_21_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16980_ _04719_ VGND VGND VPWR VPWR _04742_ sky130_fd_sc_hd__buf_4
X_24089_ _10256_ VGND VGND VPWR VPWR _02122_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_55_Left_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_88_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15931_ _14301_ VGND VGND VPWR VPWR _02060_ sky130_fd_sc_hd__clkbuf_1
X_27917_ _12155_ net1995 net47 VGND VGND VPWR VPWR _12410_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28897_ _12953_ VGND VGND VPWR VPWR _04233_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_144_3948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_552 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18650_ _05965_ _06005_ _05768_ VGND VGND VPWR VPWR _06006_ sky130_fd_sc_hd__mux2_1
X_27848_ _12371_ net2386 _12357_ VGND VGND VPWR VPWR _12372_ sky130_fd_sc_hd__mux2_1
X_15862_ _14263_ VGND VGND VPWR VPWR _02091_ sky130_fd_sc_hd__clkbuf_1
Xhold2290 rvcpu.dp.rf.reg_file_arr\[8\]\[30\] VGND VGND VPWR VPWR net3440 sky130_fd_sc_hd__dlygate4sd3_1
X_17601_ _13254_ net3163 _05068_ VGND VGND VPWR VPWR _05072_ sky130_fd_sc_hd__mux2_1
XFILLER_0_203_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14813_ _13312_ _13365_ VGND VGND VPWR VPWR _13366_ sky130_fd_sc_hd__nand2_4
XFILLER_0_189_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18581_ _05799_ _05796_ VGND VGND VPWR VPWR _05940_ sky130_fd_sc_hd__nor2_1
X_27779_ _12330_ VGND VGND VPWR VPWR _03738_ sky130_fd_sc_hd__clkbuf_1
X_15793_ _14226_ VGND VGND VPWR VPWR _02131_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_203_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17532_ _05035_ VGND VGND VPWR VPWR _01277_ sky130_fd_sc_hd__clkbuf_1
X_29518_ net880 _01253_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[28\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_14744_ _13296_ VGND VGND VPWR VPWR _13297_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_153_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_47_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30790_ clknet_leaf_172_clk _02525_ VGND VGND VPWR VPWR datamem.data_ram\[46\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17463_ _14177_ net4092 _04996_ VGND VGND VPWR VPWR _04999_ sky130_fd_sc_hd__mux2_1
X_29449_ net811 _01184_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[30\]\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_103_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14675_ _13240_ VGND VGND VPWR VPWR _13241_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_103_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19202_ _06509_ _06511_ VGND VGND VPWR VPWR _06512_ sky130_fd_sc_hd__xnor2_1
X_16414_ _14573_ VGND VGND VPWR VPWR _01833_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_64_Left_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32460_ clknet_leaf_246_clk _03882_ VGND VGND VPWR VPWR datamem.data_ram\[26\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_17394_ _04962_ VGND VGND VPWR VPWR _01342_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_144_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19133_ _06449_ _06450_ VGND VGND VPWR VPWR _06451_ sky130_fd_sc_hd__or2b_1
X_31411_ clknet_leaf_22_clk _03114_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCE\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16345_ net2497 _14442_ _14536_ VGND VGND VPWR VPWR _14537_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23222__872 clknet_1_0__leaf__10124_ VGND VGND VPWR VPWR net998 sky130_fd_sc_hd__inv_2
X_32391_ clknet_leaf_184_clk _03813_ VGND VGND VPWR VPWR datamem.data_ram\[29\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19064_ _06381_ _06390_ VGND VGND VPWR VPWR _06391_ sky130_fd_sc_hd__nor2_1
X_31342_ clknet_leaf_13_clk _03045_ VGND VGND VPWR VPWR rvcpu.dp.plde.Rs1E\[3\] sky130_fd_sc_hd__dfxtp_1
X_16276_ _14488_ VGND VGND VPWR VPWR _14500_ sky130_fd_sc_hd__buf_4
X_18015_ rvcpu.dp.plem.ALUResultM\[1\] _05175_ _05181_ _05182_ _05276_ VGND VGND VPWR
+ VPWR _05385_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_23_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23439__90 clknet_1_0__leaf__10155_ VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__inv_2
X_15227_ _13506_ _13767_ _13432_ _13357_ VGND VGND VPWR VPWR _13768_ sky130_fd_sc_hd__or4_1
XFILLER_0_164_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31273_ clknet_leaf_22_clk _02976_ VGND VGND VPWR VPWR rvcpu.dp.plfd.InstrD\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30224_ net578 _01959_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[7\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15158_ _13328_ _13330_ _13458_ _13701_ _13572_ VGND VGND VPWR VPWR _13702_ sky130_fd_sc_hd__o311a_1
XFILLER_0_196_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_199_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15089_ _13428_ _13634_ VGND VGND VPWR VPWR _13635_ sky130_fd_sc_hd__nand2_1
X_19966_ datamem.data_ram\[10\]\[18\] _06610_ _06821_ datamem.data_ram\[8\]\[18\]
+ VGND VGND VPWR VPWR _07260_ sky130_fd_sc_hd__o22a_1
X_30155_ net517 _01890_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[0\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_1047 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18917_ _05677_ _06201_ _06256_ VGND VGND VPWR VPWR _06257_ sky130_fd_sc_hd__a21o_1
X_19897_ datamem.data_ram\[6\]\[17\] _07028_ _06621_ datamem.data_ram\[4\]\[17\] VGND
+ VGND VPWR VPWR _07192_ sky130_fd_sc_hd__o22a_1
X_30086_ net448 _01821_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[11\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18848_ _05886_ _06191_ _06192_ VGND VGND VPWR VPWR _06193_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_220_5772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_220_5783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1271 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18779_ _05741_ _05658_ _06029_ _06127_ VGND VGND VPWR VPWR _06128_ sky130_fd_sc_hd__o31a_1
XFILLER_0_136_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20810_ datamem.data_ram\[41\]\[30\] _06947_ _08099_ _07867_ VGND VGND VPWR VPWR
+ _08100_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_19_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_960 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21790_ rvcpu.dp.rf.reg_file_arr\[12\]\[21\] rvcpu.dp.rf.reg_file_arr\[13\]\[21\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[21\] rvcpu.dp.rf.reg_file_arr\[15\]\[21\] _08578_
+ _08684_ VGND VGND VPWR VPWR _09031_ sky130_fd_sc_hd__mux4_1
X_30988_ clknet_leaf_90_clk _02723_ VGND VGND VPWR VPWR datamem.data_ram\[39\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_19_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_194_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20741_ datamem.data_ram\[41\]\[6\] _07839_ _07845_ _07832_ VGND VGND VPWR VPWR _08031_
+ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_154_4200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23540__165 clknet_1_0__leaf__10173_ VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__inv_2
X_32727_ clknet_leaf_184_clk _04149_ VGND VGND VPWR VPWR datamem.data_ram\[16\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32658_ clknet_leaf_81_clk _04080_ VGND VGND VPWR VPWR datamem.data_ram\[19\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_20672_ _06715_ _07946_ _07951_ _07962_ VGND VGND VPWR VPWR _07963_ sky130_fd_sc_hd__o31a_1
XFILLER_0_9_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22411_ rvcpu.dp.rf.reg_file_arr\[8\]\[5\] rvcpu.dp.rf.reg_file_arr\[10\]\[5\] rvcpu.dp.rf.reg_file_arr\[9\]\[5\]
+ rvcpu.dp.rf.reg_file_arr\[11\]\[5\] _09483_ _09485_ VGND VGND VPWR VPWR _09572_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_190_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_698 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31609_ clknet_leaf_25_clk net1223 VGND VGND VPWR VPWR rvcpu.dp.plmw.PCPlus4W\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23391_ _10146_ VGND VGND VPWR VPWR _01534_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32589_ clknet_leaf_171_clk _04011_ VGND VGND VPWR VPWR datamem.data_ram\[21\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_30_clk clknet_5_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_30_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_171_4591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25130_ _10472_ net2846 net87 VGND VGND VPWR VPWR _10797_ sky130_fd_sc_hd__mux2_1
X_22342_ rvcpu.dp.rf.reg_file_arr\[12\]\[2\] rvcpu.dp.rf.reg_file_arr\[13\]\[2\] rvcpu.dp.rf.reg_file_arr\[14\]\[2\]
+ rvcpu.dp.rf.reg_file_arr\[15\]\[2\] _09478_ _09479_ VGND VGND VPWR VPWR _09506_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_147_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25061_ _10759_ VGND VGND VPWR VPWR _02591_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22273_ _09429_ _09432_ _09436_ _09438_ VGND VGND VPWR VPWR _09439_ sky130_fd_sc_hd__a211o_1
XFILLER_0_170_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_227_5937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_227_5948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24012_ clknet_1_1__leaf__10224_ VGND VGND VPWR VPWR _10242_ sky130_fd_sc_hd__buf_1
XFILLER_0_182_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold130 rvcpu.dp.plem.ALUResultM\[8\] VGND VGND VPWR VPWR net1280 sky130_fd_sc_hd__dlygate4sd3_1
X_21224_ _08468_ _07691_ _08489_ VGND VGND VPWR VPWR _04435_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_148_4037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold141 rvcpu.dp.plfd.PCD\[17\] VGND VGND VPWR VPWR net1291 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_148_4048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold152 datamem.data_ram\[47\]\[3\] VGND VGND VPWR VPWR net1302 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_4059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold163 datamem.data_ram\[41\]\[4\] VGND VGND VPWR VPWR net1313 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold174 rvcpu.dp.plem.ALUResultM\[18\] VGND VGND VPWR VPWR net1324 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_180_4805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28820_ _12912_ VGND VGND VPWR VPWR _04197_ sky130_fd_sc_hd__clkbuf_1
Xhold185 datamem.data_ram\[44\]\[1\] VGND VGND VPWR VPWR net1335 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_180_4816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21155_ datamem.data_ram\[24\]\[23\] datamem.data_ram\[25\]\[23\] datamem.data_ram\[26\]\[23\]
+ datamem.data_ram\[27\]\[23\] _06933_ _07819_ VGND VGND VPWR VPWR _08444_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_180_4827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold196 datamem.data_ram\[47\]\[7\] VGND VGND VPWR VPWR net1346 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_6_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20106_ datamem.data_ram\[15\]\[10\] _06672_ _07396_ _07399_ VGND VGND VPWR VPWR
+ _07400_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_70_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28751_ _12875_ VGND VGND VPWR VPWR _04165_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_217_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21086_ datamem.data_ram\[32\]\[7\] _06935_ _08372_ _08374_ VGND VGND VPWR VPWR _08375_
+ sky130_fd_sc_hd__a211o_1
X_25963_ net1270 _11302_ _11300_ _11304_ VGND VGND VPWR VPWR _02948_ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_97_clk clknet_5_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_97_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27702_ _12279_ _12106_ _12260_ VGND VGND VPWR VPWR _12289_ sky130_fd_sc_hd__a21oi_4
X_20037_ datamem.data_ram\[18\]\[26\] _06690_ _06662_ datamem.data_ram\[21\]\[26\]
+ _06678_ VGND VGND VPWR VPWR _07331_ sky130_fd_sc_hd__o221a_1
X_24914_ _10396_ net3049 _10669_ VGND VGND VPWR VPWR _10675_ sky130_fd_sc_hd__mux2_1
X_28682_ _12764_ net2954 _12832_ VGND VGND VPWR VPWR _12839_ sky130_fd_sc_hd__mux2_1
X_25894_ net1884 _11263_ VGND VGND VPWR VPWR _11265_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_107_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27633_ _12125_ net2507 _12251_ VGND VGND VPWR VPWR _12252_ sky130_fd_sc_hd__mux2_1
XFILLER_0_225_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24845_ _10637_ VGND VGND VPWR VPWR _02497_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_217_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_178_4756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_178_4767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_4778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23165__837 clknet_1_1__leaf__10110_ VGND VGND VPWR VPWR net963 sky130_fd_sc_hd__inv_2
X_27564_ _10741_ _10898_ _12168_ VGND VGND VPWR VPWR _12215_ sky130_fd_sc_hd__a21oi_1
X_21988_ rvcpu.dp.plem.MemWriteM _06911_ _09217_ VGND VGND VPWR VPWR _09218_ sky130_fd_sc_hd__and3_1
X_24776_ _07125_ VGND VGND VPWR VPWR _10598_ sky130_fd_sc_hd__buf_8
XFILLER_0_179_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29303_ clknet_leaf_1_clk _01038_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD1E\[10\] sky130_fd_sc_hd__dfxtp_1
X_23703__297 clknet_1_0__leaf__10196_ VGND VGND VPWR VPWR net423 sky130_fd_sc_hd__inv_2
XFILLER_0_90_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20939_ datamem.data_ram\[50\]\[22\] datamem.data_ram\[51\]\[22\] _07835_ VGND VGND
+ VPWR VPWR _08229_ sky130_fd_sc_hd__mux2_1
X_27495_ _07132_ VGND VGND VPWR VPWR _12178_ sky130_fd_sc_hd__buf_8
XFILLER_0_113_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29234_ _09317_ net3920 _13132_ VGND VGND VPWR VPWR _13137_ sky130_fd_sc_hd__mux2_1
X_26446_ net4454 _11573_ _11575_ _11570_ VGND VGND VPWR VPWR _03160_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_42_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29165_ _13099_ VGND VGND VPWR VPWR _04355_ sky130_fd_sc_hd__clkbuf_1
X_22609_ _09759_ VGND VGND VPWR VPWR _01139_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26377_ _08620_ _08621_ _11151_ VGND VGND VPWR VPWR _11525_ sky130_fd_sc_hd__a21o_1
XFILLER_0_153_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_3774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_21_clk clknet_5_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_21_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_137_3785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_221_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28116_ _12523_ VGND VGND VPWR VPWR _03882_ sky130_fd_sc_hd__clkbuf_1
X_16130_ net2434 _13244_ _14407_ VGND VGND VPWR VPWR _14408_ sky130_fd_sc_hd__mux2_1
X_25328_ _10751_ net4217 _10909_ VGND VGND VPWR VPWR _10910_ sky130_fd_sc_hd__mux2_1
X_29096_ _09317_ net2958 net40 VGND VGND VPWR VPWR _13063_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28047_ _12454_ net3485 net96 VGND VGND VPWR VPWR _12487_ sky130_fd_sc_hd__mux2_1
X_16061_ _14348_ VGND VGND VPWR VPWR _14371_ sky130_fd_sc_hd__clkbuf_4
X_25259_ _10410_ _10868_ VGND VGND VPWR VPWR _10871_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15012_ _13305_ _13323_ VGND VGND VPWR VPWR _13560_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_209_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19820_ datamem.data_ram\[29\]\[9\] _06703_ _07113_ _07114_ VGND VGND VPWR VPWR _07115_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29998_ net368 _01733_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[14\]\[25\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_36_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19751_ datamem.data_ram\[43\]\[25\] _06863_ _07042_ _07045_ VGND VGND VPWR VPWR
+ _07046_ sky130_fd_sc_hd__o211a_1
XFILLER_0_159_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28949_ _12981_ VGND VGND VPWR VPWR _04257_ sky130_fd_sc_hd__clkbuf_1
X_16963_ _04733_ VGND VGND VPWR VPWR _01560_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24003__536 clknet_1_0__leaf__10241_ VGND VGND VPWR VPWR net662 sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_88_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_88_clk sky130_fd_sc_hd__clkbuf_8
X_18702_ _05809_ VGND VGND VPWR VPWR _06055_ sky130_fd_sc_hd__clkbuf_4
X_15914_ _14292_ VGND VGND VPWR VPWR _02068_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_217_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31960_ clknet_leaf_122_clk _03382_ VGND VGND VPWR VPWR datamem.data_ram\[28\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_19682_ _06951_ VGND VGND VPWR VPWR _06978_ sky130_fd_sc_hd__buf_4
XFILLER_0_204_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16894_ net2456 _14445_ _04695_ VGND VGND VPWR VPWR _04697_ sky130_fd_sc_hd__mux2_1
XFILLER_0_200_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18633_ _05363_ _05692_ VGND VGND VPWR VPWR _05990_ sky130_fd_sc_hd__nand2_2
X_30911_ clknet_leaf_263_clk _02646_ VGND VGND VPWR VPWR datamem.data_ram\[41\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15845_ _14254_ VGND VGND VPWR VPWR _02099_ sky130_fd_sc_hd__clkbuf_1
X_31891_ clknet_leaf_114_clk _03345_ VGND VGND VPWR VPWR datamem.data_ram\[36\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18564_ _05790_ _05917_ _05919_ _05921_ _05923_ VGND VGND VPWR VPWR _05924_ sky130_fd_sc_hd__o2111a_1
X_30842_ clknet_leaf_180_clk _02577_ VGND VGND VPWR VPWR datamem.data_ram\[44\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_15776_ _14217_ VGND VGND VPWR VPWR _02139_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_176_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_72_Left_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17515_ _05026_ VGND VGND VPWR VPWR _01285_ sky130_fd_sc_hd__clkbuf_1
X_14727_ rvcpu.dp.pcreg.q\[2\] VGND VGND VPWR VPWR _13280_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_169_470 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18495_ _05855_ _05856_ _05676_ VGND VGND VPWR VPWR _05857_ sky130_fd_sc_hd__mux2_1
X_30773_ clknet_leaf_220_clk _02508_ VGND VGND VPWR VPWR datamem.data_ram\[46\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_570 rvcpu.dp.plmw.ReadDataW\[24\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32512_ clknet_leaf_185_clk _03934_ VGND VGND VPWR VPWR datamem.data_ram\[24\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17446_ _14160_ net3676 _04985_ VGND VGND VPWR VPWR _04990_ sky130_fd_sc_hd__mux2_1
X_14658_ rvcpu.dp.plmw.ALUResultW\[16\] rvcpu.dp.plmw.ReadDataW\[16\] rvcpu.dp.plmw.PCPlus4W\[16\]
+ rvcpu.dp.plmw.lAuiPCW\[16\] _13192_ _13193_ VGND VGND VPWR VPWR _13228_ sky130_fd_sc_hd__mux4_2
XFILLER_0_129_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_200_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32443_ clknet_leaf_77_clk _03865_ VGND VGND VPWR VPWR datamem.data_ram\[27\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17377_ _04953_ VGND VGND VPWR VPWR _01350_ sky130_fd_sc_hd__clkbuf_1
X_14589_ rvcpu.dp.plmw.RdW\[2\] VGND VGND VPWR VPWR _13174_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_12_clk clknet_5_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_131_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19116_ _06434_ _06435_ VGND VGND VPWR VPWR _06436_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16328_ net2403 _14426_ _14525_ VGND VGND VPWR VPWR _14528_ sky130_fd_sc_hd__mux2_1
X_32374_ clknet_leaf_278_clk _03796_ VGND VGND VPWR VPWR datamem.data_ram\[2\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19047_ _06368_ _06370_ _06367_ VGND VGND VPWR VPWR _06376_ sky130_fd_sc_hd__a21boi_2
X_31325_ clknet_leaf_23_clk _03028_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCPlus4E\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16259_ _14491_ VGND VGND VPWR VPWR _01906_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_81_Left_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31256_ clknet_leaf_20_clk _02959_ VGND VGND VPWR VPWR rvcpu.dp.plfd.InstrD\[14\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_207_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__10104_ clknet_0__10104_ VGND VGND VPWR VPWR clknet_1_0__leaf__10104_
+ sky130_fd_sc_hd__clkbuf_16
X_30207_ net561 _01942_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[8\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_222_5812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31187_ clknet_leaf_38_clk _02890_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCPlus4D\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_222_5823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_222_5834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30138_ net500 _01873_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[10\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_19949_ _07242_ VGND VGND VPWR VPWR _07243_ sky130_fd_sc_hd__clkbuf_8
Xclkbuf_leaf_79_clk clknet_5_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_79_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_96_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30069_ net431 _01804_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[12\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21911_ rvcpu.dp.rf.reg_file_arr\[20\]\[28\] rvcpu.dp.rf.reg_file_arr\[21\]\[28\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[28\] rvcpu.dp.rf.reg_file_arr\[23\]\[28\] _08516_
+ _08518_ VGND VGND VPWR VPWR _09145_ sky130_fd_sc_hd__mux4_1
XFILLER_0_218_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22891_ _09398_ _10025_ VGND VGND VPWR VPWR _10026_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_90_Left_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_222_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24630_ _10452_ net2263 _10511_ VGND VGND VPWR VPWR _10518_ sky130_fd_sc_hd__mux2_1
X_21842_ rvcpu.dp.rf.reg_file_arr\[24\]\[24\] rvcpu.dp.rf.reg_file_arr\[25\]\[24\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[24\] rvcpu.dp.rf.reg_file_arr\[27\]\[24\] _08525_
+ _08528_ VGND VGND VPWR VPWR _09080_ sky130_fd_sc_hd__mux4_1
X_23622__240 clknet_1_0__leaf__10180_ VGND VGND VPWR VPWR net366 sky130_fd_sc_hd__inv_2
XFILLER_0_195_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23229__878 clknet_1_0__leaf__10125_ VGND VGND VPWR VPWR net1004 sky130_fd_sc_hd__inv_2
XFILLER_0_167_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24561_ _09329_ VGND VGND VPWR VPWR _10480_ sky130_fd_sc_hd__clkbuf_2
X_21773_ _08813_ _09014_ _08689_ VGND VGND VPWR VPWR _09015_ sky130_fd_sc_hd__a21o_1
XFILLER_0_176_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26300_ net1326 _11478_ VGND VGND VPWR VPWR _11483_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_173_4642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20724_ _07823_ datamem.data_ram\[18\]\[6\] datamem.data_ram\[19\]\[6\] _07837_ _07840_
+ VGND VGND VPWR VPWR _08014_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_173_4653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23512_ _10164_ VGND VGND VPWR VPWR _01637_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24492_ _10436_ VGND VGND VPWR VPWR _02345_ sky130_fd_sc_hd__clkbuf_1
X_27280_ _12051_ VGND VGND VPWR VPWR _03518_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_190_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26231_ rvcpu.dp.plfd.InstrD\[7\] _06573_ _11371_ VGND VGND VPWR VPWR _11456_ sky130_fd_sc_hd__and3_1
XFILLER_0_135_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_190_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20655_ datamem.data_ram\[33\]\[29\] _06783_ _07942_ _07945_ VGND VGND VPWR VPWR
+ _07946_ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_184_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26162_ net4448 _11408_ VGND VGND VPWR VPWR _11418_ sky130_fd_sc_hd__and2_1
XFILLER_0_184_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20586_ _07821_ _07873_ _07876_ _06940_ VGND VGND VPWR VPWR _07877_ sky130_fd_sc_hd__a22o_1
XFILLER_0_225_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22325_ _09476_ _09480_ _09487_ _09489_ VGND VGND VPWR VPWR _09490_ sky130_fd_sc_hd__o211a_1
X_25113_ _10731_ net3483 net88 VGND VGND VPWR VPWR _10788_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_76_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26093_ _11381_ VGND VGND VPWR VPWR _03000_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_225_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_3671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29921_ net291 _01656_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[16\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_25044_ _10748_ VGND VGND VPWR VPWR _02585_ sky130_fd_sc_hd__clkbuf_1
X_23418__71 clknet_1_0__leaf__10153_ VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__inv_2
XFILLER_0_182_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_72_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22256_ _09421_ VGND VGND VPWR VPWR _09422_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_72_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21207_ _06987_ _08298_ _08471_ _08486_ VGND VGND VPWR VPWR _04421_ sky130_fd_sc_hd__a211o_1
X_29852_ net230 _01587_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[18\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_22187_ _09244_ net4400 _09362_ VGND VGND VPWR VPWR _09366_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_218_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28803_ _12903_ VGND VGND VPWR VPWR _04189_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_109_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21138_ _08424_ _08425_ _08426_ _07820_ _07866_ VGND VGND VPWR VPWR _08427_ sky130_fd_sc_hd__a221o_1
X_29783_ net1129 _01518_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[20\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26995_ _10764_ net3463 _11875_ VGND VGND VPWR VPWR _11882_ sky130_fd_sc_hd__mux2_1
X_28734_ _12866_ VGND VGND VPWR VPWR _04157_ sky130_fd_sc_hd__clkbuf_1
X_21069_ _06666_ datamem.data_ram\[63\]\[7\] _06944_ datamem.data_ram\[62\]\[7\] _07838_
+ VGND VGND VPWR VPWR _08358_ sky130_fd_sc_hd__a221o_1
X_25946_ net1819 _11155_ VGND VGND VPWR VPWR _11295_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_31_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28665_ _12700_ net1940 _12823_ VGND VGND VPWR VPWR _12830_ sky130_fd_sc_hd__mux2_1
X_25877_ rvcpu.dp.plfd.PCPlus4D\[31\] _11253_ _08598_ VGND VGND VPWR VPWR _11254_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27616_ _12080_ net3103 net80 VGND VGND VPWR VPWR _12243_ sky130_fd_sc_hd__mux2_1
X_15630_ _14123_ VGND VGND VPWR VPWR _02191_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_213_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24828_ _10398_ net2566 _10621_ VGND VGND VPWR VPWR _10628_ sky130_fd_sc_hd__mux2_1
XFILLER_0_216_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28596_ _12747_ net2224 _12786_ VGND VGND VPWR VPWR _12793_ sky130_fd_sc_hd__mux2_1
XFILLER_0_213_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15561_ _13398_ _13767_ _13458_ _13378_ VGND VGND VPWR VPWR _14085_ sky130_fd_sc_hd__a211o_1
X_27547_ _10542_ _12106_ _12168_ VGND VGND VPWR VPWR _12206_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_139_3825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24759_ _10297_ _10327_ _10501_ VGND VGND VPWR VPWR _10589_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_96_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_3836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17300_ _04912_ VGND VGND VPWR VPWR _01394_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18280_ _05561_ _05644_ VGND VGND VPWR VPWR _05645_ sky130_fd_sc_hd__or2_1
X_15492_ _13308_ _13654_ VGND VGND VPWR VPWR _14020_ sky130_fd_sc_hd__nor2_1
X_27478_ _10113_ _10908_ _12168_ VGND VGND VPWR VPWR _12169_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_29_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29217_ _10066_ _13123_ VGND VGND VPWR VPWR _13128_ sky130_fd_sc_hd__and2_1
XFILLER_0_194_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17231_ _04875_ VGND VGND VPWR VPWR _01426_ sky130_fd_sc_hd__clkbuf_1
X_26429_ net1904 _11542_ _11563_ _11534_ VGND VGND VPWR VPWR _03155_ sky130_fd_sc_hd__o211a_1
XFILLER_0_193_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_495 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17162_ _14149_ net4287 _04829_ VGND VGND VPWR VPWR _04839_ sky130_fd_sc_hd__mux2_1
X_29148_ _13090_ VGND VGND VPWR VPWR _04347_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16113_ net2160 _13220_ _14396_ VGND VGND VPWR VPWR _14399_ sky130_fd_sc_hd__mux2_1
X_29079_ _12760_ net2818 _13049_ VGND VGND VPWR VPWR _13054_ sky130_fd_sc_hd__mux2_1
X_17093_ _04802_ VGND VGND VPWR VPWR _01491_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31110_ clknet_leaf_60_clk _02845_ VGND VGND VPWR VPWR datamem.data_ram\[43\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_16044_ _14362_ VGND VGND VPWR VPWR _02000_ sky130_fd_sc_hd__clkbuf_1
X_32090_ clknet_leaf_212_clk _03512_ VGND VGND VPWR VPWR datamem.data_ram\[8\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31041_ clknet_leaf_98_clk _02776_ VGND VGND VPWR VPWR datamem.data_ram\[41\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23334__973 clknet_1_0__leaf__10135_ VGND VGND VPWR VPWR net1099 sky130_fd_sc_hd__inv_2
X_19803_ datamem.data_ram\[13\]\[9\] _06865_ _06688_ datamem.data_ram\[12\]\[9\] _07097_
+ VGND VGND VPWR VPWR _07098_ sky130_fd_sc_hd__o221a_1
X_17995_ rvcpu.dp.plde.RD1E\[4\] _05291_ _05364_ VGND VGND VPWR VPWR _05365_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_208_168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16946_ _04724_ VGND VGND VPWR VPWR _01568_ sky130_fd_sc_hd__clkbuf_1
X_19734_ datamem.data_ram\[0\]\[25\] _06698_ _06688_ datamem.data_ram\[4\]\[25\] VGND
+ VGND VPWR VPWR _07029_ sky130_fd_sc_hd__o22a_1
XFILLER_0_223_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_1_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_8
X_32992_ clknet_leaf_202_clk _04414_ VGND VGND VPWR VPWR datamem.data_ram\[62\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19665_ _06941_ VGND VGND VPWR VPWR _06961_ sky130_fd_sc_hd__buf_4
X_31943_ clknet_leaf_115_clk _03365_ VGND VGND VPWR VPWR datamem.data_ram\[32\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_223_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16877_ net2728 _14428_ _04684_ VGND VGND VPWR VPWR _04688_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_216_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23113__791 clknet_1_1__leaf__10104_ VGND VGND VPWR VPWR net917 sky130_fd_sc_hd__inv_2
XFILLER_0_79_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_189_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18616_ _05808_ VGND VGND VPWR VPWR _05974_ sky130_fd_sc_hd__buf_2
XFILLER_0_204_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15828_ _14245_ VGND VGND VPWR VPWR _02107_ sky130_fd_sc_hd__clkbuf_1
X_31874_ clknet_leaf_111_clk _03328_ VGND VGND VPWR VPWR datamem.data_ram\[56\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19596_ datamem.data_ram\[53\]\[8\] _06815_ _06670_ datamem.data_ram\[55\]\[8\] VGND
+ VGND VPWR VPWR _06892_ sky130_fd_sc_hd__o22a_1
XFILLER_0_59_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18547_ _05889_ _05894_ _05899_ _05837_ _05907_ VGND VGND VPWR VPWR _05908_ sky130_fd_sc_hd__a32o_1
XFILLER_0_48_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30825_ clknet_leaf_220_clk _02560_ VGND VGND VPWR VPWR datamem.data_ram\[44\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_15759_ _14208_ VGND VGND VPWR VPWR _02147_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18478_ _05839_ _05760_ _05668_ VGND VGND VPWR VPWR _05840_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30756_ clknet_leaf_178_clk _02491_ VGND VGND VPWR VPWR datamem.data_ram\[48\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_215_5660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17429_ _14143_ net4346 _04974_ VGND VGND VPWR VPWR _04981_ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30687_ clknet_leaf_264_clk _02422_ VGND VGND VPWR VPWR datamem.data_ram\[4\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_211_5557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_211_5568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20440_ datamem.data_ram\[30\]\[12\] _06743_ _06617_ datamem.data_ram\[28\]\[12\]
+ _07731_ VGND VGND VPWR VPWR _07732_ sky130_fd_sc_hd__o221a_1
X_32426_ clknet_leaf_258_clk _03848_ VGND VGND VPWR VPWR datamem.data_ram\[28\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32357_ clknet_leaf_242_clk _03779_ VGND VGND VPWR VPWR datamem.data_ram\[30\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_20371_ datamem.data_ram\[44\]\[28\] _06685_ _06655_ datamem.data_ram\[41\]\[28\]
+ VGND VGND VPWR VPWR _07663_ sky130_fd_sc_hd__o22a_1
Xclkload320 clknet_1_1__leaf__10158_ VGND VGND VPWR VPWR clkload320/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_141_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload331 clknet_1_0__leaf__10140_ VGND VGND VPWR VPWR clkload331/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_3_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload342 clknet_1_1__leaf__10126_ VGND VGND VPWR VPWR clkload342/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload50 clknet_leaf_69_clk VGND VGND VPWR VPWR clkload50/Y sky130_fd_sc_hd__clkinvlp_2
X_22110_ _09319_ VGND VGND VPWR VPWR _01080_ sky130_fd_sc_hd__clkbuf_1
Xclkload353 clknet_1_0__leaf__10088_ VGND VGND VPWR VPWR clkload353/Y sky130_fd_sc_hd__clkinvlp_4
X_31308_ clknet_leaf_49_clk _03011_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCPlus4E\[14\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload61 clknet_leaf_76_clk VGND VGND VPWR VPWR clkload61/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_30_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload72 clknet_leaf_54_clk VGND VGND VPWR VPWR clkload72/Y sky130_fd_sc_hd__clkinvlp_2
X_32288_ clknet_leaf_277_clk _03710_ VGND VGND VPWR VPWR datamem.data_ram\[33\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload83 clknet_leaf_46_clk VGND VGND VPWR VPWR clkload83/Y sky130_fd_sc_hd__inv_6
XFILLER_0_3_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload94 clknet_leaf_75_clk VGND VGND VPWR VPWR clkload94/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22041_ rvcpu.dp.plem.ALUResultM\[0\] net117 _09262_ VGND VGND VPWR VPWR _09263_
+ sky130_fd_sc_hd__and3_1
X_31239_ clknet_leaf_35_clk _02942_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCD\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_166_4490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2801 datamem.data_ram\[26\]\[24\] VGND VGND VPWR VPWR net3951 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2812 datamem.data_ram\[27\]\[13\] VGND VGND VPWR VPWR net3962 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2823 rvcpu.dp.rf.reg_file_arr\[26\]\[14\] VGND VGND VPWR VPWR net3973 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2834 datamem.data_ram\[0\]\[14\] VGND VGND VPWR VPWR net3984 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25800_ rvcpu.dp.pcreg.q\[16\] _11188_ VGND VGND VPWR VPWR _11192_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_215_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_162_4376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2845 datamem.data_ram\[11\]\[17\] VGND VGND VPWR VPWR net3995 sky130_fd_sc_hd__dlygate4sd3_1
X_26780_ _11735_ net1719 _11748_ _11751_ VGND VGND VPWR VPWR _03318_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_162_4387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2856 datamem.data_ram\[57\]\[23\] VGND VGND VPWR VPWR net4006 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2867 datamem.data_ram\[17\]\[12\] VGND VGND VPWR VPWR net4017 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2878 rvcpu.dp.rf.reg_file_arr\[0\]\[4\] VGND VGND VPWR VPWR net4028 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2889 datamem.data_ram\[42\]\[9\] VGND VGND VPWR VPWR net4039 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_104_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25731_ _11139_ VGND VGND VPWR VPWR _02881_ sky130_fd_sc_hd__clkbuf_1
X_22943_ _10056_ net1554 _10046_ _10071_ VGND VGND VPWR VPWR _01161_ sky130_fd_sc_hd__a31o_1
X_23546__171 clknet_1_0__leaf__10173_ VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__inv_2
XFILLER_0_39_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28450_ _12435_ net4149 _12704_ VGND VGND VPWR VPWR _12707_ sky130_fd_sc_hd__mux2_1
X_25662_ _11085_ net1861 _11097_ _11099_ VGND VGND VPWR VPWR _02852_ sky130_fd_sc_hd__a31o_1
XFILLER_0_190_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_175_4704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22874_ rvcpu.dp.rf.reg_file_arr\[24\]\[30\] rvcpu.dp.rf.reg_file_arr\[25\]\[30\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[30\] rvcpu.dp.rf.reg_file_arr\[27\]\[30\] _08592_
+ _08595_ VGND VGND VPWR VPWR _10010_ sky130_fd_sc_hd__mux4_1
XFILLER_0_218_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27401_ _12120_ VGND VGND VPWR VPWR _03570_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_65_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24613_ _10478_ net1949 _10502_ VGND VGND VPWR VPWR _10509_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28381_ _12369_ net3641 _12659_ VGND VGND VPWR VPWR _12666_ sky130_fd_sc_hd__mux2_1
X_21825_ _08795_ _09059_ _09061_ _09063_ VGND VGND VPWR VPWR _09064_ sky130_fd_sc_hd__o2bb2a_1
X_25593_ _10413_ _11055_ VGND VGND VPWR VPWR _11060_ sky130_fd_sc_hd__and2_1
XFILLER_0_167_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_3394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27332_ _10783_ _12076_ _12077_ net1764 VGND VGND VPWR VPWR _03542_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_210_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21756_ rvcpu.dp.rf.reg_file_arr\[8\]\[19\] rvcpu.dp.rf.reg_file_arr\[10\]\[19\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[19\] rvcpu.dp.rf.reg_file_arr\[11\]\[19\] _08534_
+ _08818_ VGND VGND VPWR VPWR _08999_ sky130_fd_sc_hd__mux4_1
X_24544_ _10468_ net3860 net60 VGND VGND VPWR VPWR _10469_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20707_ _07992_ _07997_ _07154_ VGND VGND VPWR VPWR _07998_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_1022 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27263_ _10783_ _12041_ _12042_ net1346 VGND VGND VPWR VPWR _03510_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_134_3700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_3711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24475_ _10427_ VGND VGND VPWR VPWR _02337_ sky130_fd_sc_hd__clkbuf_1
X_21687_ _08672_ _08925_ _08929_ _08933_ VGND VGND VPWR VPWR _08934_ sky130_fd_sc_hd__and4_1
XFILLER_0_110_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29002_ _10057_ _13010_ VGND VGND VPWR VPWR _13012_ sky130_fd_sc_hd__and2_1
XFILLER_0_191_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_134_3722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26214_ net1296 _11436_ _11444_ VGND VGND VPWR VPWR _11445_ sky130_fd_sc_hd__and3_1
Xclkload0 clknet_5_0__leaf_clk VGND VGND VPWR VPWR clkload0/Y sky130_fd_sc_hd__clkinv_4
Xwire115 _05171_ VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_4_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20638_ _06602_ _07926_ _07928_ VGND VGND VPWR VPWR _07929_ sky130_fd_sc_hd__and3_1
X_27194_ _11918_ VGND VGND VPWR VPWR _12005_ sky130_fd_sc_hd__buf_2
XFILLER_0_191_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_1276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23815__398 clknet_1_1__leaf__10207_ VGND VGND VPWR VPWR net524 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_130_3608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_190_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26145_ net1770 _11408_ VGND VGND VPWR VPWR _11409_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_130_3619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20569_ _07859_ VGND VGND VPWR VPWR _07860_ sky130_fd_sc_hd__buf_6
XFILLER_0_116_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22308_ rvcpu.dp.plfd.InstrD\[24\] _09472_ VGND VGND VPWR VPWR _09473_ sky130_fd_sc_hd__nor2_1
X_26076_ rvcpu.dp.plfd.InstrD\[3\] rvcpu.dp.plfd.InstrD\[2\] rvcpu.dp.plfd.InstrD\[0\]
+ _11366_ VGND VGND VPWR VPWR _11369_ sky130_fd_sc_hd__and4_1
XFILLER_0_46_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29904_ clknet_leaf_141_clk _01639_ VGND VGND VPWR VPWR datamem.data_ram\[59\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_25027_ _10738_ VGND VGND VPWR VPWR _02578_ sky130_fd_sc_hd__clkbuf_1
X_22239_ _09399_ _09403_ _09404_ VGND VGND VPWR VPWR _09405_ sky130_fd_sc_hd__o21a_1
Xclkbuf_5_29__f_clk clknet_2_3_0_clk VGND VGND VPWR VPWR clknet_5_29__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_29835_ net213 _01570_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[1\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23629__246 clknet_1_0__leaf__10181_ VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_128_3559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16800_ _04646_ VGND VGND VPWR VPWR _01644_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_206_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17780_ _05177_ VGND VGND VPWR VPWR _05178_ sky130_fd_sc_hd__clkbuf_4
X_29766_ net1112 _01501_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[20\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_54_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14992_ _13384_ _13319_ _13537_ _13539_ VGND VGND VPWR VPWR _13540_ sky130_fd_sc_hd__a211o_1
X_26978_ _11835_ _11866_ VGND VGND VPWR VPWR _11873_ sky130_fd_sc_hd__and2_1
X_16731_ _14195_ net3827 _04575_ VGND VGND VPWR VPWR _04610_ sky130_fd_sc_hd__mux2_1
X_28717_ _12857_ VGND VGND VPWR VPWR _04149_ sky130_fd_sc_hd__clkbuf_1
X_25929_ net1862 _11275_ _11273_ _11284_ VGND VGND VPWR VPWR _02934_ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_221_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29697_ net1043 _01432_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[23\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_50_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19450_ datamem.data_ram\[42\]\[16\] _06728_ _06726_ datamem.data_ram\[47\]\[16\]
+ _06745_ VGND VGND VPWR VPWR _06746_ sky130_fd_sc_hd__o221a_1
XFILLER_0_72_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16662_ _04573_ VGND VGND VPWR VPWR _01709_ sky130_fd_sc_hd__clkbuf_1
X_28648_ _12747_ net2406 net71 VGND VGND VPWR VPWR _12821_ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18401_ _05754_ _05764_ _05693_ VGND VGND VPWR VPWR _05765_ sky130_fd_sc_hd__mux2_1
XFILLER_0_213_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15613_ net2274 _13244_ _14114_ VGND VGND VPWR VPWR _14115_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19381_ _06676_ VGND VGND VPWR VPWR _06677_ sky130_fd_sc_hd__clkbuf_16
X_28579_ _12764_ net2249 _12777_ VGND VGND VPWR VPWR _12784_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16593_ _04536_ VGND VGND VPWR VPWR _01749_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18332_ _05696_ VGND VGND VPWR VPWR _05697_ sky130_fd_sc_hd__clkbuf_4
X_30610_ clknet_leaf_218_clk _02345_ VGND VGND VPWR VPWR datamem.data_ram\[52\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_15544_ _13767_ _13488_ _13401_ _13477_ _13672_ VGND VGND VPWR VPWR _14070_ sky130_fd_sc_hd__o32a_1
XFILLER_0_56_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31590_ clknet_leaf_51_clk net1245 VGND VGND VPWR VPWR rvcpu.dp.plmw.PCPlus4W\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_189_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18263_ _05625_ _05457_ _05461_ _05627_ VGND VGND VPWR VPWR _05628_ sky130_fd_sc_hd__o22a_1
X_30541_ clknet_leaf_143_clk _02276_ VGND VGND VPWR VPWR datamem.data_ram\[55\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_15475_ _13372_ _13867_ VGND VGND VPWR VPWR _14004_ sky130_fd_sc_hd__and2_1
XFILLER_0_170_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17214_ _14133_ net3123 _04865_ VGND VGND VPWR VPWR _04867_ sky130_fd_sc_hd__mux2_1
X_18194_ _05290_ _05298_ _05558_ _05288_ VGND VGND VPWR VPWR _05559_ sky130_fd_sc_hd__o31ai_2
X_30472_ net150 _02207_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[19\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32211_ clknet_leaf_242_clk _03633_ VGND VGND VPWR VPWR datamem.data_ram\[36\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_17145_ _04830_ VGND VGND VPWR VPWR _01467_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold707 datamem.data_ram\[1\]\[4\] VGND VGND VPWR VPWR net1857 sky130_fd_sc_hd__dlygate4sd3_1
Xhold718 rvcpu.dp.rf.reg_file_arr\[1\]\[30\] VGND VGND VPWR VPWR net1868 sky130_fd_sc_hd__dlygate4sd3_1
X_32142_ clknet_leaf_276_clk _03564_ VGND VGND VPWR VPWR datamem.data_ram\[39\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_17076_ _14127_ net3270 _04793_ VGND VGND VPWR VPWR _04794_ sky130_fd_sc_hd__mux2_1
Xhold729 rvcpu.dp.rf.reg_file_arr\[1\]\[6\] VGND VGND VPWR VPWR net1879 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24009__542 clknet_1_1__leaf__10241_ VGND VGND VPWR VPWR net668 sky130_fd_sc_hd__inv_2
X_16027_ _14353_ VGND VGND VPWR VPWR _02008_ sky130_fd_sc_hd__clkbuf_1
X_32073_ clknet_leaf_114_clk _03495_ VGND VGND VPWR VPWR datamem.data_ram\[33\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_209_422 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31024_ clknet_leaf_59_clk _02759_ VGND VGND VPWR VPWR datamem.data_ram\[40\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2108 datamem.data_ram\[48\]\[16\] VGND VGND VPWR VPWR net3258 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2119 datamem.data_ram\[57\]\[21\] VGND VGND VPWR VPWR net3269 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1407 rvcpu.dp.rf.reg_file_arr\[21\]\[25\] VGND VGND VPWR VPWR net2557 sky130_fd_sc_hd__dlygate4sd3_1
X_17978_ rvcpu.dp.plde.RD1E\[6\] _05267_ _05271_ _13259_ _05348_ VGND VGND VPWR VPWR
+ _05349_ sky130_fd_sc_hd__a221o_4
XPHY_EDGE_ROW_127_Right_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1418 rvcpu.dp.rf.reg_file_arr\[4\]\[5\] VGND VGND VPWR VPWR net2568 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_204_5383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1429 rvcpu.dp.rf.reg_file_arr\[23\]\[19\] VGND VGND VPWR VPWR net2579 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_204_5394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19717_ datamem.data_ram\[29\]\[0\] _06970_ _07009_ _07012_ VGND VGND VPWR VPWR _07013_
+ sky130_fd_sc_hd__a211o_1
X_16929_ net2874 _14480_ _04706_ VGND VGND VPWR VPWR _04715_ sky130_fd_sc_hd__mux2_1
X_32975_ clknet_leaf_140_clk _04397_ VGND VGND VPWR VPWR datamem.data_ram\[63\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19648_ _06639_ VGND VGND VPWR VPWR _06944_ sky130_fd_sc_hd__buf_6
X_31926_ _04439_ net119 VGND VGND VPWR VPWR datamem.rd_data_mem\[31\] sky130_fd_sc_hd__dlxtn_1
XTAP_TAPCELL_ROW_217_5700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_196_5195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_217_5711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31857_ clknet_leaf_124_clk _03311_ VGND VGND VPWR VPWR datamem.data_ram\[62\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_19579_ _06864_ _06866_ _06869_ _06874_ VGND VGND VPWR VPWR _06875_ sky130_fd_sc_hd__a31o_1
X_21610_ rvcpu.dp.rf.reg_file_arr\[12\]\[11\] rvcpu.dp.rf.reg_file_arr\[13\]\[11\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[11\] rvcpu.dp.rf.reg_file_arr\[15\]\[11\] _08696_
+ _08568_ VGND VGND VPWR VPWR _08861_ sky130_fd_sc_hd__mux4_1
XFILLER_0_47_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_213_5608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30808_ clknet_leaf_149_clk _02543_ VGND VGND VPWR VPWR datamem.data_ram\[45\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_213_5619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22590_ _09476_ _09739_ _09741_ _09474_ VGND VGND VPWR VPWR _09742_ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31788_ clknet_leaf_53_clk _03242_ VGND VGND VPWR VPWR datamem.data_ram\[8\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_192_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21541_ _08786_ _08790_ _08794_ _08625_ VGND VGND VPWR VPWR _01036_ sky130_fd_sc_hd__o31a_1
X_30739_ clknet_leaf_195_clk _02474_ VGND VGND VPWR VPWR datamem.data_ram\[47\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24260_ _10302_ VGND VGND VPWR VPWR _02247_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_209_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21472_ _08515_ _08728_ _08513_ VGND VGND VPWR VPWR _08729_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_117_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32409_ clknet_leaf_231_clk _03831_ VGND VGND VPWR VPWR datamem.data_ram\[28\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_20423_ datamem.data_ram\[7\]\[12\] _06706_ _07230_ datamem.data_ram\[4\]\[12\] VGND
+ VGND VPWR VPWR _07715_ sky130_fd_sc_hd__o22a_1
XFILLER_0_16_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_168_4530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20354_ _07610_ _07621_ _07645_ VGND VGND VPWR VPWR _07646_ sky130_fd_sc_hd__o21ai_2
Xclkload150 clknet_leaf_272_clk VGND VGND VPWR VPWR clkload150/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_222_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload161 clknet_leaf_180_clk VGND VGND VPWR VPWR clkload161/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload172 clknet_leaf_215_clk VGND VGND VPWR VPWR clkload172/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_105_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload183 clknet_leaf_216_clk VGND VGND VPWR VPWR clkload183/Y sky130_fd_sc_hd__clkinv_4
X_27950_ _12427_ VGND VGND VPWR VPWR _03812_ sky130_fd_sc_hd__clkbuf_1
X_23073_ _10098_ VGND VGND VPWR VPWR _01264_ sky130_fd_sc_hd__clkbuf_1
Xclkload194 clknet_leaf_182_clk VGND VGND VPWR VPWR clkload194/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_222_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_164_4427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20285_ datamem.data_ram\[27\]\[19\] _06739_ _07577_ _06967_ VGND VGND VPWR VPWR
+ _07578_ sky130_fd_sc_hd__o211a_1
XFILLER_0_178_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_164_4438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26901_ _10057_ VGND VGND VPWR VPWR _11825_ sky130_fd_sc_hd__clkbuf_4
X_22024_ _09249_ VGND VGND VPWR VPWR _01064_ sky130_fd_sc_hd__clkbuf_1
X_27881_ _12389_ VGND VGND VPWR VPWR _03781_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_216_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold12 rvcpu.dp.plde.PCPlus4E\[20\] VGND VGND VPWR VPWR net1162 sky130_fd_sc_hd__dlygate4sd3_1
X_29620_ net974 _01355_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[25\]\[23\] sky130_fd_sc_hd__dfxtp_1
Xhold2620 rvcpu.dp.rf.reg_file_arr\[28\]\[20\] VGND VGND VPWR VPWR net3770 sky130_fd_sc_hd__dlygate4sd3_1
X_26832_ _11781_ net1400 _11773_ _11782_ VGND VGND VPWR VPWR _03339_ sky130_fd_sc_hd__a31o_1
Xhold23 rvcpu.dp.plem.PCPlus4M\[28\] VGND VGND VPWR VPWR net1173 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2631 datamem.data_ram\[13\]\[10\] VGND VGND VPWR VPWR net3781 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2642 datamem.data_ram\[44\]\[12\] VGND VGND VPWR VPWR net3792 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 rvcpu.dp.plem.lAuiPCM\[18\] VGND VGND VPWR VPWR net1184 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2653 datamem.data_ram\[29\]\[12\] VGND VGND VPWR VPWR net3803 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold45 rvcpu.dp.plem.PCPlus4M\[25\] VGND VGND VPWR VPWR net1195 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 rvcpu.dp.plem.lAuiPCM\[3\] VGND VGND VPWR VPWR net1206 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2664 datamem.data_ram\[32\]\[18\] VGND VGND VPWR VPWR net3814 sky130_fd_sc_hd__dlygate4sd3_1
X_22990__696 clknet_1_0__leaf__10084_ VGND VGND VPWR VPWR net822 sky130_fd_sc_hd__inv_2
XFILLER_0_215_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold67 rvcpu.dp.plde.PCPlus4E\[28\] VGND VGND VPWR VPWR net1217 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1930 datamem.data_ram\[33\]\[16\] VGND VGND VPWR VPWR net3080 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2675 datamem.data_ram\[45\]\[27\] VGND VGND VPWR VPWR net3825 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_67_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29551_ net905 _01286_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[27\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_26763_ _11735_ net1745 _11737_ _11741_ VGND VGND VPWR VPWR _03311_ sky130_fd_sc_hd__a31o_1
Xhold78 rvcpu.dp.plem.lAuiPCM\[12\] VGND VGND VPWR VPWR net1228 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2686 datamem.data_ram\[27\]\[18\] VGND VGND VPWR VPWR net3836 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1941 datamem.data_ram\[5\]\[27\] VGND VGND VPWR VPWR net3091 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1952 datamem.data_ram\[10\]\[17\] VGND VGND VPWR VPWR net3102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2697 datamem.data_ram\[54\]\[28\] VGND VGND VPWR VPWR net3847 sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 rvcpu.dp.plde.PCPlus4E\[12\] VGND VGND VPWR VPWR net1239 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_123_3445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1963 rvcpu.dp.rf.reg_file_arr\[21\]\[19\] VGND VGND VPWR VPWR net3113 sky130_fd_sc_hd__dlygate4sd3_1
X_28502_ _12736_ VGND VGND VPWR VPWR _04055_ sky130_fd_sc_hd__clkbuf_1
Xhold1974 rvcpu.dp.rf.reg_file_arr\[27\]\[19\] VGND VGND VPWR VPWR net3124 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_123_3456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25714_ _11130_ VGND VGND VPWR VPWR _02873_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22926_ _10058_ _10053_ VGND VGND VPWR VPWR _10059_ sky130_fd_sc_hd__and2_1
Xhold1985 datamem.data_ram\[34\]\[18\] VGND VGND VPWR VPWR net3135 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f__10263_ clknet_0__10263_ VGND VGND VPWR VPWR clknet_1_1__leaf__10263_
+ sky130_fd_sc_hd__clkbuf_16
X_29482_ net844 _01217_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[2\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_26694_ _11700_ net1831 _11693_ _11701_ VGND VGND VPWR VPWR _03282_ sky130_fd_sc_hd__a31o_1
Xhold1996 datamem.data_ram\[59\]\[28\] VGND VGND VPWR VPWR net3146 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28433_ _09317_ VGND VGND VPWR VPWR _12696_ sky130_fd_sc_hd__clkbuf_2
X_25645_ _11085_ net1813 _11077_ _11092_ VGND VGND VPWR VPWR _02842_ sky130_fd_sc_hd__a31o_1
XFILLER_0_211_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22857_ _09516_ _09991_ _09993_ _09523_ VGND VGND VPWR VPWR _09994_ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__10194_ clknet_0__10194_ VGND VGND VPWR VPWR clknet_1_1__leaf__10194_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_156_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26510__62 clknet_1_0__leaf__11602_ VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__inv_2
X_21808_ rvcpu.dp.rf.reg_file_arr\[0\]\[22\] rvcpu.dp.rf.reg_file_arr\[1\]\[22\] rvcpu.dp.rf.reg_file_arr\[2\]\[22\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[22\] _08810_ _08811_ VGND VGND VPWR VPWR _09048_
+ sky130_fd_sc_hd__mux4_1
X_28364_ _12460_ net3972 net95 VGND VGND VPWR VPWR _12657_ sky130_fd_sc_hd__mux2_1
X_25576_ _10416_ _11042_ VGND VGND VPWR VPWR _11049_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_26_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22788_ rvcpu.dp.rf.reg_file_arr\[8\]\[25\] rvcpu.dp.rf.reg_file_arr\[10\]\[25\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[25\] rvcpu.dp.rf.reg_file_arr\[11\]\[25\] _09443_
+ _09453_ VGND VGND VPWR VPWR _09929_ sky130_fd_sc_hd__mux4_1
XFILLER_0_213_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27315_ _12061_ net1792 _12065_ _12072_ VGND VGND VPWR VPWR _03532_ sky130_fd_sc_hd__a31o_1
XFILLER_0_54_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24527_ _10390_ datamem.data_ram\[52\]\[10\] _10456_ VGND VGND VPWR VPWR _10459_
+ sky130_fd_sc_hd__mux2_1
X_28295_ _12443_ net3127 _12613_ VGND VGND VPWR VPWR _12620_ sky130_fd_sc_hd__mux2_1
X_21739_ rvcpu.dp.rf.reg_file_arr\[0\]\[18\] rvcpu.dp.rf.reg_file_arr\[1\]\[18\] rvcpu.dp.rf.reg_file_arr\[2\]\[18\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[18\] _08566_ _08569_ VGND VGND VPWR VPWR _08983_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_94_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15260_ _13320_ _13434_ VGND VGND VPWR VPWR _13800_ sky130_fd_sc_hd__or2_1
X_27246_ _11946_ _12031_ VGND VGND VPWR VPWR _12037_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_97_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24458_ _10072_ VGND VGND VPWR VPWR _10418_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_152_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15191_ _13336_ _13703_ _13581_ VGND VGND VPWR VPWR _13734_ sky130_fd_sc_hd__a21oi_1
X_27177_ _09226_ _11112_ _11898_ VGND VGND VPWR VPWR _11996_ sky130_fd_sc_hd__and3_1
XFILLER_0_151_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_229_Right_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24389_ _10373_ VGND VGND VPWR VPWR _02305_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_9 _06594_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26128_ net1761 _11397_ VGND VGND VPWR VPWR _11400_ sky130_fd_sc_hd__and2_1
XFILLER_0_105_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26059_ _11353_ net1826 _11350_ _11358_ VGND VGND VPWR VPWR _02990_ sky130_fd_sc_hd__a31o_1
X_18950_ _05275_ _05733_ _06285_ _06287_ VGND VGND VPWR VPWR _06288_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_56_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23863__425 clknet_1_1__leaf__10220_ VGND VGND VPWR VPWR net551 sky130_fd_sc_hd__inv_2
XFILLER_0_120_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17901_ rvcpu.dp.plde.RD1E\[31\] _05267_ _05271_ _13172_ _05273_ VGND VGND VPWR VPWR
+ _05274_ sky130_fd_sc_hd__a221o_1
XFILLER_0_30_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18881_ _05623_ _06212_ _06214_ _06223_ VGND VGND VPWR VPWR _06224_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_52_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17832_ rvcpu.dp.plem.ALUResultM\[22\] _05215_ _05177_ VGND VGND VPWR VPWR _05216_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29818_ net196 _01553_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[1\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17763_ _05156_ _05158_ _05159_ _05160_ VGND VGND VPWR VPWR _05161_ sky130_fd_sc_hd__and4bb_4
X_14975_ rvcpu.dp.pcreg.q\[5\] _13322_ VGND VGND VPWR VPWR _13523_ sky130_fd_sc_hd__nor2_4
X_29749_ net1095 _01484_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[21\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_221_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19502_ _06713_ _06749_ _06773_ _06795_ _06797_ VGND VGND VPWR VPWR _06798_ sky130_fd_sc_hd__a32o_1
XFILLER_0_117_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16714_ _04601_ VGND VGND VPWR VPWR _01685_ sky130_fd_sc_hd__clkbuf_1
X_32760_ clknet_leaf_177_clk _04182_ VGND VGND VPWR VPWR datamem.data_ram\[15\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_17694_ _05121_ VGND VGND VPWR VPWR _01193_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24039__568 clknet_1_0__leaf__10245_ VGND VGND VPWR VPWR net694 sky130_fd_sc_hd__inv_2
X_31711_ clknet_leaf_31_clk _03169_ VGND VGND VPWR VPWR rvcpu.dp.pcreg.q\[29\] sky130_fd_sc_hd__dfxtp_1
X_19433_ _06631_ VGND VGND VPWR VPWR _06729_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_57_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16645_ _14177_ net2494 _04562_ VGND VGND VPWR VPWR _04565_ sky130_fd_sc_hd__mux2_1
X_32691_ clknet_leaf_251_clk _04113_ VGND VGND VPWR VPWR datamem.data_ram\[18\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_201_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_201_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31642_ clknet_leaf_29_clk net1220 VGND VGND VPWR VPWR rvcpu.dp.plmw.lAuiPCW\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_19364_ net122 _06615_ VGND VGND VPWR VPWR _06660_ sky130_fd_sc_hd__nand2_8
XFILLER_0_69_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_191_5070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16576_ _14177_ net4195 _04525_ VGND VGND VPWR VPWR _04528_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_191_5081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18315_ _05342_ _05349_ _05358_ _05679_ _05664_ _05669_ VGND VGND VPWR VPWR _05680_
+ sky130_fd_sc_hd__mux4_2
X_15527_ _13665_ _13451_ _13985_ VGND VGND VPWR VPWR _14053_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_174_549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31573_ clknet_leaf_71_clk datamem.rd_data_mem\[23\] VGND VGND VPWR VPWR rvcpu.dp.plmw.ReadDataW\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_19295_ net1 VGND VGND VPWR VPWR _06591_ sky130_fd_sc_hd__buf_8
XFILLER_0_127_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_218_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18246_ _05610_ _05330_ _05438_ _05323_ _05437_ VGND VGND VPWR VPWR _05611_ sky130_fd_sc_hd__o32a_1
XFILLER_0_127_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30524_ clknet_leaf_195_clk _02259_ VGND VGND VPWR VPWR datamem.data_ram\[56\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_15458_ _13682_ _13573_ _13321_ _13402_ VGND VGND VPWR VPWR _13988_ sky130_fd_sc_hd__or4_1
XFILLER_0_155_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18177_ _05539_ _05540_ VGND VGND VPWR VPWR _05542_ sky130_fd_sc_hd__and2_1
X_30455_ net133 _02190_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[19\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_15389_ _13496_ _13443_ VGND VGND VPWR VPWR _13922_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold504 datamem.data_ram\[63\]\[4\] VGND VGND VPWR VPWR net1654 sky130_fd_sc_hd__dlygate4sd3_1
X_17128_ _14183_ net3918 _04815_ VGND VGND VPWR VPWR _04821_ sky130_fd_sc_hd__mux2_1
Xhold515 datamem.data_ram\[57\]\[3\] VGND VGND VPWR VPWR net1665 sky130_fd_sc_hd__dlygate4sd3_1
X_30386_ clknet_leaf_269_clk _02121_ VGND VGND VPWR VPWR datamem.data_ram\[58\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold526 rvcpu.dp.plfd.PCPlus4D\[13\] VGND VGND VPWR VPWR net1676 sky130_fd_sc_hd__dlygate4sd3_1
Xhold537 datamem.data_ram\[25\]\[5\] VGND VGND VPWR VPWR net1687 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_229_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold548 datamem.data_ram\[58\]\[2\] VGND VGND VPWR VPWR net1698 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32125_ clknet_leaf_234_clk _03547_ VGND VGND VPWR VPWR datamem.data_ram\[7\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold559 datamem.data_ram\[61\]\[5\] VGND VGND VPWR VPWR net1709 sky130_fd_sc_hd__dlygate4sd3_1
X_17059_ _04784_ VGND VGND VPWR VPWR _01507_ sky130_fd_sc_hd__clkbuf_1
X_23039__740 clknet_1_1__leaf__10089_ VGND VGND VPWR VPWR net866 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_206_5434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_206_5445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32056_ clknet_leaf_131_clk _03478_ VGND VGND VPWR VPWR datamem.data_ram\[30\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_20070_ _06678_ _07361_ _07363_ _06750_ VGND VGND VPWR VPWR _07364_ sky130_fd_sc_hd__a31o_1
Xclkbuf_5_12__f_clk clknet_2_1_0_clk VGND VGND VPWR VPWR clknet_5_12__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_148_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31007_ clknet_leaf_164_clk _02742_ VGND VGND VPWR VPWR datamem.data_ram\[11\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1204 rvcpu.dp.rf.reg_file_arr\[30\]\[25\] VGND VGND VPWR VPWR net2354 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_198_5246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1215 datamem.data_ram\[7\]\[30\] VGND VGND VPWR VPWR net2365 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_198_5257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1226 datamem.data_ram\[59\]\[15\] VGND VGND VPWR VPWR net2376 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1237 rvcpu.dp.rf.reg_file_arr\[23\]\[31\] VGND VGND VPWR VPWR net2387 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1248 rvcpu.dp.rf.reg_file_arr\[26\]\[0\] VGND VGND VPWR VPWR net2398 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1259 rvcpu.dp.rf.reg_file_arr\[19\]\[9\] VGND VGND VPWR VPWR net2409 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_164_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20972_ datamem.data_ram\[33\]\[15\] _06945_ _08260_ _06598_ VGND VGND VPWR VPWR
+ _08261_ sky130_fd_sc_hd__a211o_1
X_32958_ clknet_leaf_98_clk _04380_ VGND VGND VPWR VPWR datamem.data_ram\[6\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22711_ _09422_ _09855_ _09472_ VGND VGND VPWR VPWR _09856_ sky130_fd_sc_hd__o21ai_1
X_31909_ _04420_ net121 VGND VGND VPWR VPWR datamem.rd_data_mem\[14\] sky130_fd_sc_hd__dlxtn_1
XFILLER_0_95_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_177_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32889_ clknet_leaf_158_clk _04311_ VGND VGND VPWR VPWR datamem.data_ram\[10\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_157_4253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_4264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25430_ _10971_ VGND VGND VPWR VPWR _02748_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_193_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22642_ _09622_ _09787_ _09790_ VGND VGND VPWR VPWR _09791_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_157_4275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_177_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25361_ _10876_ net1411 _10920_ _10929_ VGND VGND VPWR VPWR _02721_ sky130_fd_sc_hd__a31o_1
X_22573_ _09725_ VGND VGND VPWR VPWR _01137_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27100_ _11946_ _11941_ VGND VGND VPWR VPWR _11947_ sky130_fd_sc_hd__and2_1
X_24312_ _10331_ VGND VGND VPWR VPWR _02270_ sky130_fd_sc_hd__clkbuf_1
X_28080_ _12504_ VGND VGND VPWR VPWR _03865_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21524_ _08535_ VGND VGND VPWR VPWR _08778_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_69_1034 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25292_ _10754_ net3727 _10887_ VGND VGND VPWR VPWR _10889_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27031_ _11752_ VGND VGND VPWR VPWR _11904_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_133_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24243_ _09282_ net3271 _10288_ VGND VGND VPWR VPWR _10293_ sky130_fd_sc_hd__mux2_1
X_21455_ rvcpu.dp.rf.reg_file_arr\[4\]\[4\] rvcpu.dp.rf.reg_file_arr\[5\]\[4\] rvcpu.dp.rf.reg_file_arr\[6\]\[4\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[4\] _08551_ _08555_ VGND VGND VPWR VPWR _08713_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_116_3271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23274__919 clknet_1_0__leaf__10129_ VGND VGND VPWR VPWR net1045 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_116_3282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20406_ datamem.data_ram\[46\]\[12\] _06744_ _06690_ datamem.data_ram\[42\]\[12\]
+ _07697_ VGND VGND VPWR VPWR _07698_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_92_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21386_ _08547_ _08644_ _08646_ _08575_ VGND VGND VPWR VPWR _08647_ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_187_4972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_187_4983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_283_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_283_clk
+ sky130_fd_sc_hd__clkbuf_8
X_20337_ datamem.data_ram\[32\]\[4\] _06990_ _07628_ _06967_ VGND VGND VPWR VPWR _07629_
+ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_187_4994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput13 net13 VGND VGND VPWR VPWR Instr[1] sky130_fd_sc_hd__buf_2
Xoutput24 net24 VGND VGND VPWR VPWR Instr[2] sky130_fd_sc_hd__buf_2
X_28982_ _13000_ VGND VGND VPWR VPWR _04271_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__11602_ _11602_ VGND VGND VPWR VPWR clknet_0__11602_ sky130_fd_sc_hd__clkbuf_16
X_27933_ _12418_ VGND VGND VPWR VPWR _03804_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20268_ _06967_ _07558_ _07560_ VGND VGND VPWR VPWR _07561_ sky130_fd_sc_hd__and3_1
Xhold3140 rvcpu.dp.rf.reg_file_arr\[18\]\[2\] VGND VGND VPWR VPWR net4290 sky130_fd_sc_hd__dlygate4sd3_1
X_22007_ _09235_ VGND VGND VPWR VPWR _09236_ sky130_fd_sc_hd__clkbuf_2
Xhold3151 rvcpu.dp.rf.reg_file_arr\[13\]\[14\] VGND VGND VPWR VPWR net4301 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3162 rvcpu.dp.rf.reg_file_arr\[24\]\[31\] VGND VGND VPWR VPWR net4312 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_125_3507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27864_ _12380_ VGND VGND VPWR VPWR _03773_ sky130_fd_sc_hd__clkbuf_1
Xhold3173 datamem.data_ram\[30\]\[28\] VGND VGND VPWR VPWR net4323 sky130_fd_sc_hd__dlygate4sd3_1
X_20199_ datamem.data_ram\[34\]\[11\] _07023_ _07488_ _07491_ VGND VGND VPWR VPWR
+ _07492_ sky130_fd_sc_hd__o211a_1
Xhold3184 datamem.data_ram\[41\]\[28\] VGND VGND VPWR VPWR net4334 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3195 datamem.data_ram\[24\]\[22\] VGND VGND VPWR VPWR net4345 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2450 datamem.data_ram\[0\]\[9\] VGND VGND VPWR VPWR net3600 sky130_fd_sc_hd__dlygate4sd3_1
X_26815_ _07808_ _11725_ _11494_ VGND VGND VPWR VPWR _11772_ sky130_fd_sc_hd__or3_1
Xhold2461 datamem.data_ram\[49\]\[16\] VGND VGND VPWR VPWR net3611 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_3990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29603_ net957 _01338_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[25\]\[6\] sky130_fd_sc_hd__dfxtp_1
Xhold2472 datamem.data_ram\[32\]\[14\] VGND VGND VPWR VPWR net3622 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27795_ _12339_ VGND VGND VPWR VPWR _03745_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2483 rvcpu.dp.rf.reg_file_arr\[2\]\[12\] VGND VGND VPWR VPWR net3633 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2494 rvcpu.dp.rf.reg_file_arr\[19\]\[18\] VGND VGND VPWR VPWR net3644 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1760 rvcpu.dp.rf.reg_file_arr\[31\]\[8\] VGND VGND VPWR VPWR net2910 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29534_ net888 _01269_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[27\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_26746_ _11645_ _11726_ VGND VGND VPWR VPWR _11731_ sky130_fd_sc_hd__and2_1
X_14760_ rvcpu.dp.pcreg.q\[7\] VGND VGND VPWR VPWR _13313_ sky130_fd_sc_hd__clkbuf_4
Xhold1771 datamem.data_ram\[30\]\[18\] VGND VGND VPWR VPWR net2921 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_86_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23958_ _09244_ net4222 _10229_ VGND VGND VPWR VPWR _10233_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1782 datamem.data_ram\[26\]\[31\] VGND VGND VPWR VPWR net2932 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_86_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1793 rvcpu.dp.rf.reg_file_arr\[0\]\[15\] VGND VGND VPWR VPWR net2943 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22909_ _09217_ _09262_ _09220_ VGND VGND VPWR VPWR _10043_ sky130_fd_sc_hd__a21oi_4
Xclkbuf_1_1__f__10246_ clknet_0__10246_ VGND VGND VPWR VPWR clknet_1_1__leaf__10246_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_98_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29465_ net827 _01200_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[2\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_26677_ _11672_ _11677_ VGND VGND VPWR VPWR _11691_ sky130_fd_sc_hd__and2_1
X_14691_ rvcpu.dp.plmw.ALUResultW\[8\] rvcpu.dp.plmw.ReadDataW\[8\] rvcpu.dp.plmw.PCPlus4W\[8\]
+ rvcpu.dp.plmw.lAuiPCW\[8\] _13169_ _13171_ VGND VGND VPWR VPWR _13253_ sky130_fd_sc_hd__mux4_2
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16430_ _14581_ VGND VGND VPWR VPWR _01825_ sky130_fd_sc_hd__clkbuf_1
X_28416_ _12460_ net3736 _12678_ VGND VGND VPWR VPWR _12685_ sky130_fd_sc_hd__mux2_1
X_25628_ _10057_ VGND VGND VPWR VPWR _11081_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_168_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_224_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29396_ clknet_leaf_1_clk _01131_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD2E\[7\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__10177_ clknet_0__10177_ VGND VGND VPWR VPWR clknet_1_1__leaf__10177_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_156_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_706 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28347_ _12443_ net2530 _12641_ VGND VGND VPWR VPWR _12648_ sky130_fd_sc_hd__mux2_1
X_16361_ net2225 _14459_ _14536_ VGND VGND VPWR VPWR _14545_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25559_ _10766_ net2690 _11030_ VGND VGND VPWR VPWR _11038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18100_ rvcpu.dp.plem.ALUResultM\[21\] _05339_ _05340_ _13212_ VGND VGND VPWR VPWR
+ _05468_ sky130_fd_sc_hd__o22a_1
X_15312_ _13823_ _13420_ _13693_ _13848_ VGND VGND VPWR VPWR _13849_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_45_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19080_ _06404_ rvcpu.dp.plde.ImmExtE\[8\] _06355_ VGND VGND VPWR VPWR _06405_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16292_ _14508_ VGND VGND VPWR VPWR _01890_ sky130_fd_sc_hd__clkbuf_1
X_28278_ _12610_ VGND VGND VPWR VPWR _03957_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_227_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23672__269 clknet_1_0__leaf__10193_ VGND VGND VPWR VPWR net395 sky130_fd_sc_hd__inv_2
X_18031_ _05378_ _05400_ _05374_ VGND VGND VPWR VPWR _05401_ sky130_fd_sc_hd__a21bo_1
X_15243_ _13352_ _13779_ _13781_ _13782_ VGND VGND VPWR VPWR _13783_ sky130_fd_sc_hd__a31o_1
X_27229_ _12022_ net1438 _12018_ _12026_ VGND VGND VPWR VPWR _03492_ sky130_fd_sc_hd__a31o_1
XFILLER_0_83_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30240_ net594 _01975_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[7\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_15174_ _13320_ _13349_ VGND VGND VPWR VPWR _13717_ sky130_fd_sc_hd__nand2_2
XFILLER_0_50_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_205_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_274_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_274_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30171_ net533 _01906_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[0\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_19982_ _07253_ _07275_ VGND VGND VPWR VPWR _07276_ sky130_fd_sc_hd__nor2_2
X_18933_ _06217_ _06271_ _05707_ VGND VGND VPWR VPWR _06272_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18864_ _05619_ _05655_ _06207_ VGND VGND VPWR VPWR _06208_ sky130_fd_sc_hd__or3_1
X_24186__26 clknet_1_0__leaf__10266_ VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_201_5320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_201_5331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17815_ _05204_ VGND VGND VPWR VPWR rvcpu.dp.SrcBFW_Mux.y\[28\] sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_118_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18795_ _05706_ _06078_ _06142_ VGND VGND VPWR VPWR _06143_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32812_ clknet_leaf_257_clk _04234_ VGND VGND VPWR VPWR datamem.data_ram\[13\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_17746_ _05148_ VGND VGND VPWR VPWR _01168_ sky130_fd_sc_hd__clkbuf_1
X_14958_ _13296_ _13506_ VGND VGND VPWR VPWR _13507_ sky130_fd_sc_hd__nor2_2
XFILLER_0_168_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_193_5121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_193_5132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_221_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32743_ clknet_leaf_284_clk _04165_ VGND VGND VPWR VPWR datamem.data_ram\[16\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_17677_ net3120 _13265_ _05104_ VGND VGND VPWR VPWR _05112_ sky130_fd_sc_hd__mux2_1
X_14889_ _13325_ _13411_ _13440_ _13406_ VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__o31a_1
XFILLER_0_159_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16628_ _14160_ net3602 _04551_ VGND VGND VPWR VPWR _04556_ sky130_fd_sc_hd__mux2_1
X_19416_ _06594_ VGND VGND VPWR VPWR _06712_ sky130_fd_sc_hd__buf_4
XFILLER_0_202_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32674_ clknet_leaf_266_clk _04096_ VGND VGND VPWR VPWR datamem.data_ram\[18\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31625_ clknet_leaf_65_clk net1215 VGND VGND VPWR VPWR rvcpu.dp.plmw.lAuiPCW\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19347_ _06639_ _06642_ VGND VGND VPWR VPWR _06643_ sky130_fd_sc_hd__nand2_4
X_16559_ _14160_ net3235 _04514_ VGND VGND VPWR VPWR _04519_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_210_1060 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31556_ clknet_leaf_64_clk datamem.rd_data_mem\[6\] VGND VGND VPWR VPWR rvcpu.dp.plmw.ReadDataW\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_19278_ rvcpu.dp.plfd.InstrD\[14\] _06574_ _06576_ _06567_ VGND VGND VPWR VPWR _04448_
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_152_4150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18229_ _05353_ _05349_ VGND VGND VPWR VPWR _05594_ sky130_fd_sc_hd__or2b_1
X_30507_ clknet_leaf_174_clk _02242_ VGND VGND VPWR VPWR datamem.data_ram\[57\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31487_ clknet_leaf_48_clk rvcpu.dp.lAuiPCE\[13\] VGND VGND VPWR VPWR rvcpu.dp.plem.lAuiPCM\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21240_ datamem.data_ram\[52\]\[24\] datamem.data_ram\[52\]\[16\] VGND VGND VPWR
+ VPWR _08503_ sky130_fd_sc_hd__nand2_1
XFILLER_0_142_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30438_ net776 _02173_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[29\]\[17\] sky130_fd_sc_hd__dfxtp_1
Xhold301 datamem.data_ram\[50\]\[0\] VGND VGND VPWR VPWR net1451 sky130_fd_sc_hd__dlygate4sd3_1
Xhold312 datamem.data_ram\[59\]\[7\] VGND VGND VPWR VPWR net1462 sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 datamem.data_ram\[39\]\[1\] VGND VGND VPWR VPWR net1473 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__10266_ clknet_0__10266_ VGND VGND VPWR VPWR clknet_1_0__leaf__10266_
+ sky130_fd_sc_hd__clkbuf_16
Xhold334 datamem.data_ram\[4\]\[2\] VGND VGND VPWR VPWR net1484 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_265_clk clknet_5_19__leaf_clk VGND VGND VPWR VPWR clknet_leaf_265_clk
+ sky130_fd_sc_hd__clkbuf_8
X_21171_ _07859_ _08459_ _06598_ VGND VGND VPWR VPWR _08460_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_229_5990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold345 datamem.data_ram\[7\]\[2\] VGND VGND VPWR VPWR net1495 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30369_ net715 _02104_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[3\]\[20\] sky130_fd_sc_hd__dfxtp_1
Xhold356 datamem.data_ram\[3\]\[1\] VGND VGND VPWR VPWR net1506 sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 datamem.data_ram\[13\]\[3\] VGND VGND VPWR VPWR net1517 sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 datamem.data_ram\[24\]\[5\] VGND VGND VPWR VPWR net1528 sky130_fd_sc_hd__dlygate4sd3_1
X_32108_ clknet_leaf_116_clk _03530_ VGND VGND VPWR VPWR datamem.data_ram\[58\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_20122_ _07277_ _07322_ _07415_ _06583_ VGND VGND VPWR VPWR _07416_ sky130_fd_sc_hd__o22a_1
Xclkbuf_1_0__f__10197_ clknet_0__10197_ VGND VGND VPWR VPWR clknet_1_0__leaf__10197_
+ sky130_fd_sc_hd__clkbuf_16
Xhold389 datamem.data_ram\[20\]\[6\] VGND VGND VPWR VPWR net1539 sky130_fd_sc_hd__dlygate4sd3_1
X_23649__249 clknet_1_1__leaf__10181_ VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__inv_2
XFILLER_0_102_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_225_5887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_225_5898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32039_ clknet_leaf_132_clk _03461_ VGND VGND VPWR VPWR datamem.data_ram\[50\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_24930_ _10683_ VGND VGND VPWR VPWR _02536_ sky130_fd_sc_hd__clkbuf_1
X_20053_ datamem.data_ram\[35\]\[26\] _06729_ _07242_ datamem.data_ram\[33\]\[26\]
+ _07346_ VGND VGND VPWR VPWR _07347_ sky130_fd_sc_hd__o221a_1
XFILLER_0_102_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1001 datamem.data_ram\[35\]\[18\] VGND VGND VPWR VPWR net2151 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1012 rvcpu.dp.rf.reg_file_arr\[10\]\[2\] VGND VGND VPWR VPWR net2162 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_225_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1023 datamem.data_ram\[50\]\[23\] VGND VGND VPWR VPWR net2173 sky130_fd_sc_hd__dlygate4sd3_1
X_24861_ _10646_ VGND VGND VPWR VPWR _02504_ sky130_fd_sc_hd__clkbuf_1
Xhold1034 datamem.data_ram\[43\]\[31\] VGND VGND VPWR VPWR net2184 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1045 rvcpu.dp.rf.reg_file_arr\[4\]\[14\] VGND VGND VPWR VPWR net2195 sky130_fd_sc_hd__dlygate4sd3_1
X_26600_ _11618_ net1642 _11639_ _11647_ VGND VGND VPWR VPWR _03242_ sky130_fd_sc_hd__a31o_1
Xhold1056 datamem.data_ram\[63\]\[26\] VGND VGND VPWR VPWR net2206 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_159_4304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1067 datamem.data_ram\[47\]\[14\] VGND VGND VPWR VPWR net2217 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_1_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_4315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27580_ _12223_ VGND VGND VPWR VPWR _03646_ sky130_fd_sc_hd__clkbuf_1
X_24792_ _10608_ VGND VGND VPWR VPWR _02473_ sky130_fd_sc_hd__clkbuf_1
Xhold1078 rvcpu.dp.rf.reg_file_arr\[0\]\[5\] VGND VGND VPWR VPWR net2228 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_213_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1089 datamem.data_ram\[44\]\[9\] VGND VGND VPWR VPWR net2239 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__10200_ _10200_ VGND VGND VPWR VPWR clknet_0__10200_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_217_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_207 _09560_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26531_ _11607_ VGND VGND VPWR VPWR _11608_ sky130_fd_sc_hd__clkbuf_2
XANTENNA_218 _09813_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_229 _10072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_178_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20955_ datamem.data_ram\[48\]\[15\] _06933_ _06606_ VGND VGND VPWR VPWR _08244_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_36_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0__10131_ _10131_ VGND VGND VPWR VPWR clknet_0__10131_ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_81_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29250_ _13145_ VGND VGND VPWR VPWR _04394_ sky130_fd_sc_hd__clkbuf_1
X_26462_ net1900 _11573_ _11586_ _11570_ VGND VGND VPWR VPWR _03165_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_81_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20886_ datamem.data_ram\[63\]\[14\] _07831_ _08175_ _07821_ VGND VGND VPWR VPWR
+ _08176_ sky130_fd_sc_hd__o211a_1
X_28201_ _12568_ VGND VGND VPWR VPWR _03922_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25413_ _10962_ VGND VGND VPWR VPWR _02740_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_187_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29181_ _09247_ net3568 net63 VGND VGND VPWR VPWR _13108_ sky130_fd_sc_hd__mux2_1
X_22625_ _09534_ _09774_ VGND VGND VPWR VPWR _09775_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26393_ _13682_ _11329_ _11537_ _11534_ VGND VGND VPWR VPWR _03145_ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_3322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_3333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28132_ _12437_ net2996 _12528_ VGND VGND VPWR VPWR _12532_ sky130_fd_sc_hd__mux2_1
XFILLER_0_187_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25344_ _10043_ VGND VGND VPWR VPWR _10918_ sky130_fd_sc_hd__buf_2
XFILLER_0_10_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23591__212 clknet_1_1__leaf__10177_ VGND VGND VPWR VPWR net338 sky130_fd_sc_hd__inv_2
X_22556_ rvcpu.dp.rf.reg_file_arr\[24\]\[13\] rvcpu.dp.rf.reg_file_arr\[25\]\[13\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[13\] rvcpu.dp.rf.reg_file_arr\[27\]\[13\] _09393_
+ _09465_ VGND VGND VPWR VPWR _09709_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_101_Left_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_889 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21507_ _08760_ _08761_ _08743_ VGND VGND VPWR VPWR _08762_ sky130_fd_sc_hd__mux2_2
X_28063_ _12495_ VGND VGND VPWR VPWR _03857_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25275_ _10727_ net4050 _10878_ VGND VGND VPWR VPWR _10880_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22487_ rvcpu.dp.rf.reg_file_arr\[12\]\[9\] rvcpu.dp.rf.reg_file_arr\[13\]\[9\] rvcpu.dp.rf.reg_file_arr\[14\]\[9\]
+ rvcpu.dp.rf.reg_file_arr\[15\]\[9\] _09464_ _09467_ VGND VGND VPWR VPWR _09644_
+ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_40_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27014_ _11889_ net1751 _11885_ _11893_ VGND VGND VPWR VPWR _03410_ sky130_fd_sc_hd__a31o_1
XFILLER_0_133_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24226_ _09248_ net4139 _10279_ VGND VGND VPWR VPWR _10284_ sky130_fd_sc_hd__mux2_1
XFILLER_0_224_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21438_ rvcpu.dp.rf.reg_file_arr\[12\]\[3\] rvcpu.dp.rf.reg_file_arr\[13\]\[3\] rvcpu.dp.rf.reg_file_arr\[14\]\[3\]
+ rvcpu.dp.rf.reg_file_arr\[15\]\[3\] _08696_ _08568_ VGND VGND VPWR VPWR _08697_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_161_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_298 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_256_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_256_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_20_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21369_ rvcpu.dp.rf.reg_file_arr\[16\]\[1\] rvcpu.dp.rf.reg_file_arr\[17\]\[1\] rvcpu.dp.rf.reg_file_arr\[18\]\[1\]
+ rvcpu.dp.rf.reg_file_arr\[19\]\[1\] _08628_ _08629_ VGND VGND VPWR VPWR _08630_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_120_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28965_ _10057_ _12989_ VGND VGND VPWR VPWR _12991_ sky130_fd_sc_hd__and2_1
XFILLER_0_102_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24088_ _09288_ net3837 _10249_ VGND VGND VPWR VPWR _10256_ sky130_fd_sc_hd__mux2_1
Xhold890 rvcpu.dp.rf.reg_file_arr\[18\]\[5\] VGND VGND VPWR VPWR net2040 sky130_fd_sc_hd__dlygate4sd3_1
X_23708__302 clknet_1_1__leaf__10196_ VGND VGND VPWR VPWR net428 sky130_fd_sc_hd__inv_2
XFILLER_0_21_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15930_ net2326 _13254_ _14297_ VGND VGND VPWR VPWR _14301_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_88_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27916_ _12409_ VGND VGND VPWR VPWR _03796_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_194_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28896_ _12739_ net3781 net68 VGND VGND VPWR VPWR _12953_ sky130_fd_sc_hd__mux2_1
XFILLER_0_219_88 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_110_Left_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_216_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_144_3949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27847_ _09329_ VGND VGND VPWR VPWR _12371_ sky130_fd_sc_hd__clkbuf_2
X_15861_ net2198 _13257_ _14258_ VGND VGND VPWR VPWR _14263_ sky130_fd_sc_hd__mux2_1
XFILLER_0_216_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2280 datamem.data_ram\[59\]\[22\] VGND VGND VPWR VPWR net3430 sky130_fd_sc_hd__dlygate4sd3_1
X_17600_ _05071_ VGND VGND VPWR VPWR _01237_ sky130_fd_sc_hd__clkbuf_1
X_14812_ _13313_ rvcpu.dp.pcreg.q\[6\] VGND VGND VPWR VPWR _13365_ sky130_fd_sc_hd__and2_1
Xhold2291 datamem.data_ram\[61\]\[8\] VGND VGND VPWR VPWR net3441 sky130_fd_sc_hd__dlygate4sd3_1
X_18580_ _05669_ _05687_ _05938_ VGND VGND VPWR VPWR _05939_ sky130_fd_sc_hd__a21o_1
X_27778_ _12087_ net3172 _12326_ VGND VGND VPWR VPWR _12330_ sky130_fd_sc_hd__mux2_1
X_15792_ _14181_ net3274 _14221_ VGND VGND VPWR VPWR _14226_ sky130_fd_sc_hd__mux2_1
Xhold1590 datamem.data_ram\[15\]\[22\] VGND VGND VPWR VPWR net2740 sky130_fd_sc_hd__dlygate4sd3_1
X_17531_ _13251_ net3071 _05032_ VGND VGND VPWR VPWR _05035_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14743_ _13295_ VGND VGND VPWR VPWR _13296_ sky130_fd_sc_hd__buf_4
X_26729_ _11720_ VGND VGND VPWR VPWR _03298_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29517_ net879 _01252_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[28\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_197_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17462_ _04998_ VGND VGND VPWR VPWR _01310_ sky130_fd_sc_hd__clkbuf_1
X_29448_ net810 _01183_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[30\]\[19\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_103_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14674_ rvcpu.dp.plmw.ALUResultW\[12\] rvcpu.dp.plmw.ReadDataW\[12\] rvcpu.dp.plmw.PCPlus4W\[12\]
+ rvcpu.dp.plmw.lAuiPCW\[12\] _13168_ _13170_ VGND VGND VPWR VPWR _13240_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_103_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19201_ _06501_ _06510_ VGND VGND VPWR VPWR _06511_ sky130_fd_sc_hd__nand2_1
X_16413_ net2000 _14442_ _14572_ VGND VGND VPWR VPWR _14573_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_200_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29379_ clknet_leaf_139_clk _01114_ VGND VGND VPWR VPWR datamem.data_ram\[60\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17393_ _14175_ net3159 _04960_ VGND VGND VPWR VPWR _04962_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_82_Right_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19132_ rvcpu.dp.plde.ImmExtE\[15\] rvcpu.dp.plde.PCE\[15\] VGND VGND VPWR VPWR _06450_
+ sky130_fd_sc_hd__nand2_1
X_31410_ clknet_leaf_23_clk _03113_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCE\[27\] sky130_fd_sc_hd__dfxtp_1
X_23754__344 clknet_1_0__leaf__10200_ VGND VGND VPWR VPWR net470 sky130_fd_sc_hd__inv_2
XFILLER_0_229_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16344_ _14524_ VGND VGND VPWR VPWR _14536_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_183_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32390_ clknet_leaf_246_clk _03812_ VGND VGND VPWR VPWR datamem.data_ram\[29\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19063_ _06374_ _06376_ _06389_ _06379_ VGND VGND VPWR VPWR _06390_ sky130_fd_sc_hd__o211a_1
X_31341_ clknet_leaf_17_clk _03044_ VGND VGND VPWR VPWR rvcpu.dp.plde.Rs1E\[2\] sky130_fd_sc_hd__dfxtp_1
X_16275_ _14499_ VGND VGND VPWR VPWR _01898_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_180_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18014_ _05321_ rvcpu.dp.plde.ImmExtE\[1\] VGND VGND VPWR VPWR _05384_ sky130_fd_sc_hd__nand2_1
X_15226_ _13285_ VGND VGND VPWR VPWR _13767_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_120_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23869__431 clknet_1_0__leaf__10220_ VGND VGND VPWR VPWR net557 sky130_fd_sc_hd__inv_2
X_31272_ clknet_leaf_35_clk _02975_ VGND VGND VPWR VPWR rvcpu.c.ad.funct7b5 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_247_clk clknet_5_17__leaf_clk VGND VGND VPWR VPWR clknet_leaf_247_clk
+ sky130_fd_sc_hd__clkbuf_8
X_30223_ net577 _01958_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[7\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_15157_ _13410_ _13691_ _13695_ _13700_ VGND VGND VPWR VPWR _13701_ sky130_fd_sc_hd__o211a_1
XFILLER_0_164_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30154_ net516 _01889_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[0\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_15088_ _13389_ _13484_ VGND VGND VPWR VPWR _13634_ sky130_fd_sc_hd__nor2_2
X_19965_ datamem.data_ram\[14\]\[18\] _06763_ _06663_ datamem.data_ram\[13\]\[18\]
+ _07258_ VGND VGND VPWR VPWR _07259_ sky130_fd_sc_hd__o221a_1
XFILLER_0_120_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_91_Right_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18916_ _05707_ _06255_ _06109_ VGND VGND VPWR VPWR _06256_ sky130_fd_sc_hd__a21o_1
X_30085_ net447 _01820_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[11\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_19896_ _06698_ VGND VGND VPWR VPWR _07191_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_219_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18847_ _05494_ _06167_ _05563_ VGND VGND VPWR VPWR _06192_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_222_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_220_5773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_220_5784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18778_ _05990_ _05986_ _05989_ _06109_ VGND VGND VPWR VPWR _06127_ sky130_fd_sc_hd__o22a_1
XFILLER_0_222_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23460__109 clknet_1_1__leaf__10157_ VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__inv_2
XFILLER_0_54_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17729_ _05139_ VGND VGND VPWR VPWR _01176_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30987_ clknet_leaf_91_clk _02722_ VGND VGND VPWR VPWR datamem.data_ram\[39\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_19_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20740_ datamem.data_ram\[42\]\[6\] _07000_ _07137_ datamem.data_ram\[43\]\[6\] _06777_
+ VGND VGND VPWR VPWR _08030_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_154_4201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32726_ clknet_leaf_243_clk _04148_ VGND VGND VPWR VPWR datamem.data_ram\[16\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20671_ _06752_ _07956_ _07961_ _06594_ VGND VGND VPWR VPWR _07962_ sky130_fd_sc_hd__o31a_1
X_32657_ clknet_leaf_79_clk _04079_ VGND VGND VPWR VPWR datamem.data_ram\[19\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_23082__763 clknet_1_1__leaf__10091_ VGND VGND VPWR VPWR net889 sky130_fd_sc_hd__inv_2
XFILLER_0_162_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22410_ rvcpu.dp.rf.reg_file_arr\[12\]\[5\] rvcpu.dp.rf.reg_file_arr\[13\]\[5\] rvcpu.dp.rf.reg_file_arr\[14\]\[5\]
+ rvcpu.dp.rf.reg_file_arr\[15\]\[5\] _09478_ _09479_ VGND VGND VPWR VPWR _09571_
+ sky130_fd_sc_hd__mux4_1
X_31608_ clknet_leaf_26_clk net1191 VGND VGND VPWR VPWR rvcpu.dp.plmw.PCPlus4W\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_32588_ clknet_leaf_80_clk _04010_ VGND VGND VPWR VPWR datamem.data_ram\[21\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_23390_ _09310_ net1921 _10143_ VGND VGND VPWR VPWR _10146_ sky130_fd_sc_hd__mux2_1
X_23004__709 clknet_1_1__leaf__10085_ VGND VGND VPWR VPWR net835 sky130_fd_sc_hd__inv_2
XFILLER_0_18_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_171_4592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22341_ _09461_ _09502_ _09504_ _09474_ VGND VGND VPWR VPWR _09505_ sky130_fd_sc_hd__o211a_1
X_31539_ clknet_leaf_75_clk net1263 VGND VGND VPWR VPWR rvcpu.dp.plem.funct3M\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25060_ _10758_ net3739 _10752_ VGND VGND VPWR VPWR _10759_ sky130_fd_sc_hd__mux2_1
X_22272_ _09437_ VGND VGND VPWR VPWR _09438_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_60_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_227_5938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21223_ _08468_ _07461_ _08489_ VGND VGND VPWR VPWR _04434_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_238_clk clknet_5_20__leaf_clk VGND VGND VPWR VPWR clknet_leaf_238_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_103_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_227_5949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_184_4920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold120 rvcpu.dp.plfd.InstrD\[3\] VGND VGND VPWR VPWR net1270 sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 rvcpu.dp.plem.ALUResultM\[14\] VGND VGND VPWR VPWR net1281 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_4038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold142 datamem.data_ram\[0\]\[2\] VGND VGND VPWR VPWR net1292 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_4049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold153 rvcpu.dp.plem.ALUResultM\[31\] VGND VGND VPWR VPWR net1303 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold164 datamem.data_ram\[41\]\[5\] VGND VGND VPWR VPWR net1314 sky130_fd_sc_hd__dlygate4sd3_1
X_21154_ datamem.data_ram\[30\]\[23\] datamem.data_ram\[31\]\[23\] _07824_ VGND VGND
+ VPWR VPWR _08443_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_74_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold175 datamem.data_ram\[46\]\[1\] VGND VGND VPWR VPWR net1325 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_180_4806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold186 datamem.data_ram\[46\]\[5\] VGND VGND VPWR VPWR net1336 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_180_4817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_306 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold197 datamem.data_ram\[40\]\[3\] VGND VGND VPWR VPWR net1347 sky130_fd_sc_hd__dlygate4sd3_1
X_20105_ datamem.data_ram\[10\]\[10\] _06754_ _06810_ _07398_ VGND VGND VPWR VPWR
+ _07399_ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28750_ _12747_ net2501 net41 VGND VGND VPWR VPWR _12875_ sky130_fd_sc_hd__mux2_1
X_21085_ datamem.data_ram\[33\]\[7\] _06946_ _08373_ _06615_ VGND VGND VPWR VPWR _08374_
+ sky130_fd_sc_hd__a22o_1
X_25962_ net27 _11289_ VGND VGND VPWR VPWR _11304_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_6_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27701_ _12288_ VGND VGND VPWR VPWR _03702_ sky130_fd_sc_hd__clkbuf_1
X_20036_ datamem.data_ram\[22\]\[26\] _07085_ _06705_ datamem.data_ram\[23\]\[26\]
+ VGND VGND VPWR VPWR _07330_ sky130_fd_sc_hd__o22a_1
X_24913_ _10674_ VGND VGND VPWR VPWR _02528_ sky130_fd_sc_hd__clkbuf_1
X_28681_ _12838_ VGND VGND VPWR VPWR _04132_ sky130_fd_sc_hd__clkbuf_1
X_25893_ _13387_ _11256_ _11258_ _11264_ VGND VGND VPWR VPWR _02918_ sky130_fd_sc_hd__o211a_1
XFILLER_0_137_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_225_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27632_ _10520_ _10908_ _12168_ VGND VGND VPWR VPWR _12251_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_77_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24844_ _10450_ net3214 _10631_ VGND VGND VPWR VPWR _10637_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_178_4757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27563_ _12214_ VGND VGND VPWR VPWR _03638_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_178_4768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24775_ _10597_ VGND VGND VPWR VPWR _02467_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_213_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_178_4779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21987_ _05391_ net117 _09216_ VGND VGND VPWR VPWR _09217_ sky130_fd_sc_hd__a21o_1
X_29302_ clknet_leaf_1_clk _01037_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD1E\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_197_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20938_ datamem.data_ram\[48\]\[22\] _07828_ _07839_ VGND VGND VPWR VPWR _08228_
+ sky130_fd_sc_hd__o21a_1
X_27494_ _12177_ VGND VGND VPWR VPWR _03606_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29233_ _13136_ VGND VGND VPWR VPWR _04386_ sky130_fd_sc_hd__clkbuf_1
X_26445_ _06492_ _11539_ _11529_ _11205_ _11574_ VGND VGND VPWR VPWR _11575_ sky130_fd_sc_hd__a221o_1
XFILLER_0_193_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23206__857 clknet_1_1__leaf__10112_ VGND VGND VPWR VPWR net983 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_42_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20869_ _07833_ _08155_ _08158_ VGND VGND VPWR VPWR _08159_ sky130_fd_sc_hd__a21o_1
XFILLER_0_187_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29164_ _09247_ net2779 net64 VGND VGND VPWR VPWR _13099_ sky130_fd_sc_hd__mux2_1
X_22608_ _09705_ _09750_ _09754_ _09758_ VGND VGND VPWR VPWR _09759_ sky130_fd_sc_hd__and4_1
X_26376_ rvcpu.dp.plde.JalrE VGND VGND VPWR VPWR _11524_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_187_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_3775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_3786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28115_ _12363_ net4127 net74 VGND VGND VPWR VPWR _12523_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25327_ _10598_ _10908_ _10828_ VGND VGND VPWR VPWR _10909_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_180_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29095_ _13062_ VGND VGND VPWR VPWR _04322_ sky130_fd_sc_hd__clkbuf_1
X_22539_ rvcpu.dp.rf.reg_file_arr\[28\]\[12\] rvcpu.dp.rf.reg_file_arr\[30\]\[12\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[12\] rvcpu.dp.rf.reg_file_arr\[31\]\[12\] _09400_
+ _09484_ VGND VGND VPWR VPWR _09693_ sky130_fd_sc_hd__mux4_1
XFILLER_0_221_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_228_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28046_ _12486_ VGND VGND VPWR VPWR _03849_ sky130_fd_sc_hd__clkbuf_1
X_16060_ _14370_ VGND VGND VPWR VPWR _01992_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_224_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25258_ _10538_ net1506 _10867_ _10870_ VGND VGND VPWR VPWR _02677_ sky130_fd_sc_hd__a31o_1
XFILLER_0_224_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15011_ _13558_ VGND VGND VPWR VPWR _13559_ sky130_fd_sc_hd__buf_2
XFILLER_0_20_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_229_clk clknet_5_20__leaf_clk VGND VGND VPWR VPWR clknet_leaf_229_clk
+ sky130_fd_sc_hd__clkbuf_8
X_24209_ _09318_ net4052 _10270_ VGND VGND VPWR VPWR _10275_ sky130_fd_sc_hd__mux2_1
X_25189_ _10832_ VGND VGND VPWR VPWR _02646_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29997_ net367 _01732_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[14\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_19750_ datamem.data_ram\[42\]\[25\] _06754_ _06810_ _07044_ VGND VGND VPWR VPWR
+ _07045_ sky130_fd_sc_hd__o211a_1
X_28948_ _12739_ net4033 net67 VGND VGND VPWR VPWR _12981_ sky130_fd_sc_hd__mux2_1
X_16962_ net3396 _14445_ _04731_ VGND VGND VPWR VPWR _04733_ sky130_fd_sc_hd__mux2_1
X_23252__899 clknet_1_1__leaf__10127_ VGND VGND VPWR VPWR net1025 sky130_fd_sc_hd__inv_2
X_18701_ _05410_ _06053_ VGND VGND VPWR VPWR _06054_ sky130_fd_sc_hd__xnor2_1
X_15913_ net2345 _13229_ _14286_ VGND VGND VPWR VPWR _14292_ sky130_fd_sc_hd__mux2_1
X_19681_ _06976_ VGND VGND VPWR VPWR _06977_ sky130_fd_sc_hd__buf_4
X_16893_ _04696_ VGND VGND VPWR VPWR _01593_ sky130_fd_sc_hd__clkbuf_1
X_28879_ _12756_ net3145 _12941_ VGND VGND VPWR VPWR _12944_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18632_ _05901_ _05892_ _05799_ VGND VGND VPWR VPWR _05989_ sky130_fd_sc_hd__mux2_1
X_30910_ clknet_leaf_281_clk _02645_ VGND VGND VPWR VPWR datamem.data_ram\[41\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_15844_ net2402 _13232_ _14247_ VGND VGND VPWR VPWR _14254_ sky130_fd_sc_hd__mux2_1
X_31890_ clknet_leaf_113_clk _03344_ VGND VGND VPWR VPWR datamem.data_ram\[36\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30841_ clknet_leaf_261_clk _02576_ VGND VGND VPWR VPWR datamem.data_ram\[44\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_18563_ _05782_ _05922_ VGND VGND VPWR VPWR _05923_ sky130_fd_sc_hd__or2_1
X_15775_ _14164_ net2847 _14210_ VGND VGND VPWR VPWR _14217_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23598__218 clknet_1_0__leaf__10178_ VGND VGND VPWR VPWR net344 sky130_fd_sc_hd__inv_2
XFILLER_0_8_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14726_ _13279_ VGND VGND VPWR VPWR _03172_ sky130_fd_sc_hd__clkbuf_1
X_17514_ _13226_ net2782 _05021_ VGND VGND VPWR VPWR _05026_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18494_ _05313_ _05334_ _05500_ _05506_ _05684_ _05668_ VGND VGND VPWR VPWR _05856_
+ sky130_fd_sc_hd__mux4_1
X_30772_ clknet_leaf_172_clk _02507_ VGND VGND VPWR VPWR datamem.data_ram\[47\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_482 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_560 _09401_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_571 _06610_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_185_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32511_ clknet_leaf_184_clk _03933_ VGND VGND VPWR VPWR datamem.data_ram\[24\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_17445_ _04989_ VGND VGND VPWR VPWR _01318_ sky130_fd_sc_hd__clkbuf_1
X_14657_ _13227_ VGND VGND VPWR VPWR _03189_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_184_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_200_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_185_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32442_ clknet_leaf_87_clk _03864_ VGND VGND VPWR VPWR datamem.data_ram\[27\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17376_ _14158_ net3514 _04949_ VGND VGND VPWR VPWR _04953_ sky130_fd_sc_hd__mux2_1
X_14588_ _13172_ VGND VGND VPWR VPWR _13173_ sky130_fd_sc_hd__buf_4
XFILLER_0_171_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19115_ rvcpu.dp.plde.ImmExtE\[13\] rvcpu.dp.plde.PCE\[13\] VGND VGND VPWR VPWR _06435_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_171_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16327_ _14527_ VGND VGND VPWR VPWR _01874_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_171_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32373_ clknet_leaf_263_clk _03795_ VGND VGND VPWR VPWR datamem.data_ram\[2\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19046_ _06373_ _06374_ VGND VGND VPWR VPWR _06375_ sky130_fd_sc_hd__nor2_1
X_31324_ clknet_leaf_18_clk _03027_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCPlus4E\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16258_ net4082 _14424_ _14489_ VGND VGND VPWR VPWR _14491_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15209_ _13493_ VGND VGND VPWR VPWR _13751_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31255_ clknet_leaf_20_clk _02958_ VGND VGND VPWR VPWR rvcpu.dp.plfd.InstrD\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16189_ _14444_ VGND VGND VPWR VPWR _01937_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__10103_ clknet_0__10103_ VGND VGND VPWR VPWR clknet_1_0__leaf__10103_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_3_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30206_ net560 _01941_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[8\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31186_ clknet_leaf_40_clk _02889_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCPlus4D\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_222_5813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_206_Left_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_227_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_222_5824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_222_5835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30137_ net499 _01872_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[10\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_19948_ _06653_ VGND VGND VPWR VPWR _07242_ sky130_fd_sc_hd__buf_4
XFILLER_0_208_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23311__952 clknet_1_0__leaf__10133_ VGND VGND VPWR VPWR net1078 sky130_fd_sc_hd__inv_2
XFILLER_0_177_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30068_ net430 _01803_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[12\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_19879_ datamem.data_ram\[23\]\[1\] _06927_ _07173_ _07081_ VGND VGND VPWR VPWR _07174_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_156_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21910_ rvcpu.dp.rf.reg_file_arr\[16\]\[28\] rvcpu.dp.rf.reg_file_arr\[17\]\[28\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[28\] rvcpu.dp.rf.reg_file_arr\[19\]\[28\] _08516_
+ _08518_ VGND VGND VPWR VPWR _09144_ sky130_fd_sc_hd__mux4_1
XFILLER_0_156_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22890_ rvcpu.dp.rf.reg_file_arr\[20\]\[31\] rvcpu.dp.rf.reg_file_arr\[21\]\[31\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[31\] rvcpu.dp.rf.reg_file_arr\[23\]\[31\] _09384_
+ _09577_ VGND VGND VPWR VPWR _10025_ sky130_fd_sc_hd__mux4_1
XFILLER_0_218_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21841_ _08532_ _09078_ VGND VGND VPWR VPWR _09079_ sky130_fd_sc_hd__nor2_1
XFILLER_0_179_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_194_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24560_ _10479_ VGND VGND VPWR VPWR _02370_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_215_Left_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21772_ rvcpu.dp.rf.reg_file_arr\[4\]\[20\] rvcpu.dp.rf.reg_file_arr\[5\]\[20\] rvcpu.dp.rf.reg_file_arr\[6\]\[20\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[20\] _08628_ _08856_ VGND VGND VPWR VPWR _09014_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_172_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23511_ _09236_ net4343 _10162_ VGND VGND VPWR VPWR _10164_ sky130_fd_sc_hd__mux2_1
X_20723_ datamem.data_ram\[16\]\[6\] datamem.data_ram\[17\]\[6\] _07837_ VGND VGND
+ VPWR VPWR _08013_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_173_4643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32709_ clknet_leaf_79_clk _04131_ VGND VGND VPWR VPWR datamem.data_ram\[17\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_173_4654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24491_ _09322_ datamem.data_ram\[52\]\[29\] _10430_ VGND VGND VPWR VPWR _10436_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26230_ _09478_ _11371_ _11369_ VGND VGND VPWR VPWR _11455_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20654_ datamem.data_ram\[32\]\[29\] _06647_ _07944_ _06679_ VGND VGND VPWR VPWR
+ _07945_ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26161_ _11417_ VGND VGND VPWR VPWR _03033_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_191_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20585_ _07867_ _07875_ VGND VGND VPWR VPWR _07876_ sky130_fd_sc_hd__or2_1
XFILLER_0_162_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25112_ _10787_ VGND VGND VPWR VPWR _02614_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_76_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22324_ _09488_ VGND VGND VPWR VPWR _09489_ sky130_fd_sc_hd__buf_2
X_26092_ net1660 _11372_ VGND VGND VPWR VPWR _11381_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_132_3661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_132_3672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29920_ net290 _01655_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[16\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_25043_ _10476_ net2791 net90 VGND VGND VPWR VPWR _10748_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_72_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22255_ rvcpu.dp.plfd.InstrD\[22\] VGND VGND VPWR VPWR _09421_ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_224_Left_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21206_ _06580_ _08354_ VGND VGND VPWR VPWR _08486_ sky130_fd_sc_hd__nor2_1
X_22186_ _09365_ VGND VGND VPWR VPWR _01110_ sky130_fd_sc_hd__clkbuf_1
X_29851_ net229 _01586_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[18\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28802_ _12747_ net4183 _12896_ VGND VGND VPWR VPWR _12903_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_109_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21137_ datamem.data_ram\[50\]\[23\] datamem.data_ram\[51\]\[23\] _07825_ VGND VGND
+ VPWR VPWR _08426_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_109_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26994_ _11881_ VGND VGND VPWR VPWR _03402_ sky130_fd_sc_hd__clkbuf_1
X_29782_ net1128 _01517_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[20\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_217_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21068_ datamem.data_ram\[60\]\[7\] _06944_ _08356_ _06666_ _06640_ VGND VGND VPWR
+ VPWR _08357_ sky130_fd_sc_hd__a221o_1
X_25945_ rvcpu.dp.pcreg.q\[26\] _11290_ _11286_ _11294_ VGND VGND VPWR VPWR _02940_
+ sky130_fd_sc_hd__o211a_1
X_28733_ _12764_ net2344 _12859_ VGND VGND VPWR VPWR _12866_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_31_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20019_ datamem.data_ram\[34\]\[2\] _06930_ _06600_ _07312_ VGND VGND VPWR VPWR _07313_
+ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_31_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28664_ _12829_ VGND VGND VPWR VPWR _04124_ sky130_fd_sc_hd__clkbuf_1
X_25876_ _11252_ _11247_ VGND VGND VPWR VPWR _11253_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_198_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23089__769 clknet_1_1__leaf__10102_ VGND VGND VPWR VPWR net895 sky130_fd_sc_hd__inv_2
XFILLER_0_9_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24827_ _10627_ VGND VGND VPWR VPWR _02489_ sky130_fd_sc_hd__clkbuf_1
X_27615_ _10520_ _10898_ _12168_ VGND VGND VPWR VPWR _12242_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_216_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_214_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28595_ _12792_ VGND VGND VPWR VPWR _04092_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_198_566 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15560_ _13419_ _13370_ _13301_ _13336_ VGND VGND VPWR VPWR _14084_ sky130_fd_sc_hd__o22a_1
X_27546_ _12205_ VGND VGND VPWR VPWR _03630_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24758_ _10588_ VGND VGND VPWR VPWR _02459_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_3826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_3837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15491_ _14005_ _14007_ _14013_ _14019_ VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__o31a_1
XFILLER_0_189_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27477_ _10500_ VGND VGND VPWR VPWR _12168_ sky130_fd_sc_hd__buf_6
XFILLER_0_166_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24689_ _10551_ VGND VGND VPWR VPWR _02427_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_29_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17230_ _14149_ net3506 _04865_ VGND VGND VPWR VPWR _04875_ sky130_fd_sc_hd__mux2_1
X_26428_ _06453_ _11539_ _11529_ _11190_ _11562_ VGND VGND VPWR VPWR _11563_ sky130_fd_sc_hd__a221o_1
X_29216_ _11533_ net1416 _13122_ _13127_ VGND VGND VPWR VPWR _04378_ sky130_fd_sc_hd__a31o_1
XFILLER_0_138_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17161_ _04838_ VGND VGND VPWR VPWR _01459_ sky130_fd_sc_hd__clkbuf_1
X_29147_ _09281_ net3266 net39 VGND VGND VPWR VPWR _13090_ sky130_fd_sc_hd__mux2_1
X_26359_ _11501_ net1408 _11510_ _11513_ VGND VGND VPWR VPWR _03135_ sky130_fd_sc_hd__a31o_1
XFILLER_0_37_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16112_ _14398_ VGND VGND VPWR VPWR _01968_ sky130_fd_sc_hd__clkbuf_1
X_29078_ _13053_ VGND VGND VPWR VPWR _04314_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17092_ _14147_ net4154 _04793_ VGND VGND VPWR VPWR _04802_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28029_ _12437_ net3372 _12473_ VGND VGND VPWR VPWR _12477_ sky130_fd_sc_hd__mux2_1
X_16043_ net2197 _13217_ _14360_ VGND VGND VPWR VPWR _14362_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_108_Right_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_177_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31040_ clknet_leaf_59_clk _02775_ VGND VGND VPWR VPWR datamem.data_ram\[41\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_1290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_208_103 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19802_ datamem.data_ram\[15\]\[9\] _06761_ _06783_ datamem.data_ram\[9\]\[9\] VGND
+ VGND VPWR VPWR _07097_ sky130_fd_sc_hd__o22a_1
X_17994_ rvcpu.dp.plem.ALUResultM\[4\] _05339_ _05340_ _13265_ VGND VGND VPWR VPWR
+ _05364_ sky130_fd_sc_hd__o22a_1
XFILLER_0_202_1187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19733_ _06683_ VGND VGND VPWR VPWR _07028_ sky130_fd_sc_hd__buf_8
XFILLER_0_198_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16945_ net1880 _14428_ _04720_ VGND VGND VPWR VPWR _04724_ sky130_fd_sc_hd__mux2_1
X_32991_ clknet_leaf_194_clk _04413_ VGND VGND VPWR VPWR datamem.data_ram\[62\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_23606__225 clknet_1_1__leaf__10179_ VGND VGND VPWR VPWR net351 sky130_fd_sc_hd__inv_2
X_31942_ clknet_leaf_113_clk _03364_ VGND VGND VPWR VPWR datamem.data_ram\[59\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_19664_ datamem.data_ram\[46\]\[0\] _06952_ _06958_ datamem.data_ram\[41\]\[0\] _06959_
+ VGND VGND VPWR VPWR _06960_ sky130_fd_sc_hd__a221o_1
XFILLER_0_159_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16876_ _04687_ VGND VGND VPWR VPWR _01601_ sky130_fd_sc_hd__clkbuf_1
X_18615_ _05879_ _05972_ _05957_ _05786_ VGND VGND VPWR VPWR _05973_ sky130_fd_sc_hd__o2bb2a_1
X_15827_ net4120 _13207_ _14236_ VGND VGND VPWR VPWR _14245_ sky130_fd_sc_hd__mux2_1
X_31873_ clknet_leaf_122_clk _03327_ VGND VGND VPWR VPWR datamem.data_ram\[56\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19595_ datamem.data_ram\[59\]\[8\] _06634_ _06887_ _06890_ VGND VGND VPWR VPWR _06891_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_204_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18546_ _05903_ _05906_ _05370_ VGND VGND VPWR VPWR _05907_ sky130_fd_sc_hd__mux2_1
X_30824_ clknet_leaf_224_clk _02559_ VGND VGND VPWR VPWR datamem.data_ram\[44\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_15758_ _14147_ net2908 _14199_ VGND VGND VPWR VPWR _14208_ sky130_fd_sc_hd__mux2_1
X_14709_ net2006 _13266_ _13245_ VGND VGND VPWR VPWR _13267_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_215_5650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18477_ _05456_ _05463_ _05684_ VGND VGND VPWR VPWR _05839_ sky130_fd_sc_hd__mux2_1
X_30755_ clknet_leaf_177_clk _02490_ VGND VGND VPWR VPWR datamem.data_ram\[48\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_15689_ _14163_ VGND VGND VPWR VPWR _02172_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_390 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_215_5661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17428_ _04980_ VGND VGND VPWR VPWR _01326_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30686_ clknet_leaf_174_clk _02421_ VGND VGND VPWR VPWR datamem.data_ram\[4\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_211_5558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32425_ clknet_leaf_248_clk _03847_ VGND VGND VPWR VPWR datamem.data_ram\[28\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_211_5569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_606 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17359_ _14141_ net2270 _04938_ VGND VGND VPWR VPWR _04944_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload310 clknet_1_0__leaf__10172_ VGND VGND VPWR VPWR clkload310/X sky130_fd_sc_hd__clkbuf_8
X_20370_ datamem.data_ram\[32\]\[28\] _06807_ _07658_ _07661_ VGND VGND VPWR VPWR
+ _07662_ sky130_fd_sc_hd__o211a_1
Xclkload321 clknet_1_1__leaf__10156_ VGND VGND VPWR VPWR clkload321/Y sky130_fd_sc_hd__clkinvlp_4
X_32356_ clknet_leaf_256_clk _03778_ VGND VGND VPWR VPWR datamem.data_ram\[30\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload332 clknet_1_1__leaf__10138_ VGND VGND VPWR VPWR clkload332/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload40 clknet_leaf_26_clk VGND VGND VPWR VPWR clkload40/Y sky130_fd_sc_hd__clkinv_1
XFILLER_0_141_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload343 clknet_1_0__leaf__10125_ VGND VGND VPWR VPWR clkload343/Y sky130_fd_sc_hd__clkinvlp_4
X_31307_ clknet_leaf_49_clk _03010_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCPlus4E\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_19029_ rvcpu.dp.plde.ImmExtE\[2\] rvcpu.dp.plde.PCE\[2\] VGND VGND VPWR VPWR _06360_
+ sky130_fd_sc_hd__nand2_1
Xclkload51 clknet_leaf_11_clk VGND VGND VPWR VPWR clkload51/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_3_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload354 clknet_1_0__leaf__10080_ VGND VGND VPWR VPWR clkload354/Y sky130_fd_sc_hd__inv_6
Xclkload62 clknet_leaf_77_clk VGND VGND VPWR VPWR clkload62/Y sky130_fd_sc_hd__clkinv_1
X_32287_ clknet_leaf_276_clk _03709_ VGND VGND VPWR VPWR datamem.data_ram\[33\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload73 clknet_leaf_55_clk VGND VGND VPWR VPWR clkload73/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_140_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload84 clknet_leaf_47_clk VGND VGND VPWR VPWR clkload84/Y sky130_fd_sc_hd__inv_8
X_22040_ rvcpu.dp.plem.ALUResultM\[1\] _09213_ VGND VGND VPWR VPWR _09262_ sky130_fd_sc_hd__nor2_2
X_31238_ clknet_leaf_34_clk _02941_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCD\[27\] sky130_fd_sc_hd__dfxtp_1
Xclkload95 clknet_leaf_82_clk VGND VGND VPWR VPWR clkload95/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_140_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_166_4480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_166_4491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31169_ clknet_leaf_13_clk rvcpu.ALUResultE\[28\] VGND VGND VPWR VPWR rvcpu.dp.plem.ALUResultM\[28\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2802 datamem.data_ram\[34\]\[27\] VGND VGND VPWR VPWR net3952 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2813 datamem.data_ram\[56\]\[27\] VGND VGND VPWR VPWR net3963 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2824 datamem.data_ram\[61\]\[26\] VGND VGND VPWR VPWR net3974 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2835 datamem.data_ram\[35\]\[5\] VGND VGND VPWR VPWR net3985 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_162_4377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2846 datamem.data_ram\[58\]\[10\] VGND VGND VPWR VPWR net3996 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2857 datamem.data_ram\[22\]\[21\] VGND VGND VPWR VPWR net4007 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_162_4388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2868 datamem.data_ram\[48\]\[28\] VGND VGND VPWR VPWR net4018 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2879 datamem.data_ram\[57\]\[30\] VGND VGND VPWR VPWR net4029 sky130_fd_sc_hd__dlygate4sd3_1
X_25730_ _10822_ net3292 _11133_ VGND VGND VPWR VPWR _11139_ sky130_fd_sc_hd__mux2_1
X_22942_ _10070_ _10053_ VGND VGND VPWR VPWR _10071_ sky130_fd_sc_hd__and2_1
XFILLER_0_138_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23995__529 clknet_1_1__leaf__10240_ VGND VGND VPWR VPWR net655 sky130_fd_sc_hd__inv_2
XFILLER_0_183_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25661_ _11078_ _11098_ VGND VGND VPWR VPWR _11099_ sky130_fd_sc_hd__and2_1
XFILLER_0_223_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22873_ rvcpu.dp.rf.reg_file_arr\[28\]\[30\] rvcpu.dp.rf.reg_file_arr\[30\]\[30\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[30\] rvcpu.dp.rf.reg_file_arr\[31\]\[30\] _09381_
+ _09423_ VGND VGND VPWR VPWR _10009_ sky130_fd_sc_hd__mux4_1
XFILLER_0_190_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_175_4705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27400_ _12087_ net3119 net85 VGND VGND VPWR VPWR _12120_ sky130_fd_sc_hd__mux2_1
XFILLER_0_211_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24612_ _10508_ VGND VGND VPWR VPWR _02393_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_65_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28380_ _12665_ VGND VGND VPWR VPWR _04004_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_65_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21824_ _08523_ _09062_ _08748_ VGND VGND VPWR VPWR _09063_ sky130_fd_sc_hd__o21ai_1
X_25592_ _11057_ net1563 _11053_ _11059_ VGND VGND VPWR VPWR _02822_ sky130_fd_sc_hd__a31o_1
XFILLER_0_149_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_65_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_3395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27331_ _10073_ _12076_ _12077_ net1790 VGND VGND VPWR VPWR _03541_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24543_ _09305_ VGND VGND VPWR VPWR _10468_ sky130_fd_sc_hd__clkbuf_2
X_21755_ _08692_ _08995_ _08997_ VGND VGND VPWR VPWR _08998_ sky130_fd_sc_hd__a21o_1
X_20706_ datamem.data_ram\[11\]\[5\] _07137_ _07993_ _07996_ VGND VGND VPWR VPWR _07997_
+ sky130_fd_sc_hd__a211o_1
X_27262_ _10073_ _12041_ _12042_ net1319 VGND VGND VPWR VPWR _03509_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24474_ _09322_ net3284 _10421_ VGND VGND VPWR VPWR _10427_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_3701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21686_ _08817_ _08930_ _08932_ _08700_ VGND VGND VPWR VPWR _08933_ sky130_fd_sc_hd__a211o_1
XFILLER_0_93_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24032__563 clknet_1_0__leaf__10243_ VGND VGND VPWR VPWR net689 sky130_fd_sc_hd__inv_2
XFILLER_0_110_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29001_ _12995_ net1402 _13009_ _13011_ VGND VGND VPWR VPWR _04279_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_134_3712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26213_ rvcpu.dp.plfd.InstrD\[6\] rvcpu.dp.plfd.InstrD\[3\] _11376_ rvcpu.dp.plfd.InstrD\[4\]
+ VGND VGND VPWR VPWR _11444_ sky130_fd_sc_hd__or4b_2
XTAP_TAPCELL_ROW_134_3723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload1 clknet_5_1__leaf_clk VGND VGND VPWR VPWR clkload1/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_135_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27193_ _11991_ net1570 _11995_ _12004_ VGND VGND VPWR VPWR _03478_ sky130_fd_sc_hd__a31o_1
XFILLER_0_117_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20637_ datamem.data_ram\[11\]\[29\] _06737_ _06619_ datamem.data_ram\[12\]\[29\]
+ _07927_ VGND VGND VPWR VPWR _07928_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_24_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26144_ _11371_ VGND VGND VPWR VPWR _11408_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_130_3609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20568_ _06922_ VGND VGND VPWR VPWR _07859_ sky130_fd_sc_hd__buf_4
XFILLER_0_6_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22995__701 clknet_1_1__leaf__10084_ VGND VGND VPWR VPWR net827 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_95_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22307_ rvcpu.dp.plfd.InstrD\[23\] VGND VGND VPWR VPWR _09472_ sky130_fd_sc_hd__clkbuf_4
X_26075_ _11368_ VGND VGND VPWR VPWR _02995_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23318__958 clknet_1_1__leaf__10134_ VGND VGND VPWR VPWR net1084 sky130_fd_sc_hd__inv_2
X_20499_ _07131_ _07787_ _07789_ VGND VGND VPWR VPWR _07790_ sky130_fd_sc_hd__and3_1
XFILLER_0_221_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29903_ clknet_leaf_145_clk _01638_ VGND VGND VPWR VPWR datamem.data_ram\[59\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_25026_ _10737_ net2107 _10725_ VGND VGND VPWR VPWR _10738_ sky130_fd_sc_hd__mux2_1
X_22238_ rvcpu.dp.plfd.InstrD\[23\] VGND VGND VPWR VPWR _09404_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_218_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29834_ net212 _01569_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[1\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22169_ _09314_ net2290 _09352_ VGND VGND VPWR VPWR _09356_ sky130_fd_sc_hd__mux2_1
XFILLER_0_218_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_54_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14991_ _13538_ VGND VGND VPWR VPWR _13539_ sky130_fd_sc_hd__clkbuf_4
X_29765_ net1111 _01500_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[20\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_54_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26977_ _11863_ net1787 _11865_ _11872_ VGND VGND VPWR VPWR _03394_ sky130_fd_sc_hd__a31o_1
XFILLER_0_227_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16730_ _04609_ VGND VGND VPWR VPWR _01677_ sky130_fd_sc_hd__clkbuf_1
X_28716_ _12700_ net2854 _12850_ VGND VGND VPWR VPWR _12857_ sky130_fd_sc_hd__mux2_1
X_25928_ net1295 _11279_ VGND VGND VPWR VPWR _11284_ sky130_fd_sc_hd__or2_1
X_29696_ net1042 _01431_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[23\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_50_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16661_ _14193_ net2900 _04539_ VGND VGND VPWR VPWR _04573_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25859_ rvcpu.dp.pcreg.q\[28\] _11234_ VGND VGND VPWR VPWR _11239_ sky130_fd_sc_hd__and2_1
X_28647_ _12820_ VGND VGND VPWR VPWR _04116_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18400_ _05705_ _05759_ _05763_ VGND VGND VPWR VPWR _05764_ sky130_fd_sc_hd__o21a_1
X_15612_ _14091_ VGND VGND VPWR VPWR _14114_ sky130_fd_sc_hd__buf_4
X_19380_ _06675_ VGND VGND VPWR VPWR _06676_ sky130_fd_sc_hd__buf_8
X_16592_ _14193_ net2970 _04502_ VGND VGND VPWR VPWR _04536_ sky130_fd_sc_hd__mux2_1
X_28578_ _12783_ VGND VGND VPWR VPWR _04084_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15543_ _14064_ _14065_ _14068_ _13466_ VGND VGND VPWR VPWR _14069_ sky130_fd_sc_hd__a31o_1
XFILLER_0_186_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18331_ _05375_ VGND VGND VPWR VPWR _05696_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_201_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27529_ _12196_ VGND VGND VPWR VPWR _03622_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18262_ _05626_ _05464_ VGND VGND VPWR VPWR _05627_ sky130_fd_sc_hd__or2_1
X_30540_ clknet_leaf_199_clk _02275_ VGND VGND VPWR VPWR datamem.data_ram\[55\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_15474_ _13893_ VGND VGND VPWR VPWR _14003_ sky130_fd_sc_hd__inv_2
XFILLER_0_167_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17213_ _04866_ VGND VGND VPWR VPWR _01435_ sky130_fd_sc_hd__clkbuf_1
X_18193_ _05305_ _05555_ _05557_ VGND VGND VPWR VPWR _05558_ sky130_fd_sc_hd__o21a_1
X_30471_ net149 _02206_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[19\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17144_ _14127_ net3524 _04829_ VGND VGND VPWR VPWR _04830_ sky130_fd_sc_hd__mux2_1
X_32210_ clknet_leaf_273_clk _03632_ VGND VGND VPWR VPWR datamem.data_ram\[36\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_208_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold708 rvcpu.dp.plfd.PCPlus4D\[22\] VGND VGND VPWR VPWR net1858 sky130_fd_sc_hd__dlygate4sd3_1
X_32141_ clknet_leaf_263_clk _03563_ VGND VGND VPWR VPWR datamem.data_ram\[39\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold719 rvcpu.dp.pcreg.q\[17\] VGND VGND VPWR VPWR net1869 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17075_ _04792_ VGND VGND VPWR VPWR _04793_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_204_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16026_ net2335 _13190_ _14349_ VGND VGND VPWR VPWR _14353_ sky130_fd_sc_hd__mux2_1
X_32072_ clknet_leaf_121_clk _03494_ VGND VGND VPWR VPWR datamem.data_ram\[29\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_228_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31023_ clknet_leaf_60_clk _02758_ VGND VGND VPWR VPWR datamem.data_ram\[40\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_139_Left_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_198_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2109 datamem.data_ram\[29\]\[14\] VGND VGND VPWR VPWR net3259 sky130_fd_sc_hd__dlygate4sd3_1
X_17977_ _05347_ _05339_ VGND VGND VPWR VPWR _05348_ sky130_fd_sc_hd__nor2_1
Xhold1408 rvcpu.dp.rf.reg_file_arr\[0\]\[0\] VGND VGND VPWR VPWR net2558 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_204_5384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1419 rvcpu.dp.rf.reg_file_arr\[7\]\[25\] VGND VGND VPWR VPWR net2569 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_204_5395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19716_ datamem.data_ram\[26\]\[0\] _06989_ _07010_ _07011_ VGND VGND VPWR VPWR _07012_
+ sky130_fd_sc_hd__a211o_1
X_16928_ _04714_ VGND VGND VPWR VPWR _01576_ sky130_fd_sc_hd__clkbuf_1
X_32974_ clknet_leaf_138_clk _04396_ VGND VGND VPWR VPWR datamem.data_ram\[63\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19647_ _06942_ VGND VGND VPWR VPWR _06943_ sky130_fd_sc_hd__buf_4
X_31925_ _04438_ net118 VGND VGND VPWR VPWR datamem.rd_data_mem\[30\] sky130_fd_sc_hd__dlxtn_1
XFILLER_0_79_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_205_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16859_ net3833 _14478_ _04670_ VGND VGND VPWR VPWR _04678_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_217_5701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_196_5196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_217_5712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31856_ clknet_leaf_111_clk _03310_ VGND VGND VPWR VPWR datamem.data_ram\[62\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19578_ datamem.data_ram\[14\]\[8\] _06683_ _06870_ _06873_ VGND VGND VPWR VPWR _06874_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_177_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_148_Left_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_213_5609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30807_ clknet_leaf_150_clk _02542_ VGND VGND VPWR VPWR datamem.data_ram\[45\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_18529_ _05334_ _05320_ _05327_ _05446_ _05682_ _05579_ VGND VGND VPWR VPWR _05890_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_48_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31787_ clknet_leaf_53_clk _03241_ VGND VGND VPWR VPWR datamem.data_ram\[8\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21540_ _08565_ _08791_ _08793_ _08652_ VGND VGND VPWR VPWR _08794_ sky130_fd_sc_hd__o211a_1
XFILLER_0_117_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30738_ clknet_leaf_221_clk _02473_ VGND VGND VPWR VPWR datamem.data_ram\[47\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21471_ rvcpu.dp.rf.reg_file_arr\[24\]\[5\] rvcpu.dp.rf.reg_file_arr\[25\]\[5\] rvcpu.dp.rf.reg_file_arr\[26\]\[5\]
+ rvcpu.dp.rf.reg_file_arr\[27\]\[5\] _08517_ _08519_ VGND VGND VPWR VPWR _08728_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_15_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23576__198 clknet_1_1__leaf__10176_ VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__inv_2
XFILLER_0_62_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30669_ clknet_leaf_179_clk _02404_ VGND VGND VPWR VPWR datamem.data_ram\[50\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20422_ _06715_ _07702_ _07713_ _06712_ VGND VGND VPWR VPWR _07714_ sky130_fd_sc_hd__o211a_1
X_32408_ clknet_leaf_276_clk _03830_ VGND VGND VPWR VPWR datamem.data_ram\[29\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_168_4520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_168_4531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload140 clknet_leaf_245_clk VGND VGND VPWR VPWR clkload140/Y sky130_fd_sc_hd__clkinv_4
X_20353_ _06916_ _07631_ _07644_ _06985_ VGND VGND VPWR VPWR _07645_ sky130_fd_sc_hd__a211o_1
X_32339_ clknet_leaf_240_clk _03761_ VGND VGND VPWR VPWR datamem.data_ram\[30\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload151 clknet_leaf_273_clk VGND VGND VPWR VPWR clkload151/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_144_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload162 clknet_leaf_181_clk VGND VGND VPWR VPWR clkload162/Y sky130_fd_sc_hd__bufinv_16
Xclkload173 clknet_leaf_228_clk VGND VGND VPWR VPWR clkload173/Y sky130_fd_sc_hd__clkinvlp_4
XPHY_EDGE_ROW_157_Left_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload184 clknet_leaf_217_clk VGND VGND VPWR VPWR clkload184/Y sky130_fd_sc_hd__clkinvlp_2
X_20284_ datamem.data_ram\[24\]\[19\] _06697_ _07024_ datamem.data_ram\[28\]\[19\]
+ _07576_ VGND VGND VPWR VPWR _07577_ sky130_fd_sc_hd__o221a_1
X_23072_ _09282_ net4414 _10093_ VGND VGND VPWR VPWR _10098_ sky130_fd_sc_hd__mux2_1
Xclkload195 clknet_leaf_185_clk VGND VGND VPWR VPWR clkload195/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_101_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_164_4428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3300 rvcpu.dp.pcreg.q\[11\] VGND VGND VPWR VPWR net4450 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_164_4439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26900_ _11813_ net1441 _11821_ _11824_ VGND VGND VPWR VPWR _03365_ sky130_fd_sc_hd__a31o_1
X_22023_ _09248_ net4311 _09232_ VGND VGND VPWR VPWR _09249_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_90_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27880_ _12155_ net2002 _12382_ VGND VGND VPWR VPWR _12389_ sky130_fd_sc_hd__mux2_1
X_24062__589 clknet_1_0__leaf__10247_ VGND VGND VPWR VPWR net715 sky130_fd_sc_hd__inv_2
Xhold2610 datamem.data_ram\[56\]\[21\] VGND VGND VPWR VPWR net3760 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2621 datamem.data_ram\[37\]\[10\] VGND VGND VPWR VPWR net3771 sky130_fd_sc_hd__dlygate4sd3_1
X_26831_ _11689_ _11774_ VGND VGND VPWR VPWR _11782_ sky130_fd_sc_hd__and2_1
Xhold13 rvcpu.dp.plem.PCPlus4M\[1\] VGND VGND VPWR VPWR net1163 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 rvcpu.dp.plde.PCPlus4E\[3\] VGND VGND VPWR VPWR net1174 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2632 datamem.data_ram\[61\]\[11\] VGND VGND VPWR VPWR net3782 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 rvcpu.dp.plem.PCPlus4M\[2\] VGND VGND VPWR VPWR net1185 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2643 datamem.data_ram\[62\]\[30\] VGND VGND VPWR VPWR net3793 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 rvcpu.dp.plde.PCPlus4E\[26\] VGND VGND VPWR VPWR net1196 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2654 datamem.data_ram\[44\]\[18\] VGND VGND VPWR VPWR net3804 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1920 datamem.data_ram\[43\]\[16\] VGND VGND VPWR VPWR net3070 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2665 rvcpu.dp.rf.reg_file_arr\[9\]\[8\] VGND VGND VPWR VPWR net3815 sky130_fd_sc_hd__dlygate4sd3_1
X_26762_ _11681_ _11738_ VGND VGND VPWR VPWR _11741_ sky130_fd_sc_hd__and2_1
Xhold57 rvcpu.dp.plem.ResultSrcM\[1\] VGND VGND VPWR VPWR net1207 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1931 datamem.data_ram\[23\]\[16\] VGND VGND VPWR VPWR net3081 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2676 datamem.data_ram\[27\]\[8\] VGND VGND VPWR VPWR net3826 sky130_fd_sc_hd__dlygate4sd3_1
X_29550_ net904 _01285_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[27\]\[17\] sky130_fd_sc_hd__dfxtp_1
Xhold68 rvcpu.dp.plde.PCPlus4E\[30\] VGND VGND VPWR VPWR net1218 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1942 datamem.data_ram\[55\]\[29\] VGND VGND VPWR VPWR net3092 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_67_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold79 rvcpu.dp.plem.PCPlus4M\[17\] VGND VGND VPWR VPWR net1229 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2687 datamem.data_ram\[58\]\[14\] VGND VGND VPWR VPWR net3837 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1953 datamem.data_ram\[34\]\[24\] VGND VGND VPWR VPWR net3103 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2698 rvcpu.dp.rf.reg_file_arr\[31\]\[2\] VGND VGND VPWR VPWR net3848 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_3446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1964 datamem.data_ram\[41\]\[15\] VGND VGND VPWR VPWR net3114 sky130_fd_sc_hd__dlygate4sd3_1
X_28501_ _12734_ net4108 net43 VGND VGND VPWR VPWR _12736_ sky130_fd_sc_hd__mux2_1
X_25713_ _10822_ net2576 _11124_ VGND VGND VPWR VPWR _11130_ sky130_fd_sc_hd__mux2_1
X_22925_ _10057_ VGND VGND VPWR VPWR _10058_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_123_3457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1975 rvcpu.dp.rf.reg_file_arr\[14\]\[22\] VGND VGND VPWR VPWR net3125 sky130_fd_sc_hd__dlygate4sd3_1
X_26693_ _11687_ _11694_ VGND VGND VPWR VPWR _11701_ sky130_fd_sc_hd__and2_1
XFILLER_0_196_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1986 datamem.data_ram\[45\]\[18\] VGND VGND VPWR VPWR net3136 sky130_fd_sc_hd__dlygate4sd3_1
X_29481_ net843 _01216_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[2\]\[20\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__10262_ clknet_0__10262_ VGND VGND VPWR VPWR clknet_1_1__leaf__10262_
+ sky130_fd_sc_hd__clkbuf_16
Xhold1997 rvcpu.dp.rf.reg_file_arr\[17\]\[15\] VGND VGND VPWR VPWR net3147 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25644_ _11091_ _11079_ VGND VGND VPWR VPWR _11092_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_166_Left_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28432_ _12695_ VGND VGND VPWR VPWR _04026_ sky130_fd_sc_hd__clkbuf_1
X_22856_ _09390_ _09992_ VGND VGND VPWR VPWR _09993_ sky130_fd_sc_hd__or2_1
Xclkbuf_1_1__f__10193_ clknet_0__10193_ VGND VGND VPWR VPWR clknet_1_1__leaf__10193_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21807_ _08626_ _09040_ _09042_ _09046_ _08509_ VGND VGND VPWR VPWR _09047_ sky130_fd_sc_hd__a311o_1
X_28363_ _12656_ VGND VGND VPWR VPWR _03996_ sky130_fd_sc_hd__clkbuf_1
X_25575_ _11018_ net1423 _11041_ _11048_ VGND VGND VPWR VPWR _02816_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_26_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22787_ rvcpu.dp.rf.reg_file_arr\[12\]\[25\] rvcpu.dp.rf.reg_file_arr\[13\]\[25\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[25\] rvcpu.dp.rf.reg_file_arr\[15\]\[25\] _09386_
+ _09419_ VGND VGND VPWR VPWR _09928_ sky130_fd_sc_hd__mux4_1
XFILLER_0_38_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27314_ _11976_ _12066_ VGND VGND VPWR VPWR _12072_ sky130_fd_sc_hd__and2_1
XFILLER_0_136_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24526_ _10458_ VGND VGND VPWR VPWR _02357_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_213_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28294_ _12619_ VGND VGND VPWR VPWR _03964_ sky130_fd_sc_hd__clkbuf_1
X_21738_ rvcpu.dp.rf.reg_file_arr\[4\]\[18\] rvcpu.dp.rf.reg_file_arr\[5\]\[18\] rvcpu.dp.rf.reg_file_arr\[6\]\[18\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[18\] _08839_ _08840_ VGND VGND VPWR VPWR _08982_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_66_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27245_ _11918_ VGND VGND VPWR VPWR _12036_ sky130_fd_sc_hd__buf_2
XFILLER_0_152_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24457_ _10412_ net1835 _10404_ _10417_ VGND VGND VPWR VPWR _02329_ sky130_fd_sc_hd__a31o_1
XFILLER_0_191_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21669_ _08916_ VGND VGND VPWR VPWR _01042_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_193_Right_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15190_ _13344_ _13548_ _13533_ VGND VGND VPWR VPWR _13733_ sky130_fd_sc_hd__a21oi_1
X_27176_ _11994_ VGND VGND VPWR VPWR _11995_ sky130_fd_sc_hd__buf_2
XFILLER_0_163_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24388_ _09252_ net4206 _10367_ VGND VGND VPWR VPWR _10373_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26127_ _11399_ VGND VGND VPWR VPWR _03016_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26058_ _11089_ _11351_ VGND VGND VPWR VPWR _11358_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_1079 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17900_ rvcpu.dp.plem.ALUResultM\[31\] _05272_ VGND VGND VPWR VPWR _05273_ sky130_fd_sc_hd__and2_1
X_25009_ _10726_ VGND VGND VPWR VPWR _02572_ sky130_fd_sc_hd__clkbuf_1
X_18880_ _06215_ _06219_ _06221_ _06222_ VGND VGND VPWR VPWR _06223_ sky130_fd_sc_hd__a211o_1
XFILLER_0_197_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_207_916 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17831_ _13209_ rvcpu.dp.plde.RD2E\[22\] _05196_ VGND VGND VPWR VPWR _05215_ sky130_fd_sc_hd__mux2_1
X_29817_ net195 _01552_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[1\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_17762_ _14346_ rvcpu.dp.plde.Rs2E\[0\] rvcpu.dp.plmw.RegWriteW VGND VGND VPWR VPWR
+ _05160_ sky130_fd_sc_hd__o21a_1
X_29748_ net1094 _01483_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[21\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_14974_ _13469_ _13486_ _13500_ _13522_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__o211ai_2
XFILLER_0_89_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19501_ _06796_ VGND VGND VPWR VPWR _06797_ sky130_fd_sc_hd__buf_8
X_16713_ _14177_ net3219 _04598_ VGND VGND VPWR VPWR _04601_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17693_ _13187_ net2201 _05118_ VGND VGND VPWR VPWR _05121_ sky130_fd_sc_hd__mux2_1
X_29679_ net1025 _01414_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[23\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31710_ clknet_leaf_31_clk _03168_ VGND VGND VPWR VPWR rvcpu.dp.pcreg.q\[28\] sky130_fd_sc_hd__dfxtp_1
X_19432_ _06690_ VGND VGND VPWR VPWR _06728_ sky130_fd_sc_hd__buf_6
XFILLER_0_202_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16644_ _04564_ VGND VGND VPWR VPWR _01718_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_190_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32690_ clknet_leaf_273_clk _04112_ VGND VGND VPWR VPWR datamem.data_ram\[18\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31641_ clknet_leaf_69_clk net1166 VGND VGND VPWR VPWR rvcpu.dp.plmw.lAuiPCW\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_19363_ _06658_ VGND VGND VPWR VPWR _06659_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_191_5071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16575_ _04527_ VGND VGND VPWR VPWR _01758_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_174_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_191_5082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18314_ _05365_ VGND VGND VPWR VPWR _05679_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15526_ _13572_ _14036_ _14041_ _14052_ VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__o31a_1
X_31572_ clknet_leaf_71_clk datamem.rd_data_mem\[22\] VGND VGND VPWR VPWR rvcpu.dp.plmw.ReadDataW\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_19294_ _06583_ _06589_ VGND VGND VPWR VPWR _06590_ sky130_fd_sc_hd__or2_1
X_23495__141 clknet_1_1__leaf__10160_ VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__inv_2
XFILLER_0_44_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15457_ _13985_ _13986_ _13501_ VGND VGND VPWR VPWR _13987_ sky130_fd_sc_hd__a21oi_1
X_30523_ clknet_leaf_140_clk _02258_ VGND VGND VPWR VPWR datamem.data_ram\[56\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_18245_ _05327_ VGND VGND VPWR VPWR _05610_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30454_ net132 _02189_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[19\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_15388_ _13297_ _13422_ _13586_ VGND VGND VPWR VPWR _13921_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_160_Right_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18176_ _05539_ _05540_ VGND VGND VPWR VPWR _05541_ sky130_fd_sc_hd__nor2_1
XFILLER_0_163_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17127_ _04820_ VGND VGND VPWR VPWR _01475_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold505 datamem.data_ram\[11\]\[6\] VGND VGND VPWR VPWR net1655 sky130_fd_sc_hd__dlygate4sd3_1
X_30385_ clknet_leaf_269_clk _02120_ VGND VGND VPWR VPWR datamem.data_ram\[58\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold516 datamem.data_ram\[32\]\[5\] VGND VGND VPWR VPWR net1666 sky130_fd_sc_hd__dlygate4sd3_1
Xhold527 datamem.data_ram\[2\]\[4\] VGND VGND VPWR VPWR net1677 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold538 datamem.data_ram\[9\]\[1\] VGND VGND VPWR VPWR net1688 sky130_fd_sc_hd__dlygate4sd3_1
X_17058_ net2878 _14472_ _04779_ VGND VGND VPWR VPWR _04784_ sky130_fd_sc_hd__mux2_1
X_32124_ clknet_leaf_228_clk _03546_ VGND VGND VPWR VPWR datamem.data_ram\[7\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold549 datamem.data_ram\[9\]\[4\] VGND VGND VPWR VPWR net1699 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_206_5435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16009_ _14342_ VGND VGND VPWR VPWR _02023_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_206_5446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32055_ clknet_leaf_131_clk _03477_ VGND VGND VPWR VPWR datamem.data_ram\[30\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_31006_ clknet_leaf_158_clk _02741_ VGND VGND VPWR VPWR datamem.data_ram\[11\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_198_5236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1205 rvcpu.dp.rf.reg_file_arr\[1\]\[8\] VGND VGND VPWR VPWR net2355 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_198_5247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1216 rvcpu.dp.rf.reg_file_arr\[18\]\[16\] VGND VGND VPWR VPWR net2366 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_198_5258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1227 datamem.data_ram\[43\]\[30\] VGND VGND VPWR VPWR net2377 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1238 rvcpu.dp.rf.reg_file_arr\[26\]\[13\] VGND VGND VPWR VPWR net2388 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1249 rvcpu.dp.rf.reg_file_arr\[9\]\[26\] VGND VGND VPWR VPWR net2399 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32957_ clknet_leaf_99_clk _04379_ VGND VGND VPWR VPWR datamem.data_ram\[6\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20971_ datamem.data_ram\[32\]\[15\] _06935_ _08257_ _06641_ _08259_ VGND VGND VPWR
+ VPWR _08260_ sky130_fd_sc_hd__a221o_1
XFILLER_0_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22710_ rvcpu.dp.rf.reg_file_arr\[24\]\[21\] rvcpu.dp.rf.reg_file_arr\[25\]\[21\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[21\] rvcpu.dp.rf.reg_file_arr\[27\]\[21\] _09484_
+ _09431_ VGND VGND VPWR VPWR _09855_ sky130_fd_sc_hd__mux4_1
X_31908_ _04419_ net118 VGND VGND VPWR VPWR datamem.rd_data_mem\[13\] sky130_fd_sc_hd__dlxtn_1
XFILLER_0_75_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32888_ clknet_leaf_281_clk _04310_ VGND VGND VPWR VPWR datamem.data_ram\[10\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_178_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_157_4254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22641_ _09528_ _09788_ _09789_ VGND VGND VPWR VPWR _09790_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_157_4265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31839_ clknet_leaf_162_clk _03293_ VGND VGND VPWR VPWR datamem.data_ram\[8\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25360_ _10416_ _10923_ VGND VGND VPWR VPWR _10929_ sky130_fd_sc_hd__and2_1
X_22572_ _09705_ _09713_ _09719_ _09724_ VGND VGND VPWR VPWR _09725_ sky130_fd_sc_hd__and4_1
XFILLER_0_8_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_180_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24311_ _09310_ net3374 _10328_ VGND VGND VPWR VPWR _10331_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21523_ rvcpu.dp.rf.reg_file_arr\[16\]\[8\] rvcpu.dp.rf.reg_file_arr\[17\]\[8\] rvcpu.dp.rf.reg_file_arr\[18\]\[8\]
+ rvcpu.dp.rf.reg_file_arr\[19\]\[8\] _08703_ _08721_ VGND VGND VPWR VPWR _08777_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_7_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25291_ _10888_ VGND VGND VPWR VPWR _02692_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27030_ _11889_ net1425 _11897_ _11903_ VGND VGND VPWR VPWR _03416_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_21_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24242_ _10292_ VGND VGND VPWR VPWR _02239_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_161_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21454_ _08511_ _08711_ VGND VGND VPWR VPWR _08712_ sky130_fd_sc_hd__nor2_1
XFILLER_0_133_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_116_3272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20405_ datamem.data_ram\[40\]\[12\] _06820_ _06617_ datamem.data_ram\[44\]\[12\]
+ VGND VGND VPWR VPWR _07697_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_92_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24173_ clknet_1_1__leaf__10079_ VGND VGND VPWR VPWR _10265_ sky130_fd_sc_hd__buf_1
XFILLER_0_32_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21385_ _08542_ _08645_ VGND VGND VPWR VPWR _08646_ sky130_fd_sc_hd__or2_1
XFILLER_0_142_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_187_4973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_187_4984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20336_ datamem.data_ram\[38\]\[4\] _06951_ _06954_ datamem.data_ram\[36\]\[4\] _07627_
+ VGND VGND VPWR VPWR _07628_ sky130_fd_sc_hd__a221o_1
Xoutput14 net14 VGND VGND VPWR VPWR Instr[20] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_187_4995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput25 net25 VGND VGND VPWR VPWR Instr[30] sky130_fd_sc_hd__buf_2
X_28981_ _12687_ net4024 _12999_ VGND VGND VPWR VPWR _13000_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_129_3600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__11601_ _11601_ VGND VGND VPWR VPWR clknet_0__11601_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_12_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27932_ _12136_ net3339 _12412_ VGND VGND VPWR VPWR _12418_ sky130_fd_sc_hd__mux2_1
X_23055_ clknet_1_1__leaf__10087_ VGND VGND VPWR VPWR _10091_ sky130_fd_sc_hd__buf_1
X_20267_ datamem.data_ram\[62\]\[19\] _06719_ _06738_ datamem.data_ram\[59\]\[19\]
+ _07559_ VGND VGND VPWR VPWR _07560_ sky130_fd_sc_hd__o221a_1
Xhold3130 datamem.data_ram\[10\]\[11\] VGND VGND VPWR VPWR net4280 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_179_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22006_ rvcpu.dp.plem.WriteDataM\[1\] _09215_ _09219_ _09234_ VGND VGND VPWR VPWR
+ _09235_ sky130_fd_sc_hd__a31o_4
Xhold3141 datamem.data_ram\[54\]\[18\] VGND VGND VPWR VPWR net4291 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3152 datamem.data_ram\[5\]\[20\] VGND VGND VPWR VPWR net4302 sky130_fd_sc_hd__dlygate4sd3_1
X_27863_ _12138_ net1997 _12373_ VGND VGND VPWR VPWR _12380_ sky130_fd_sc_hd__mux2_1
Xhold3163 rvcpu.dp.rf.reg_file_arr\[13\]\[7\] VGND VGND VPWR VPWR net4313 sky130_fd_sc_hd__dlygate4sd3_1
X_20198_ datamem.data_ram\[37\]\[11\] _06703_ _07489_ _07490_ VGND VGND VPWR VPWR
+ _07491_ sky130_fd_sc_hd__o211a_1
Xhold3174 rvcpu.dp.rf.reg_file_arr\[23\]\[12\] VGND VGND VPWR VPWR net4324 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2440 rvcpu.dp.rf.reg_file_arr\[4\]\[13\] VGND VGND VPWR VPWR net3590 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3185 rvcpu.dp.rf.reg_file_arr\[24\]\[16\] VGND VGND VPWR VPWR net4335 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2451 datamem.data_ram\[27\]\[17\] VGND VGND VPWR VPWR net3601 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29602_ net956 _01337_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[25\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_26814_ _11767_ net1561 _11761_ _11771_ VGND VGND VPWR VPWR _03332_ sky130_fd_sc_hd__a31o_1
XFILLER_0_192_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold3196 rvcpu.dp.rf.reg_file_arr\[26\]\[25\] VGND VGND VPWR VPWR net4346 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_192_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_146_3991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2462 datamem.data_ram\[17\]\[25\] VGND VGND VPWR VPWR net3612 sky130_fd_sc_hd__dlygate4sd3_1
X_27794_ _12130_ net2620 _12336_ VGND VGND VPWR VPWR _12339_ sky130_fd_sc_hd__mux2_1
Xhold2473 datamem.data_ram\[9\]\[8\] VGND VGND VPWR VPWR net3623 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2484 datamem.data_ram\[20\]\[20\] VGND VGND VPWR VPWR net3634 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_174_Left_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2495 datamem.data_ram\[31\]\[28\] VGND VGND VPWR VPWR net3645 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1750 rvcpu.dp.rf.reg_file_arr\[14\]\[1\] VGND VGND VPWR VPWR net2900 sky130_fd_sc_hd__dlygate4sd3_1
X_29533_ net887 _01268_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[27\]\[0\] sky130_fd_sc_hd__dfxtp_1
Xhold1761 rvcpu.dp.rf.reg_file_arr\[15\]\[17\] VGND VGND VPWR VPWR net2911 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_86_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26745_ _11700_ net1752 _11724_ _11730_ VGND VGND VPWR VPWR _03304_ sky130_fd_sc_hd__a31o_1
X_23957_ _10232_ VGND VGND VPWR VPWR _02014_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_4_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1772 datamem.data_ram\[22\]\[27\] VGND VGND VPWR VPWR net2922 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1783 rvcpu.dp.rf.reg_file_arr\[29\]\[11\] VGND VGND VPWR VPWR net2933 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_142_3899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1794 datamem.data_ram\[1\]\[26\] VGND VGND VPWR VPWR net2944 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22908_ _08144_ VGND VGND VPWR VPWR _10042_ sky130_fd_sc_hd__buf_4
XFILLER_0_86_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26676_ _11683_ net1832 _11675_ _11690_ VGND VGND VPWR VPWR _03275_ sky130_fd_sc_hd__a31o_1
X_14690_ _13252_ VGND VGND VPWR VPWR _03181_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29464_ net826 _01199_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[2\]\[3\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__10245_ clknet_0__10245_ VGND VGND VPWR VPWR clknet_1_1__leaf__10245_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_212_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_631 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28415_ _12684_ VGND VGND VPWR VPWR _04020_ sky130_fd_sc_hd__clkbuf_1
X_25627_ _11057_ net1564 _11077_ _11080_ VGND VGND VPWR VPWR _02836_ sky130_fd_sc_hd__a31o_1
X_22839_ _09442_ _09972_ _09974_ _09976_ VGND VGND VPWR VPWR _09977_ sky130_fd_sc_hd__o2bb2a_1
X_29395_ clknet_leaf_2_clk _01130_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD2E\[6\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__10176_ clknet_0__10176_ VGND VGND VPWR VPWR clknet_1_1__leaf__10176_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_49_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24112__619 clknet_1_1__leaf__10259_ VGND VGND VPWR VPWR net745 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_15_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16360_ _14544_ VGND VGND VPWR VPWR _01858_ sky130_fd_sc_hd__clkbuf_1
X_25558_ _11037_ VGND VGND VPWR VPWR _02810_ sky130_fd_sc_hd__clkbuf_1
X_28346_ _12647_ VGND VGND VPWR VPWR _03988_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15311_ _13767_ _13324_ _13847_ _13823_ _13319_ VGND VGND VPWR VPWR _13848_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_13_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24509_ _10447_ VGND VGND VPWR VPWR _02351_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16291_ net4235 _14457_ _14500_ VGND VGND VPWR VPWR _14508_ sky130_fd_sc_hd__mux2_1
X_28277_ _12369_ net2573 _12603_ VGND VGND VPWR VPWR _12610_ sky130_fd_sc_hd__mux2_1
X_25489_ _10570_ _10997_ _10998_ VGND VGND VPWR VPWR _10999_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_124_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15242_ _13428_ _13703_ _13574_ _13312_ VGND VGND VPWR VPWR _13782_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_183_Left_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18030_ _05383_ _05397_ _05399_ VGND VGND VPWR VPWR _05400_ sky130_fd_sc_hd__a21o_1
X_27228_ _11976_ _12019_ VGND VGND VPWR VPWR _12026_ sky130_fd_sc_hd__and2_1
XFILLER_0_164_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15173_ _13326_ _13714_ _13715_ _13504_ VGND VGND VPWR VPWR _13716_ sky130_fd_sc_hd__a22o_1
X_27159_ _11974_ net1491 _11983_ _11985_ VGND VGND VPWR VPWR _03463_ sky130_fd_sc_hd__a31o_1
XFILLER_0_34_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_607 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30170_ net532 _01905_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[0\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_19981_ _06716_ _07263_ _07274_ _06985_ VGND VGND VPWR VPWR _07275_ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18932_ _05714_ _06270_ _05670_ VGND VGND VPWR VPWR _06271_ sky130_fd_sc_hd__mux2_1
XFILLER_0_185_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_1174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18863_ _05481_ _05573_ _05618_ VGND VGND VPWR VPWR _06207_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_201_5310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_201_5321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_192_Left_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22973__681 clknet_1_0__leaf__10082_ VGND VGND VPWR VPWR net807 sky130_fd_sc_hd__inv_2
X_17814_ rvcpu.dp.plem.ALUResultM\[28\] _05203_ _05178_ VGND VGND VPWR VPWR _05204_
+ sky130_fd_sc_hd__mux2_1
X_18794_ _05706_ _06141_ VGND VGND VPWR VPWR _06142_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32811_ clknet_leaf_255_clk _04233_ VGND VGND VPWR VPWR datamem.data_ram\[13\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_17745_ _13266_ net3690 _05140_ VGND VGND VPWR VPWR _05148_ sky130_fd_sc_hd__mux2_1
XFILLER_0_222_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14957_ _13287_ _13281_ VGND VGND VPWR VPWR _13506_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_193_5122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_193_5133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32742_ clknet_leaf_284_clk _04164_ VGND VGND VPWR VPWR datamem.data_ram\[16\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17676_ _05111_ VGND VGND VPWR VPWR _01201_ sky130_fd_sc_hd__clkbuf_1
X_14888_ _13413_ _13418_ _13421_ _13437_ _13439_ VGND VGND VPWR VPWR _13440_ sky130_fd_sc_hd__a32o_1
XFILLER_0_43_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_212_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19415_ _06604_ _06638_ _06674_ _06710_ VGND VGND VPWR VPWR _06711_ sky130_fd_sc_hd__a31o_1
X_16627_ _04555_ VGND VGND VPWR VPWR _01726_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26486__40 clknet_1_1__leaf__10267_ VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__inv_2
X_32673_ clknet_leaf_244_clk _04095_ VGND VGND VPWR VPWR datamem.data_ram\[18\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31624_ clknet_leaf_64_clk net1169 VGND VGND VPWR VPWR rvcpu.dp.plmw.lAuiPCW\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19346_ _06640_ _06641_ VGND VGND VPWR VPWR _06642_ sky130_fd_sc_hd__nor2_4
XFILLER_0_9_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16558_ _04518_ VGND VGND VPWR VPWR _01766_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_898 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_210_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15509_ _13458_ _14035_ VGND VGND VPWR VPWR _14036_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_152_4140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1072 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31555_ clknet_leaf_63_clk datamem.rd_data_mem\[5\] VGND VGND VPWR VPWR rvcpu.dp.plmw.ReadDataW\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_19277_ _06575_ rvcpu.c.ad.funct7b5 _06574_ VGND VGND VPWR VPWR _06576_ sky130_fd_sc_hd__or3b_1
XFILLER_0_155_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_152_4151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16489_ net3474 _14449_ _04478_ VGND VGND VPWR VPWR _04482_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18228_ _05588_ _05591_ _05592_ VGND VGND VPWR VPWR _05593_ sky130_fd_sc_hd__o21ba_1
X_30506_ clknet_leaf_268_clk _02241_ VGND VGND VPWR VPWR datamem.data_ram\[57\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31486_ clknet_leaf_52_clk rvcpu.dp.lAuiPCE\[12\] VGND VGND VPWR VPWR rvcpu.dp.plem.lAuiPCM\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_23731__323 clknet_1_1__leaf__10198_ VGND VGND VPWR VPWR net449 sky130_fd_sc_hd__inv_2
XFILLER_0_143_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18159_ _05482_ _05519_ _05523_ VGND VGND VPWR VPWR _05524_ sky130_fd_sc_hd__a21o_1
X_30437_ net775 _02172_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[29\]\[16\] sky130_fd_sc_hd__dfxtp_1
Xhold302 datamem.data_ram\[43\]\[4\] VGND VGND VPWR VPWR net1452 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__10265_ clknet_0__10265_ VGND VGND VPWR VPWR clknet_1_0__leaf__10265_
+ sky130_fd_sc_hd__clkbuf_16
Xhold313 datamem.data_ram\[11\]\[2\] VGND VGND VPWR VPWR net1463 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23374__1009 clknet_1_1__leaf__10139_ VGND VGND VPWR VPWR net1135 sky130_fd_sc_hd__inv_2
Xhold324 datamem.data_ram\[48\]\[4\] VGND VGND VPWR VPWR net1474 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_229_5980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold335 datamem.data_ram\[20\]\[0\] VGND VGND VPWR VPWR net1485 sky130_fd_sc_hd__dlygate4sd3_1
X_21170_ datamem.data_ram\[14\]\[23\] datamem.data_ram\[15\]\[23\] _07824_ VGND VGND
+ VPWR VPWR _08459_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_229_5991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold346 datamem.data_ram\[49\]\[4\] VGND VGND VPWR VPWR net1496 sky130_fd_sc_hd__dlygate4sd3_1
X_30368_ net714 _02103_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[3\]\[19\] sky130_fd_sc_hd__dfxtp_1
Xhold357 datamem.data_ram\[50\]\[4\] VGND VGND VPWR VPWR net1507 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23846__410 clknet_1_1__leaf__10208_ VGND VGND VPWR VPWR net536 sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__10196_ clknet_0__10196_ VGND VGND VPWR VPWR clknet_1_0__leaf__10196_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_229_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold368 datamem.data_ram\[24\]\[0\] VGND VGND VPWR VPWR net1518 sky130_fd_sc_hd__dlygate4sd3_1
X_32107_ clknet_leaf_120_clk _03529_ VGND VGND VPWR VPWR datamem.data_ram\[58\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_20121_ _06912_ _07276_ _07323_ _07414_ VGND VGND VPWR VPWR _07415_ sky130_fd_sc_hd__o211a_1
Xhold379 datamem.data_ram\[55\]\[0\] VGND VGND VPWR VPWR net1529 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30299_ net645 _02034_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[5\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_225_5888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20052_ datamem.data_ram\[38\]\[26\] _06624_ _06616_ datamem.data_ram\[36\]\[26\]
+ VGND VGND VPWR VPWR _07346_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_225_5899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32038_ clknet_leaf_131_clk _03460_ VGND VGND VPWR VPWR datamem.data_ram\[50\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_182_4870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1002 datamem.data_ram\[6\]\[31\] VGND VGND VPWR VPWR net2152 sky130_fd_sc_hd__dlygate4sd3_1
X_24860_ _10394_ net4181 net93 VGND VGND VPWR VPWR _10646_ sky130_fd_sc_hd__mux2_1
Xhold1013 rvcpu.dp.rf.reg_file_arr\[3\]\[26\] VGND VGND VPWR VPWR net2163 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1024 rvcpu.dp.rf.reg_file_arr\[10\]\[5\] VGND VGND VPWR VPWR net2174 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1035 rvcpu.dp.rf.reg_file_arr\[4\]\[3\] VGND VGND VPWR VPWR net2185 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1046 rvcpu.dp.rf.reg_file_arr\[20\]\[12\] VGND VGND VPWR VPWR net2196 sky130_fd_sc_hd__dlygate4sd3_1
X_23811_ clknet_1_0__leaf__10203_ VGND VGND VPWR VPWR _10207_ sky130_fd_sc_hd__buf_1
XFILLER_0_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1057 rvcpu.dp.rf.reg_file_arr\[2\]\[25\] VGND VGND VPWR VPWR net2207 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_159_4305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1068 rvcpu.dp.rf.reg_file_arr\[21\]\[21\] VGND VGND VPWR VPWR net2218 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_1_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24791_ _10476_ net3886 net94 VGND VGND VPWR VPWR _10608_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_159_4316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1079 rvcpu.dp.rf.reg_file_arr\[6\]\[3\] VGND VGND VPWR VPWR net2229 sky130_fd_sc_hd__dlygate4sd3_1
X_26530_ _07203_ _10946_ _11494_ VGND VGND VPWR VPWR _11607_ sky130_fd_sc_hd__or3_1
XFILLER_0_197_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_208 _09560_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20954_ datamem.data_ram\[49\]\[15\] _06639_ VGND VGND VPWR VPWR _08243_ sky130_fd_sc_hd__or2_1
XANTENNA_219 _09813_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_221_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0__10130_ _10130_ VGND VGND VPWR VPWR clknet_0__10130_ sky130_fd_sc_hd__clkbuf_16
X_26461_ _11576_ _11228_ _11540_ _06525_ _11585_ VGND VGND VPWR VPWR _11586_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_81_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_270 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20885_ _07635_ datamem.data_ram\[62\]\[14\] VGND VGND VPWR VPWR _08175_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23892__452 clknet_1_0__leaf__10222_ VGND VGND VPWR VPWR net578 sky130_fd_sc_hd__inv_2
X_25412_ _10751_ net2528 _10961_ VGND VGND VPWR VPWR _10962_ sky130_fd_sc_hd__mux2_1
X_28200_ _12454_ net3200 net46 VGND VGND VPWR VPWR _12568_ sky130_fd_sc_hd__mux2_1
X_29180_ _13107_ VGND VGND VPWR VPWR _04362_ sky130_fd_sc_hd__clkbuf_1
X_22624_ rvcpu.dp.rf.reg_file_arr\[12\]\[16\] rvcpu.dp.rf.reg_file_arr\[13\]\[16\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[16\] rvcpu.dp.rf.reg_file_arr\[15\]\[16\] _09552_
+ _09721_ VGND VGND VPWR VPWR _09774_ sky130_fd_sc_hd__mux4_1
X_26392_ _06384_ _11522_ _11526_ _11158_ _11536_ VGND VGND VPWR VPWR _11537_ sky130_fd_sc_hd__a221o_1
XFILLER_0_187_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28131_ _12531_ VGND VGND VPWR VPWR _03889_ sky130_fd_sc_hd__clkbuf_1
X_25343_ _10917_ VGND VGND VPWR VPWR _02715_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_118_3334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22555_ _09706_ _09707_ _09421_ VGND VGND VPWR VPWR _09708_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21506_ rvcpu.dp.rf.reg_file_arr\[20\]\[7\] rvcpu.dp.rf.reg_file_arr\[21\]\[7\] rvcpu.dp.rf.reg_file_arr\[22\]\[7\]
+ rvcpu.dp.rf.reg_file_arr\[23\]\[7\] _08631_ _08632_ VGND VGND VPWR VPWR _08761_
+ sky130_fd_sc_hd__mux4_1
X_28062_ _12361_ net3412 _12492_ VGND VGND VPWR VPWR _12495_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_518 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25274_ _10879_ VGND VGND VPWR VPWR _02684_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22486_ _09441_ _09642_ VGND VGND VPWR VPWR _09643_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27013_ _11833_ _11886_ VGND VGND VPWR VPWR _11893_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_40_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24225_ _10283_ VGND VGND VPWR VPWR _02231_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_79_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21437_ _08535_ VGND VGND VPWR VPWR _08696_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_79_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_1130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21368_ _08552_ VGND VGND VPWR VPWR _08629_ sky130_fd_sc_hd__buf_4
XFILLER_0_20_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20319_ datamem.data_ram\[24\]\[4\] _07122_ _07133_ datamem.data_ram\[25\]\[4\] VGND
+ VGND VPWR VPWR _07611_ sky130_fd_sc_hd__a22o_1
X_28964_ _12727_ net1601 _12988_ _12990_ VGND VGND VPWR VPWR _04263_ sky130_fd_sc_hd__a31o_1
X_24087_ _10255_ VGND VGND VPWR VPWR _02121_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21299_ _08536_ VGND VGND VPWR VPWR _08561_ sky130_fd_sc_hd__clkbuf_4
Xhold880 rvcpu.dp.rf.reg_file_arr\[5\]\[15\] VGND VGND VPWR VPWR net2030 sky130_fd_sc_hd__dlygate4sd3_1
Xhold891 rvcpu.dp.rf.reg_file_arr\[28\]\[23\] VGND VGND VPWR VPWR net2041 sky130_fd_sc_hd__dlygate4sd3_1
X_27915_ _12153_ net2132 net47 VGND VGND VPWR VPWR _12409_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28895_ _12952_ VGND VGND VPWR VPWR _04232_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_200_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27846_ _12370_ VGND VGND VPWR VPWR _03765_ sky130_fd_sc_hd__clkbuf_1
X_15860_ _14262_ VGND VGND VPWR VPWR _02092_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_204_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2270 datamem.data_ram\[48\]\[30\] VGND VGND VPWR VPWR net3420 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14811_ _13296_ _13341_ VGND VGND VPWR VPWR _13364_ sky130_fd_sc_hd__nand2_2
XFILLER_0_204_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2281 datamem.data_ram\[41\]\[8\] VGND VGND VPWR VPWR net3431 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2292 rvcpu.dp.rf.reg_file_arr\[12\]\[3\] VGND VGND VPWR VPWR net3442 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_153_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27777_ _12329_ VGND VGND VPWR VPWR _03737_ sky130_fd_sc_hd__clkbuf_1
X_15791_ _14225_ VGND VGND VPWR VPWR _02132_ sky130_fd_sc_hd__clkbuf_1
X_24989_ _10542_ _10630_ _10705_ VGND VGND VPWR VPWR _10715_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_118_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1580 datamem.data_ram\[0\]\[25\] VGND VGND VPWR VPWR net2730 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17530_ _05034_ VGND VGND VPWR VPWR _01278_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29516_ net878 _01251_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[28\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_14742_ rvcpu.dp.pcreg.q\[5\] VGND VGND VPWR VPWR _13295_ sky130_fd_sc_hd__inv_2
X_26728_ _10762_ net4104 _11714_ VGND VGND VPWR VPWR _11720_ sky130_fd_sc_hd__mux2_1
Xhold1591 datamem.data_ram\[33\]\[24\] VGND VGND VPWR VPWR net2741 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_197_973 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17461_ _14175_ net2882 _04996_ VGND VGND VPWR VPWR _04998_ sky130_fd_sc_hd__mux2_1
X_14673_ _13239_ VGND VGND VPWR VPWR _03185_ sky130_fd_sc_hd__clkbuf_1
X_29447_ net809 _01182_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[30\]\[18\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__10228_ clknet_0__10228_ VGND VGND VPWR VPWR clknet_1_1__leaf__10228_
+ sky130_fd_sc_hd__clkbuf_16
X_26659_ _10057_ VGND VGND VPWR VPWR _11679_ sky130_fd_sc_hd__buf_2
XFILLER_0_196_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_192_clk clknet_5_28__leaf_clk VGND VGND VPWR VPWR clknet_leaf_192_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_19_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19200_ _06487_ _06491_ _06496_ _06503_ _06495_ VGND VGND VPWR VPWR _06510_ sky130_fd_sc_hd__a311o_1
XFILLER_0_184_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_103_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16412_ _14560_ VGND VGND VPWR VPWR _14572_ sky130_fd_sc_hd__clkbuf_4
X_23142__817 clknet_1_1__leaf__10107_ VGND VGND VPWR VPWR net943 sky130_fd_sc_hd__inv_2
XFILLER_0_55_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0__10259_ _10259_ VGND VGND VPWR VPWR clknet_0__10259_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_183_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29378_ clknet_leaf_139_clk _01113_ VGND VGND VPWR VPWR datamem.data_ram\[60\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17392_ _04961_ VGND VGND VPWR VPWR _01343_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1__f__10159_ clknet_0__10159_ VGND VGND VPWR VPWR clknet_1_1__leaf__10159_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_55_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_824 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19131_ rvcpu.dp.plde.ImmExtE\[15\] rvcpu.dp.plde.PCE\[15\] VGND VGND VPWR VPWR _06449_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_171_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28329_ _12638_ VGND VGND VPWR VPWR _03980_ sky130_fd_sc_hd__clkbuf_1
X_16343_ _14535_ VGND VGND VPWR VPWR _01866_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19062_ _06382_ VGND VGND VPWR VPWR _06389_ sky130_fd_sc_hd__inv_2
X_31340_ clknet_leaf_13_clk _03043_ VGND VGND VPWR VPWR rvcpu.dp.plde.Rs1E\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16274_ net2985 _14440_ _14489_ VGND VGND VPWR VPWR _14499_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23257__904 clknet_1_0__leaf__10127_ VGND VGND VPWR VPWR net1030 sky130_fd_sc_hd__inv_2
XFILLER_0_109_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_202_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15225_ _13402_ _13484_ _13692_ VGND VGND VPWR VPWR _13766_ sky130_fd_sc_hd__o21a_1
X_18013_ _05380_ _05382_ VGND VGND VPWR VPWR _05383_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_23_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31271_ clknet_leaf_35_clk _02974_ VGND VGND VPWR VPWR rvcpu.dp.plfd.InstrD\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15156_ _13327_ _13699_ VGND VGND VPWR VPWR _13700_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30222_ net576 _01957_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[7\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_196_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30153_ net515 _01888_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[0\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_15087_ _13538_ _13611_ _13629_ _13632_ VGND VGND VPWR VPWR _13633_ sky130_fd_sc_hd__or4_1
X_19964_ datamem.data_ram\[15\]\[18\] _06705_ _06781_ datamem.data_ram\[9\]\[18\]
+ VGND VGND VPWR VPWR _07258_ sky130_fd_sc_hd__o22a_1
XFILLER_0_226_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18915_ _05456_ _05469_ _05533_ _05463_ _05670_ _05769_ VGND VGND VPWR VPWR _06255_
+ sky130_fd_sc_hd__mux4_1
X_30084_ net446 _01819_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[11\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_19895_ _06604_ _07181_ _07184_ _07189_ VGND VGND VPWR VPWR _07190_ sky130_fd_sc_hd__a31o_1
XFILLER_0_129_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18846_ _05563_ _05494_ _06167_ VGND VGND VPWR VPWR _06191_ sky130_fd_sc_hd__and3_1
XFILLER_0_101_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_220_5774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_220_5785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18777_ _05318_ _05728_ _05820_ _06125_ VGND VGND VPWR VPWR _06126_ sky130_fd_sc_hd__a211o_1
XFILLER_0_136_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15989_ net2045 _13241_ _14322_ VGND VGND VPWR VPWR _14332_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17728_ _13241_ net3143 _05129_ VGND VGND VPWR VPWR _05139_ sky130_fd_sc_hd__mux2_1
XFILLER_0_188_940 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30986_ clknet_leaf_117_clk _02721_ VGND VGND VPWR VPWR datamem.data_ram\[39\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32725_ clknet_leaf_244_clk _04147_ VGND VGND VPWR VPWR datamem.data_ram\[16\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_17659_ _05102_ VGND VGND VPWR VPWR _01209_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_154_4202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_183_clk clknet_5_19__leaf_clk VGND VGND VPWR VPWR clknet_leaf_183_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_148_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20670_ datamem.data_ram\[50\]\[29\] _06804_ _07957_ _07960_ VGND VGND VPWR VPWR
+ _07961_ sky130_fd_sc_hd__o211a_1
X_32656_ clknet_leaf_183_clk _04078_ VGND VGND VPWR VPWR datamem.data_ram\[19\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31607_ clknet_leaf_27_clk net1195 VGND VGND VPWR VPWR rvcpu.dp.plmw.PCPlus4W\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_19329_ _06624_ VGND VGND VPWR VPWR _06625_ sky130_fd_sc_hd__buf_6
X_32587_ clknet_leaf_171_clk _04009_ VGND VGND VPWR VPWR datamem.data_ram\[21\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_4593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22340_ _09469_ _09503_ VGND VGND VPWR VPWR _09504_ sky130_fd_sc_hd__or2_1
X_31538_ clknet_leaf_75_clk net1269 VGND VGND VPWR VPWR rvcpu.dp.plem.funct3M\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22271_ _08589_ _09404_ VGND VGND VPWR VPWR _09437_ sky130_fd_sc_hd__nand2_2
X_31469_ clknet_leaf_5_clk rvcpu.dp.SrcBFW_Mux.y\[27\] VGND VGND VPWR VPWR rvcpu.dp.plem.WriteDataM\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_227_5939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_184_4910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21222_ _08468_ _07368_ _08489_ VGND VGND VPWR VPWR _04433_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_143_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold110 rvcpu.dp.plem.RdM\[2\] VGND VGND VPWR VPWR net1260 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_184_4921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold121 rvcpu.dp.plem.RdM\[4\] VGND VGND VPWR VPWR net1271 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold132 rvcpu.dp.plem.ALUResultM\[23\] VGND VGND VPWR VPWR net1282 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_4039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__10248_ clknet_0__10248_ VGND VGND VPWR VPWR clknet_1_0__leaf__10248_
+ sky130_fd_sc_hd__clkbuf_16
Xhold143 rvcpu.dp.plem.ALUResultM\[0\] VGND VGND VPWR VPWR net1293 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold154 datamem.data_ram\[45\]\[4\] VGND VGND VPWR VPWR net1304 sky130_fd_sc_hd__dlygate4sd3_1
X_23445__95 clknet_1_1__leaf__10156_ VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_74_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold165 rvcpu.dp.plfd.InstrD\[26\] VGND VGND VPWR VPWR net1315 sky130_fd_sc_hd__dlygate4sd3_1
X_21153_ datamem.data_ram\[28\]\[23\] datamem.data_ram\[29\]\[23\] _07825_ VGND VGND
+ VPWR VPWR _08442_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_74_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold176 rvcpu.dp.plfd.PCD\[21\] VGND VGND VPWR VPWR net1326 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_180_4807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_4818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24141__645 clknet_1_0__leaf__10262_ VGND VGND VPWR VPWR net771 sky130_fd_sc_hd__inv_2
Xhold187 datamem.data_ram\[40\]\[0\] VGND VGND VPWR VPWR net1337 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__10179_ clknet_0__10179_ VGND VGND VPWR VPWR clknet_1_0__leaf__10179_
+ sky130_fd_sc_hd__clkbuf_16
Xhold198 datamem.data_ram\[46\]\[3\] VGND VGND VPWR VPWR net1348 sky130_fd_sc_hd__dlygate4sd3_1
X_20104_ datamem.data_ram\[12\]\[10\] _06686_ _06656_ datamem.data_ram\[9\]\[10\]
+ _07397_ VGND VGND VPWR VPWR _07398_ sky130_fd_sc_hd__o221a_1
XFILLER_0_217_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21084_ datamem.data_ram\[36\]\[7\] datamem.data_ram\[37\]\[7\] _07912_ VGND VGND
+ VPWR VPWR _08373_ sky130_fd_sc_hd__mux2_1
X_25961_ net4245 _11302_ _11300_ _11303_ VGND VGND VPWR VPWR _02947_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_6_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27700_ _12140_ net1923 _12280_ VGND VGND VPWR VPWR _12288_ sky130_fd_sc_hd__mux2_1
X_20035_ datamem.data_ram\[16\]\[26\] _06778_ _06699_ datamem.data_ram\[17\]\[26\]
+ VGND VGND VPWR VPWR _07329_ sky130_fd_sc_hd__o22a_1
X_24912_ _10394_ net3702 _10669_ VGND VGND VPWR VPWR _10674_ sky130_fd_sc_hd__mux2_1
X_25892_ net1801 _11263_ VGND VGND VPWR VPWR _11264_ sky130_fd_sc_hd__or2_1
X_28680_ _12762_ net2972 _12832_ VGND VGND VPWR VPWR _12838_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27631_ _12250_ VGND VGND VPWR VPWR _03670_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_225_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24843_ _10636_ VGND VGND VPWR VPWR _02496_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_107_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_178_4758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27562_ _12157_ net2209 _12206_ VGND VGND VPWR VPWR _12214_ sky130_fd_sc_hd__mux2_1
X_24774_ _10480_ net2746 _10589_ VGND VGND VPWR VPWR _10597_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_178_4769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21986_ _08488_ VGND VGND VPWR VPWR _09216_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29301_ clknet_leaf_1_clk _01036_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD1E\[8\] sky130_fd_sc_hd__dfxtp_1
X_20937_ datamem.data_ram\[49\]\[22\] _07832_ VGND VGND VPWR VPWR _08227_ sky130_fd_sc_hd__or2_1
X_27493_ _12140_ net2667 _12169_ VGND VGND VPWR VPWR _12177_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_174_clk clknet_5_19__leaf_clk VGND VGND VPWR VPWR clknet_leaf_174_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_178_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23738__329 clknet_1_1__leaf__10199_ VGND VGND VPWR VPWR net455 sky130_fd_sc_hd__inv_2
XFILLER_0_166_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29232_ _09313_ net2460 _13132_ VGND VGND VPWR VPWR _13136_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26444_ _11545_ rvcpu.ALUResultE\[20\] VGND VGND VPWR VPWR _11574_ sky130_fd_sc_hd__and2_1
XFILLER_0_166_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20868_ datamem.data_ram\[35\]\[14\] _07851_ _07836_ _08157_ VGND VGND VPWR VPWR
+ _08158_ sky130_fd_sc_hd__o211a_1
XFILLER_0_194_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22607_ _09627_ _09755_ _09757_ _09438_ VGND VGND VPWR VPWR _09758_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_42_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26375_ _06365_ _11522_ VGND VGND VPWR VPWR _11523_ sky130_fd_sc_hd__and2_1
XFILLER_0_165_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29163_ _13098_ VGND VGND VPWR VPWR _04354_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20799_ datamem.data_ram\[50\]\[30\] _07831_ VGND VGND VPWR VPWR _08089_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_137_3776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_3787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25326_ _09228_ _10897_ VGND VGND VPWR VPWR _10908_ sky130_fd_sc_hd__nor2_8
X_28114_ _12522_ VGND VGND VPWR VPWR _03881_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_221_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22538_ _09391_ _09691_ VGND VGND VPWR VPWR _09692_ sky130_fd_sc_hd__or2_1
XFILLER_0_107_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29094_ _09313_ net2959 net40 VGND VGND VPWR VPWR _13062_ sky130_fd_sc_hd__mux2_1
XFILLER_0_228_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25257_ _10408_ _10868_ VGND VGND VPWR VPWR _10870_ sky130_fd_sc_hd__and2_1
X_28045_ _12452_ net4162 net96 VGND VGND VPWR VPWR _12486_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22469_ _09399_ VGND VGND VPWR VPWR _09627_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_228_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_224_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15010_ _13305_ _13346_ VGND VGND VPWR VPWR _13558_ sky130_fd_sc_hd__or2_1
X_24208_ _10274_ VGND VGND VPWR VPWR _02223_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25188_ _10729_ net2639 net57 VGND VGND VPWR VPWR _10832_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29996_ net366 _01731_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[14\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28947_ _12980_ VGND VGND VPWR VPWR _04256_ sky130_fd_sc_hd__clkbuf_1
X_16961_ _04732_ VGND VGND VPWR VPWR _01561_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_217_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18700_ _05419_ _06036_ _05416_ VGND VGND VPWR VPWR _06053_ sky130_fd_sc_hd__a21oi_1
X_15912_ _14291_ VGND VGND VPWR VPWR _02069_ sky130_fd_sc_hd__clkbuf_1
X_19680_ _06954_ VGND VGND VPWR VPWR _06976_ sky130_fd_sc_hd__buf_4
X_28878_ _12943_ VGND VGND VPWR VPWR _04224_ sky130_fd_sc_hd__clkbuf_1
X_16892_ net3445 _14442_ _04695_ VGND VGND VPWR VPWR _04696_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_217_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18631_ _05692_ _05986_ _05987_ VGND VGND VPWR VPWR _05988_ sky130_fd_sc_hd__o21a_1
X_23899__458 clknet_1_0__leaf__10223_ VGND VGND VPWR VPWR net584 sky130_fd_sc_hd__inv_2
X_27829_ _09305_ VGND VGND VPWR VPWR _12359_ sky130_fd_sc_hd__clkbuf_2
X_15843_ _14253_ VGND VGND VPWR VPWR _02100_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_189_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18562_ _05779_ _05751_ _05674_ VGND VGND VPWR VPWR _05922_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30840_ clknet_leaf_258_clk _02575_ VGND VGND VPWR VPWR datamem.data_ram\[44\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_15774_ _14216_ VGND VGND VPWR VPWR _02140_ sky130_fd_sc_hd__clkbuf_1
X_17513_ _05025_ VGND VGND VPWR VPWR _01286_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23373__1008 clknet_1_0__leaf__10139_ VGND VGND VPWR VPWR net1134 sky130_fd_sc_hd__inv_2
X_14725_ net2232 _13278_ _13180_ VGND VGND VPWR VPWR _13279_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18493_ _05320_ _05327_ _05446_ _05412_ _05769_ _05689_ VGND VGND VPWR VPWR _05855_
+ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_165_clk clknet_5_25__leaf_clk VGND VGND VPWR VPWR clknet_leaf_165_clk
+ sky130_fd_sc_hd__clkbuf_8
X_30771_ clknet_leaf_172_clk _02506_ VGND VGND VPWR VPWR datamem.data_ram\[47\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_197_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_550 _07177_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32510_ clknet_leaf_246_clk _03932_ VGND VGND VPWR VPWR datamem.data_ram\[24\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_561 _09401_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_196_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_572 _06610_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17444_ _14158_ net3866 _04985_ VGND VGND VPWR VPWR _04989_ sky130_fd_sc_hd__mux2_1
X_14656_ net3559 _13226_ _13214_ VGND VGND VPWR VPWR _13227_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32441_ clknet_leaf_77_clk _03863_ VGND VGND VPWR VPWR datamem.data_ram\[27\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17375_ _04952_ VGND VGND VPWR VPWR _01351_ sky130_fd_sc_hd__clkbuf_1
X_14587_ rvcpu.dp.plmw.ALUResultW\[31\] rvcpu.dp.plmw.ReadDataW\[31\] rvcpu.dp.plmw.PCPlus4W\[31\]
+ rvcpu.dp.plmw.lAuiPCW\[31\] _13169_ _13171_ VGND VGND VPWR VPWR _13172_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_188_5010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19114_ rvcpu.dp.plde.ImmExtE\[13\] rvcpu.dp.plde.PCE\[13\] VGND VGND VPWR VPWR _06434_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_172_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16326_ net2517 _14424_ _14525_ VGND VGND VPWR VPWR _14527_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32372_ clknet_leaf_257_clk _03794_ VGND VGND VPWR VPWR datamem.data_ram\[2\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19045_ rvcpu.dp.plde.ImmExtE\[4\] rvcpu.dp.plde.PCE\[4\] VGND VGND VPWR VPWR _06374_
+ sky130_fd_sc_hd__nor2_1
X_31323_ clknet_leaf_18_clk _03026_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCPlus4E\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_16257_ _14490_ VGND VGND VPWR VPWR _01907_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15208_ _13296_ _13393_ VGND VGND VPWR VPWR _13750_ sky130_fd_sc_hd__nand2_1
X_31254_ clknet_leaf_21_clk _02957_ VGND VGND VPWR VPWR rvcpu.dp.plfd.InstrD\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__10102_ clknet_0__10102_ VGND VGND VPWR VPWR clknet_1_0__leaf__10102_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_207_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16188_ net1957 _14442_ _14443_ VGND VGND VPWR VPWR _14444_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30205_ net559 _01940_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[8\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_15139_ _13335_ _13526_ _13681_ _13573_ _13682_ VGND VGND VPWR VPWR _13683_ sky130_fd_sc_hd__a311o_1
XFILLER_0_2_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31185_ clknet_leaf_40_clk _02888_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCPlus4D\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_222_5814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_222_5825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19947_ datamem.data_ram\[54\]\[18\] _07085_ _06646_ datamem.data_ram\[48\]\[18\]
+ VGND VGND VPWR VPWR _07241_ sky130_fd_sc_hd__o22a_1
X_30136_ net498 _01871_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[10\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30067_ net429 _01802_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[12\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_19878_ datamem.data_ram\[22\]\[1\] _06978_ _06973_ datamem.data_ram\[16\]\[1\] _07172_
+ VGND VGND VPWR VPWR _07173_ sky130_fd_sc_hd__a221o_1
XFILLER_0_177_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18829_ _05697_ _06004_ _05872_ _05702_ VGND VGND VPWR VPWR _06175_ sky130_fd_sc_hd__a31o_1
XFILLER_0_65_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21840_ rvcpu.dp.rf.reg_file_arr\[28\]\[24\] rvcpu.dp.rf.reg_file_arr\[30\]\[24\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[24\] rvcpu.dp.rf.reg_file_arr\[31\]\[24\] _08534_
+ _08537_ VGND VGND VPWR VPWR _09078_ sky130_fd_sc_hd__mux4_1
XFILLER_0_222_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21771_ rvcpu.dp.rf.reg_file_arr\[0\]\[20\] rvcpu.dp.rf.reg_file_arr\[1\]\[20\] rvcpu.dp.rf.reg_file_arr\[2\]\[20\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[20\] _08810_ _08811_ VGND VGND VPWR VPWR _09013_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_210_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_188_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_156_clk clknet_5_30__leaf_clk VGND VGND VPWR VPWR clknet_leaf_156_clk
+ sky130_fd_sc_hd__clkbuf_8
X_30969_ clknet_leaf_222_clk _02704_ VGND VGND VPWR VPWR datamem.data_ram\[39\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23510_ _10163_ VGND VGND VPWR VPWR _01636_ sky130_fd_sc_hd__clkbuf_1
X_20722_ _07227_ _07857_ _08012_ VGND VGND VPWR VPWR _04442_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_147_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32708_ clknet_leaf_80_clk _04130_ VGND VGND VPWR VPWR datamem.data_ram\[17\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_173_4644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24490_ _10435_ VGND VGND VPWR VPWR _02344_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_173_4655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20653_ datamem.data_ram\[34\]\[29\] _06610_ _06618_ datamem.data_ram\[36\]\[29\]
+ _07943_ VGND VGND VPWR VPWR _07944_ sky130_fd_sc_hd__o221a_1
XFILLER_0_74_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32639_ clknet_leaf_282_clk _04061_ VGND VGND VPWR VPWR datamem.data_ram\[1\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26160_ net4446 _11408_ VGND VGND VPWR VPWR _11417_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20584_ datamem.data_ram\[48\]\[13\] datamem.data_ram\[49\]\[13\] _07874_ VGND VGND
+ VPWR VPWR _07875_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25111_ _10729_ net2931 net88 VGND VGND VPWR VPWR _10787_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_76_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22323_ rvcpu.dp.plfd.InstrD\[24\] _09411_ VGND VGND VPWR VPWR _09488_ sky130_fd_sc_hd__nor2_2
X_26091_ _11380_ VGND VGND VPWR VPWR _02999_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_171_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23930__485 clknet_1_1__leaf__10227_ VGND VGND VPWR VPWR net611 sky130_fd_sc_hd__inv_2
XFILLER_0_225_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25042_ _10747_ VGND VGND VPWR VPWR _02584_ sky130_fd_sc_hd__clkbuf_1
X_22254_ rvcpu.dp.rf.reg_file_arr\[0\]\[0\] rvcpu.dp.rf.reg_file_arr\[1\]\[0\] rvcpu.dp.rf.reg_file_arr\[2\]\[0\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[0\] _09417_ _09419_ VGND VGND VPWR VPWR _09420_ sky130_fd_sc_hd__mux4_1
XFILLER_0_170_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_72_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21205_ _08485_ VGND VGND VPWR VPWR _04420_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29850_ net228 _01585_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[18\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_22185_ _09240_ net4399 _09362_ VGND VGND VPWR VPWR _09365_ sky130_fd_sc_hd__mux2_1
XFILLER_0_223_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23171__843 clknet_1_0__leaf__10110_ VGND VGND VPWR VPWR net969 sky130_fd_sc_hd__inv_2
X_28801_ _12902_ VGND VGND VPWR VPWR _04188_ sky130_fd_sc_hd__clkbuf_1
X_21136_ datamem.data_ram\[48\]\[23\] _07874_ _07838_ VGND VGND VPWR VPWR _08425_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_109_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29781_ net1127 _01516_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[20\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_109_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26993_ _10762_ net3170 _11875_ VGND VGND VPWR VPWR _11881_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_35_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28732_ _12865_ VGND VGND VPWR VPWR _04156_ sky130_fd_sc_hd__clkbuf_1
X_25944_ net1871 _11155_ VGND VGND VPWR VPWR _11294_ sky130_fd_sc_hd__or2_1
X_21067_ _06585_ datamem.data_ram\[61\]\[7\] VGND VGND VPWR VPWR _08356_ sky130_fd_sc_hd__and2_1
XFILLER_0_214_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20018_ datamem.data_ram\[32\]\[2\] _06935_ _06953_ datamem.data_ram\[36\]\[2\] _07311_
+ VGND VGND VPWR VPWR _07312_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_31_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28663_ _12698_ net3535 _12823_ VGND VGND VPWR VPWR _12829_ sky130_fd_sc_hd__mux2_1
XFILLER_0_226_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25875_ net1795 VGND VGND VPWR VPWR _11252_ sky130_fd_sc_hd__inv_2
XFILLER_0_225_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27614_ _12241_ VGND VGND VPWR VPWR _03662_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_193_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24826_ _10396_ net2013 _10621_ VGND VGND VPWR VPWR _10627_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28594_ _12745_ net3850 _12786_ VGND VGND VPWR VPWR _12792_ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_198_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23972__508 clknet_1_1__leaf__10238_ VGND VGND VPWR VPWR net634 sky130_fd_sc_hd__inv_2
XFILLER_0_201_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27545_ _12140_ net2063 _12197_ VGND VGND VPWR VPWR _12205_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_147_clk clknet_5_29__leaf_clk VGND VGND VPWR VPWR clknet_leaf_147_clk
+ sky130_fd_sc_hd__clkbuf_8
X_24757_ _10400_ net2192 _10580_ VGND VGND VPWR VPWR _10588_ sky130_fd_sc_hd__mux2_1
X_21969_ rvcpu.dp.rf.reg_file_arr\[20\]\[31\] rvcpu.dp.rf.reg_file_arr\[21\]\[31\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[31\] rvcpu.dp.rf.reg_file_arr\[23\]\[31\] _08548_
+ _08552_ VGND VGND VPWR VPWR _09200_ sky130_fd_sc_hd__mux4_1
XFILLER_0_201_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_100_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_3827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15490_ _13439_ _14016_ _14018_ _13776_ _13638_ VGND VGND VPWR VPWR _14019_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_139_3838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24688_ _10400_ net1938 _10543_ VGND VGND VPWR VPWR _10551_ sky130_fd_sc_hd__mux2_1
X_27476_ _12167_ VGND VGND VPWR VPWR _03598_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29215_ _10063_ _13123_ VGND VGND VPWR VPWR _13127_ sky130_fd_sc_hd__and2_1
XFILLER_0_193_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_182_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26427_ _11545_ rvcpu.ALUResultE\[15\] VGND VGND VPWR VPWR _11562_ sky130_fd_sc_hd__and2_1
XFILLER_0_166_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23639_ _09279_ net3490 _10182_ VGND VGND VPWR VPWR _10186_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17160_ _14147_ net3387 _04829_ VGND VGND VPWR VPWR _04838_ sky130_fd_sc_hd__mux2_1
X_29146_ _13089_ VGND VGND VPWR VPWR _04346_ sky130_fd_sc_hd__clkbuf_1
X_23790__375 clknet_1_0__leaf__10205_ VGND VGND VPWR VPWR net501 sky130_fd_sc_hd__inv_2
X_26358_ _11081_ _11511_ VGND VGND VPWR VPWR _11513_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_1022 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16111_ net1939 _13217_ _14396_ VGND VGND VPWR VPWR _14398_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25309_ _10598_ _10898_ _10828_ VGND VGND VPWR VPWR _10899_ sky130_fd_sc_hd__a21oi_4
X_26289_ net1815 _11467_ VGND VGND VPWR VPWR _11477_ sky130_fd_sc_hd__and2_1
X_29077_ _12758_ net3055 _13049_ VGND VGND VPWR VPWR _13053_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17091_ _04801_ VGND VGND VPWR VPWR _01492_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28028_ _12476_ VGND VGND VPWR VPWR _03841_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16042_ _14361_ VGND VGND VPWR VPWR _02001_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19801_ _07071_ _07076_ _07083_ _07095_ VGND VGND VPWR VPWR _07096_ sky130_fd_sc_hd__o31a_1
XFILLER_0_20_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23424__76 clknet_1_0__leaf__10154_ VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__inv_2
XFILLER_0_62_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_208_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17993_ _05321_ rvcpu.dp.SrcBFW_Mux.y\[4\] _05362_ VGND VGND VPWR VPWR _05363_ sky130_fd_sc_hd__o21ai_4
X_29979_ net349 _01714_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[14\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_19732_ datamem.data_ram\[8\]\[25\] _06649_ _07026_ _06603_ VGND VGND VPWR VPWR _07027_
+ sky130_fd_sc_hd__o211a_1
X_16944_ _04723_ VGND VGND VPWR VPWR _01569_ sky130_fd_sc_hd__clkbuf_1
X_23684__280 clknet_1_0__leaf__10194_ VGND VGND VPWR VPWR net406 sky130_fd_sc_hd__inv_2
X_32990_ clknet_leaf_207_clk _04412_ VGND VGND VPWR VPWR datamem.data_ram\[62\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31941_ clknet_leaf_116_clk _03363_ VGND VGND VPWR VPWR datamem.data_ram\[59\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_19663_ datamem.data_ram\[42\]\[0\] _06931_ _06925_ datamem.data_ram\[47\]\[0\] VGND
+ VGND VPWR VPWR _06959_ sky130_fd_sc_hd__a22o_1
XFILLER_0_217_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16875_ net2681 _14426_ _04684_ VGND VGND VPWR VPWR _04687_ sky130_fd_sc_hd__mux2_1
X_18614_ _05675_ _05709_ VGND VGND VPWR VPWR _05972_ sky130_fd_sc_hd__or2_1
X_15826_ _14244_ VGND VGND VPWR VPWR _02108_ sky130_fd_sc_hd__clkbuf_1
X_31872_ clknet_leaf_112_clk _03326_ VGND VGND VPWR VPWR datamem.data_ram\[56\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_19594_ datamem.data_ram\[63\]\[8\] _06670_ _06889_ _06851_ VGND VGND VPWR VPWR _06890_
+ sky130_fd_sc_hd__o211a_1
X_23148__823 clknet_1_1__leaf__10107_ VGND VGND VPWR VPWR net949 sky130_fd_sc_hd__inv_2
XFILLER_0_126_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_220_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18545_ _05704_ _05904_ _05905_ VGND VGND VPWR VPWR _05906_ sky130_fd_sc_hd__a21oi_2
X_30823_ clknet_leaf_203_clk _02558_ VGND VGND VPWR VPWR datamem.data_ram\[44\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_138_clk clknet_5_31__leaf_clk VGND VGND VPWR VPWR clknet_leaf_138_clk
+ sky130_fd_sc_hd__clkbuf_8
X_15757_ _14207_ VGND VGND VPWR VPWR _02148_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_220_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14708_ _13265_ VGND VGND VPWR VPWR _13266_ sky130_fd_sc_hd__clkbuf_8
X_18476_ _05469_ _05475_ _05484_ _05490_ _05769_ _05689_ VGND VGND VPWR VPWR _05838_
+ sky130_fd_sc_hd__mux4_1
X_30754_ clknet_leaf_189_clk _02489_ VGND VGND VPWR VPWR datamem.data_ram\[48\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15688_ _14162_ net4394 _14152_ VGND VGND VPWR VPWR _14163_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_215_5651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_380 rvcpu.dp.plmw.ReadDataW\[29\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_215_5662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_391 net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17427_ _14141_ net3509 _04974_ VGND VGND VPWR VPWR _04980_ sky130_fd_sc_hd__mux2_1
X_23341__979 clknet_1_0__leaf__10136_ VGND VGND VPWR VPWR net1105 sky130_fd_sc_hd__inv_2
XFILLER_0_28_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14639_ _13180_ VGND VGND VPWR VPWR _13214_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_157_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30685_ clknet_leaf_261_clk _02420_ VGND VGND VPWR VPWR datamem.data_ram\[4\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_211_5548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32424_ clknet_leaf_78_clk _03846_ VGND VGND VPWR VPWR datamem.data_ram\[28\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_211_5559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_979 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17358_ _04943_ VGND VGND VPWR VPWR _01359_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_144_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16309_ _14517_ VGND VGND VPWR VPWR _01882_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32355_ clknet_leaf_249_clk _03777_ VGND VGND VPWR VPWR datamem.data_ram\[30\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload300 clknet_1_0__leaf__10205_ VGND VGND VPWR VPWR clkload300/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_181_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17289_ net4248 _13194_ _04902_ VGND VGND VPWR VPWR _04907_ sky130_fd_sc_hd__mux2_1
Xclkload311 clknet_1_0__leaf__10191_ VGND VGND VPWR VPWR clkload311/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_3_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload322 clknet_1_0__leaf__10154_ VGND VGND VPWR VPWR clkload322/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload30 clknet_leaf_20_clk VGND VGND VPWR VPWR clkload30/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_113_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload333 clknet_1_1__leaf__10137_ VGND VGND VPWR VPWR clkload333/Y sky130_fd_sc_hd__clkinvlp_4
X_31306_ clknet_leaf_52_clk _03009_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCPlus4E\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_19028_ _06359_ VGND VGND VPWR VPWR rvcpu.dp.lAuiPCE\[1\] sky130_fd_sc_hd__clkbuf_1
Xclkload41 clknet_leaf_27_clk VGND VGND VPWR VPWR clkload41/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_67_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload344 clknet_1_1__leaf__10124_ VGND VGND VPWR VPWR clkload344/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_207_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23120__797 clknet_1_1__leaf__10105_ VGND VGND VPWR VPWR net923 sky130_fd_sc_hd__inv_2
Xclkload52 clknet_leaf_290_clk VGND VGND VPWR VPWR clkload52/Y sky130_fd_sc_hd__inv_6
Xclkload355 clknet_1_0__leaf__10086_ VGND VGND VPWR VPWR clkload355/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_70_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32286_ clknet_leaf_272_clk _03708_ VGND VGND VPWR VPWR datamem.data_ram\[33\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload63 clknet_leaf_79_clk VGND VGND VPWR VPWR clkload63/Y sky130_fd_sc_hd__clkinv_1
XFILLER_0_3_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload74 clknet_leaf_56_clk VGND VGND VPWR VPWR clkload74/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_144_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload85 clknet_leaf_49_clk VGND VGND VPWR VPWR clkload85/Y sky130_fd_sc_hd__inv_12
XFILLER_0_101_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31237_ clknet_leaf_31_clk _02940_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCD\[26\] sky130_fd_sc_hd__dfxtp_1
Xclkload96 clknet_leaf_83_clk VGND VGND VPWR VPWR clkload96/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_140_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23767__355 clknet_1_1__leaf__10202_ VGND VGND VPWR VPWR net481 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_166_4470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_4481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31168_ clknet_leaf_9_clk rvcpu.ALUResultE\[27\] VGND VGND VPWR VPWR rvcpu.dp.plem.ALUResultM\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23235__884 clknet_1_1__leaf__10125_ VGND VGND VPWR VPWR net1010 sky130_fd_sc_hd__inv_2
Xhold2803 datamem.data_ram\[44\]\[13\] VGND VGND VPWR VPWR net3953 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2814 rvcpu.dp.rf.reg_file_arr\[31\]\[30\] VGND VGND VPWR VPWR net3964 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2825 datamem.data_ram\[48\]\[27\] VGND VGND VPWR VPWR net3975 sky130_fd_sc_hd__dlygate4sd3_1
X_30119_ net481 _01854_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[10\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2836 rvcpu.dp.rf.reg_file_arr\[20\]\[0\] VGND VGND VPWR VPWR net3986 sky130_fd_sc_hd__dlygate4sd3_1
X_23990_ clknet_1_1__leaf__10224_ VGND VGND VPWR VPWR _10240_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_162_4378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2847 rvcpu.dp.rf.reg_file_arr\[25\]\[6\] VGND VGND VPWR VPWR net3997 sky130_fd_sc_hd__dlygate4sd3_1
X_31099_ clknet_leaf_279_clk _02834_ VGND VGND VPWR VPWR datamem.data_ram\[9\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_162_4389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2858 datamem.data_ram\[42\]\[18\] VGND VGND VPWR VPWR net4008 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2869 rvcpu.dp.rf.reg_file_arr\[3\]\[10\] VGND VGND VPWR VPWR net4019 sky130_fd_sc_hd__dlygate4sd3_1
X_22941_ _10069_ VGND VGND VPWR VPWR _10070_ sky130_fd_sc_hd__buf_2
XFILLER_0_98_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_223_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25660_ _10142_ _10921_ _10922_ VGND VGND VPWR VPWR _11098_ sky130_fd_sc_hd__and3_2
X_22872_ _09398_ _10007_ VGND VGND VPWR VPWR _10008_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_175_4706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_214_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24611_ _10476_ net4059 _10502_ VGND VGND VPWR VPWR _10508_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21823_ rvcpu.dp.rf.reg_file_arr\[28\]\[23\] rvcpu.dp.rf.reg_file_arr\[30\]\[23\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[23\] rvcpu.dp.rf.reg_file_arr\[31\]\[23\] _08568_
+ _08683_ VGND VGND VPWR VPWR _09062_ sky130_fd_sc_hd__mux4_1
X_25591_ _10410_ _11055_ VGND VGND VPWR VPWR _11059_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_129_clk clknet_5_31__leaf_clk VGND VGND VPWR VPWR clknet_leaf_129_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_214_1048 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27330_ _10070_ _12076_ _12077_ net1359 VGND VGND VPWR VPWR _03540_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_174_Right_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_121_3396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24542_ _10467_ VGND VGND VPWR VPWR _02364_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21754_ _08813_ _08996_ _08689_ VGND VGND VPWR VPWR _08997_ sky130_fd_sc_hd__a21o_1
XFILLER_0_149_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20705_ datamem.data_ram\[13\]\[5\] _06921_ _07994_ _07995_ VGND VGND VPWR VPWR _07996_
+ sky130_fd_sc_hd__a211o_1
X_27261_ _10070_ net52 _12042_ net1366 VGND VGND VPWR VPWR _03508_ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24473_ _10426_ VGND VGND VPWR VPWR _02336_ sky130_fd_sc_hd__clkbuf_1
X_21685_ _08695_ _08931_ VGND VGND VPWR VPWR _08932_ sky130_fd_sc_hd__and2_1
X_29000_ _10047_ _13010_ VGND VGND VPWR VPWR _13011_ sky130_fd_sc_hd__and2_1
XFILLER_0_149_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_134_3702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26212_ net1705 _11442_ _03041_ _11443_ VGND VGND VPWR VPWR _03058_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_3713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27192_ _11980_ _11996_ VGND VGND VPWR VPWR _12004_ sky130_fd_sc_hd__and2_1
X_20636_ datamem.data_ram\[10\]\[29\] _06610_ _06821_ datamem.data_ram\[8\]\[29\]
+ VGND VGND VPWR VPWR _07927_ sky130_fd_sc_hd__o22a_1
Xclkload2 clknet_5_3__leaf_clk VGND VGND VPWR VPWR clkload2/Y sky130_fd_sc_hd__inv_6
XFILLER_0_151_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26143_ _11407_ VGND VGND VPWR VPWR _03024_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20567_ rvcpu.dp.plem.ALUResultM\[6\] _06860_ VGND VGND VPWR VPWR _07858_ sky130_fd_sc_hd__nor2_4
XFILLER_0_149_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24147__651 clknet_1_1__leaf__10262_ VGND VGND VPWR VPWR net777 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_95_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22306_ _09469_ _09470_ VGND VGND VPWR VPWR _09471_ sky130_fd_sc_hd__or2_1
X_26074_ _08622_ _11367_ VGND VGND VPWR VPWR _11368_ sky130_fd_sc_hd__and2_1
XFILLER_0_132_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23553__177 clknet_1_1__leaf__10174_ VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_95_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20498_ datamem.data_ram\[32\]\[21\] _06649_ _07077_ datamem.data_ram\[35\]\[21\]
+ _07788_ VGND VGND VPWR VPWR _07789_ sky130_fd_sc_hd__o221a_1
XFILLER_0_225_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29902_ clknet_leaf_140_clk _01637_ VGND VGND VPWR VPWR datamem.data_ram\[59\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_25025_ _09287_ VGND VGND VPWR VPWR _10737_ sky130_fd_sc_hd__buf_2
X_22237_ rvcpu.dp.rf.reg_file_arr\[28\]\[0\] rvcpu.dp.rf.reg_file_arr\[30\]\[0\] rvcpu.dp.rf.reg_file_arr\[29\]\[0\]
+ rvcpu.dp.rf.reg_file_arr\[31\]\[0\] _09400_ _09402_ VGND VGND VPWR VPWR _09403_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_104_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23372__1007 clknet_1_0__leaf__10139_ VGND VGND VPWR VPWR net1133 sky130_fd_sc_hd__inv_2
XFILLER_0_218_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29833_ net211 _01568_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[1\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_22168_ _09355_ VGND VGND VPWR VPWR _01102_ sky130_fd_sc_hd__clkbuf_1
X_21119_ _08369_ _08380_ _08407_ VGND VGND VPWR VPWR _08408_ sky130_fd_sc_hd__a21oi_2
X_29764_ net1110 _01499_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[21\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_14990_ rvcpu.dp.pcreg.q\[9\] VGND VGND VPWR VPWR _13538_ sky130_fd_sc_hd__inv_2
X_26976_ _11833_ _11866_ VGND VGND VPWR VPWR _11872_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22099_ _09310_ net3974 _09302_ VGND VGND VPWR VPWR _09311_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28715_ _12856_ VGND VGND VPWR VPWR _04148_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_205_129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25927_ net2078 _11275_ _11273_ _11283_ VGND VGND VPWR VPWR _02933_ sky130_fd_sc_hd__o211a_1
XFILLER_0_191_1107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29695_ net1041 _01430_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[23\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16660_ _04572_ VGND VGND VPWR VPWR _01710_ sky130_fd_sc_hd__clkbuf_1
X_28646_ _12745_ net3068 _12814_ VGND VGND VPWR VPWR _12820_ sky130_fd_sc_hd__mux2_1
X_25858_ _11238_ VGND VGND VPWR VPWR _02909_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15611_ _14113_ VGND VGND VPWR VPWR _02200_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24809_ _10450_ net3929 _10612_ VGND VGND VPWR VPWR _10618_ sky130_fd_sc_hd__mux2_1
X_28577_ _12762_ net2575 _12777_ VGND VGND VPWR VPWR _12783_ sky130_fd_sc_hd__mux2_1
X_16591_ _04535_ VGND VGND VPWR VPWR _01750_ sky130_fd_sc_hd__clkbuf_1
X_25789_ _11182_ _11183_ _11149_ VGND VGND VPWR VPWR _11184_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_201_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18330_ _05678_ _05691_ _05694_ VGND VGND VPWR VPWR _05695_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15542_ _13374_ _14066_ _14067_ _13513_ VGND VGND VPWR VPWR _14068_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_141_Right_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27528_ _12095_ net1894 _12188_ VGND VGND VPWR VPWR _12196_ sky130_fd_sc_hd__mux2_1
XFILLER_0_189_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18261_ rvcpu.dp.plde.RD1E\[22\] _05564_ _05462_ VGND VGND VPWR VPWR _05626_ sky130_fd_sc_hd__o21ai_2
X_15473_ _14002_ VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__inv_2
XFILLER_0_38_952 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27459_ _12158_ VGND VGND VPWR VPWR _03590_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_182_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_1312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17212_ _14127_ net2387 _04865_ VGND VGND VPWR VPWR _04866_ sky130_fd_sc_hd__mux2_1
X_18192_ _05302_ _05556_ VGND VGND VPWR VPWR _05557_ sky130_fd_sc_hd__nor2_1
X_30470_ net148 _02205_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[19\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_730 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29129_ _13080_ VGND VGND VPWR VPWR _04338_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17143_ _04828_ VGND VGND VPWR VPWR _04829_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_13_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23178__849 clknet_1_1__leaf__10111_ VGND VGND VPWR VPWR net975 sky130_fd_sc_hd__inv_2
XFILLER_0_53_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32140_ clknet_leaf_256_clk _03562_ VGND VGND VPWR VPWR datamem.data_ram\[39\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold709 rvcpu.dp.pcreg.q\[24\] VGND VGND VPWR VPWR net1859 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17074_ _14128_ _04755_ VGND VGND VPWR VPWR _04792_ sky130_fd_sc_hd__nand2_4
XFILLER_0_126_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_690 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16025_ _14352_ VGND VGND VPWR VPWR _02009_ sky130_fd_sc_hd__clkbuf_1
X_32071_ clknet_leaf_121_clk _03493_ VGND VGND VPWR VPWR datamem.data_ram\[29\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31022_ clknet_leaf_60_clk _02757_ VGND VGND VPWR VPWR datamem.data_ram\[40\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17976_ rvcpu.dp.plem.ALUResultM\[6\] VGND VGND VPWR VPWR _05347_ sky130_fd_sc_hd__inv_6
Xhold1409 rvcpu.dp.rf.reg_file_arr\[5\]\[26\] VGND VGND VPWR VPWR net2559 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19715_ datamem.data_ram\[24\]\[0\] _06936_ _06942_ datamem.data_ram\[27\]\[0\] _06769_
+ VGND VGND VPWR VPWR _07011_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_204_5385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_204_5396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16927_ net1883 _14478_ _04706_ VGND VGND VPWR VPWR _04714_ sky130_fd_sc_hd__mux2_1
X_32973_ clknet_leaf_145_clk _04395_ VGND VGND VPWR VPWR datamem.data_ram\[63\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19646_ _06941_ VGND VGND VPWR VPWR _06942_ sky130_fd_sc_hd__buf_4
X_31924_ _04436_ net118 VGND VGND VPWR VPWR datamem.rd_data_mem\[29\] sky130_fd_sc_hd__dlxtn_1
XFILLER_0_79_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16858_ _04677_ VGND VGND VPWR VPWR _01609_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_215_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_217_5702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_196_5197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_217_5713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15809_ _14090_ _14234_ VGND VGND VPWR VPWR _14235_ sky130_fd_sc_hd__nor2_2
X_31855_ clknet_leaf_125_clk _03309_ VGND VGND VPWR VPWR datamem.data_ram\[62\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_19577_ datamem.data_ram\[10\]\[8\] _06754_ _06871_ _06872_ VGND VGND VPWR VPWR _06873_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_215_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16789_ net3424 _14476_ _04634_ VGND VGND VPWR VPWR _04641_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_1110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30806_ clknet_leaf_137_clk _02541_ VGND VGND VPWR VPWR datamem.data_ram\[45\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_18528_ _05866_ _05805_ VGND VGND VPWR VPWR _05889_ sky130_fd_sc_hd__nor2_1
XFILLER_0_133_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31786_ clknet_leaf_53_clk _03240_ VGND VGND VPWR VPWR datamem.data_ram\[8\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_24016__548 clknet_1_1__leaf__10242_ VGND VGND VPWR VPWR net674 sky130_fd_sc_hd__inv_2
XFILLER_0_220_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18459_ _05622_ _05574_ _05570_ _05565_ _05682_ _05579_ VGND VGND VPWR VPWR _05822_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_118_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30737_ clknet_leaf_219_clk _02472_ VGND VGND VPWR VPWR datamem.data_ram\[47\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21470_ _08725_ _08726_ VGND VGND VPWR VPWR _08727_ sky130_fd_sc_hd__nor2_1
X_30668_ clknet_leaf_130_clk _02403_ VGND VGND VPWR VPWR datamem.data_ram\[50\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_356 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32407_ clknet_leaf_274_clk _03829_ VGND VGND VPWR VPWR datamem.data_ram\[29\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_20421_ _06751_ _07707_ _07712_ VGND VGND VPWR VPWR _07713_ sky130_fd_sc_hd__or3_1
XFILLER_0_16_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23472__120 clknet_1_0__leaf__10158_ VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__inv_2
XFILLER_0_132_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30599_ clknet_leaf_197_clk _02334_ VGND VGND VPWR VPWR datamem.data_ram\[53\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20352_ _07633_ _07638_ _07643_ _06716_ VGND VGND VPWR VPWR _07644_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_168_4521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32338_ clknet_leaf_239_clk _03760_ VGND VGND VPWR VPWR datamem.data_ram\[30\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload130 clknet_leaf_258_clk VGND VGND VPWR VPWR clkload130/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_168_4532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload141 clknet_leaf_246_clk VGND VGND VPWR VPWR clkload141/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload152 clknet_leaf_275_clk VGND VGND VPWR VPWR clkload152/Y sky130_fd_sc_hd__clkinv_4
Xclkload163 clknet_leaf_183_clk VGND VGND VPWR VPWR clkload163/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_222_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload174 clknet_leaf_229_clk VGND VGND VPWR VPWR clkload174/Y sky130_fd_sc_hd__bufinv_16
X_23071_ _10097_ VGND VGND VPWR VPWR _01263_ sky130_fd_sc_hd__clkbuf_1
X_20283_ datamem.data_ram\[30\]\[19\] _06763_ _06699_ datamem.data_ram\[25\]\[19\]
+ VGND VGND VPWR VPWR _07576_ sky130_fd_sc_hd__o22a_1
X_32269_ clknet_leaf_223_clk _03691_ VGND VGND VPWR VPWR datamem.data_ram\[33\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload185 clknet_leaf_218_clk VGND VGND VPWR VPWR clkload185/Y sky130_fd_sc_hd__bufinv_16
Xclkload196 clknet_leaf_186_clk VGND VGND VPWR VPWR clkload196/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_164_4429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3301 rvcpu.dp.plfd.InstrD\[7\] VGND VGND VPWR VPWR net4451 sky130_fd_sc_hd__dlygate4sd3_1
X_22022_ _09247_ VGND VGND VPWR VPWR _09248_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_90_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2600 rvcpu.dp.rf.reg_file_arr\[15\]\[8\] VGND VGND VPWR VPWR net3750 sky130_fd_sc_hd__dlygate4sd3_1
X_26830_ _11752_ VGND VGND VPWR VPWR _11781_ sky130_fd_sc_hd__buf_2
Xhold2611 datamem.data_ram\[10\]\[10\] VGND VGND VPWR VPWR net3761 sky130_fd_sc_hd__dlygate4sd3_1
X_23016__720 clknet_1_1__leaf__10086_ VGND VGND VPWR VPWR net846 sky130_fd_sc_hd__inv_2
Xhold14 rvcpu.dp.plem.lAuiPCM\[25\] VGND VGND VPWR VPWR net1164 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2622 datamem.data_ram\[24\]\[26\] VGND VGND VPWR VPWR net3772 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2633 rvcpu.dp.rf.reg_file_arr\[10\]\[14\] VGND VGND VPWR VPWR net3783 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 rvcpu.dp.plde.PCPlus4E\[31\] VGND VGND VPWR VPWR net1175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2644 rvcpu.dp.rf.reg_file_arr\[25\]\[2\] VGND VGND VPWR VPWR net3794 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 rvcpu.dp.plde.PCPlus4E\[9\] VGND VGND VPWR VPWR net1186 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_127_3550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1910 datamem.data_ram\[1\]\[30\] VGND VGND VPWR VPWR net3060 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 rvcpu.dp.plem.PCPlus4M\[23\] VGND VGND VPWR VPWR net1197 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2655 datamem.data_ram\[17\]\[11\] VGND VGND VPWR VPWR net3805 sky130_fd_sc_hd__dlygate4sd3_1
X_26761_ _11735_ net1754 _11737_ _11740_ VGND VGND VPWR VPWR _03310_ sky130_fd_sc_hd__a31o_1
Xhold2666 datamem.data_ram\[32\]\[21\] VGND VGND VPWR VPWR net3816 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 rvcpu.dp.plde.MemWriteE VGND VGND VPWR VPWR net1208 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1921 rvcpu.dp.rf.reg_file_arr\[27\]\[9\] VGND VGND VPWR VPWR net3071 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold69 rvcpu.dp.plde.PCPlus4E\[27\] VGND VGND VPWR VPWR net1219 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1932 rvcpu.dp.rf.reg_file_arr\[31\]\[26\] VGND VGND VPWR VPWR net3082 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2677 rvcpu.dp.rf.reg_file_arr\[15\]\[0\] VGND VGND VPWR VPWR net3827 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_67_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1943 datamem.data_ram\[24\]\[24\] VGND VGND VPWR VPWR net3093 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2688 datamem.data_ram\[12\]\[28\] VGND VGND VPWR VPWR net3838 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_123_3436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2699 rvcpu.dp.rf.reg_file_arr\[27\]\[15\] VGND VGND VPWR VPWR net3849 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1954 rvcpu.dp.rf.reg_file_arr\[30\]\[21\] VGND VGND VPWR VPWR net3104 sky130_fd_sc_hd__dlygate4sd3_1
X_28500_ _12279_ _10092_ _12668_ VGND VGND VPWR VPWR _12735_ sky130_fd_sc_hd__a21oi_4
X_25712_ _11129_ VGND VGND VPWR VPWR _02872_ sky130_fd_sc_hd__clkbuf_1
Xhold1965 datamem.data_ram\[40\]\[10\] VGND VGND VPWR VPWR net3115 sky130_fd_sc_hd__dlygate4sd3_1
X_22924_ rvcpu.dp.plem.WriteDataM\[1\] VGND VGND VPWR VPWR _10057_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_123_3447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29480_ net842 _01215_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[2\]\[19\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__10261_ clknet_0__10261_ VGND VGND VPWR VPWR clknet_1_1__leaf__10261_
+ sky130_fd_sc_hd__clkbuf_16
X_26692_ _11104_ VGND VGND VPWR VPWR _11700_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_123_3458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1976 datamem.data_ram\[3\]\[24\] VGND VGND VPWR VPWR net3126 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_600 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1987 datamem.data_ram\[16\]\[28\] VGND VGND VPWR VPWR net3137 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1998 datamem.data_ram\[3\]\[27\] VGND VGND VPWR VPWR net3148 sky130_fd_sc_hd__dlygate4sd3_1
X_28431_ _12694_ net3956 _12688_ VGND VGND VPWR VPWR _12695_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25643_ _10072_ VGND VGND VPWR VPWR _11091_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_151_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22855_ rvcpu.dp.rf.reg_file_arr\[24\]\[29\] rvcpu.dp.rf.reg_file_arr\[25\]\[29\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[29\] rvcpu.dp.rf.reg_file_arr\[27\]\[29\] _08592_
+ _09394_ VGND VGND VPWR VPWR _09992_ sky130_fd_sc_hd__mux4_1
Xclkbuf_1_1__f__10192_ clknet_0__10192_ VGND VGND VPWR VPWR clknet_1_1__leaf__10192_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_210_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28362_ _12458_ net3603 _12650_ VGND VGND VPWR VPWR _12656_ sky130_fd_sc_hd__mux2_1
X_21806_ _08798_ _09043_ _09045_ _08512_ VGND VGND VPWR VPWR _09046_ sky130_fd_sc_hd__o211a_1
X_25574_ _11047_ _11042_ VGND VGND VPWR VPWR _11048_ sky130_fd_sc_hd__and2_1
X_22786_ _09441_ _09926_ VGND VGND VPWR VPWR _09927_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_26_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27313_ _12061_ net1584 _12065_ _12071_ VGND VGND VPWR VPWR _03531_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_26_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24525_ _10388_ datamem.data_ram\[52\]\[9\] _10456_ VGND VGND VPWR VPWR _10458_ sky130_fd_sc_hd__mux2_1
X_21737_ _08663_ _08978_ _08980_ _08558_ VGND VGND VPWR VPWR _08981_ sky130_fd_sc_hd__o211a_1
X_28293_ _12441_ net3871 _12613_ VGND VGND VPWR VPWR _12619_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23936__491 clknet_1_1__leaf__10227_ VGND VGND VPWR VPWR net617 sky130_fd_sc_hd__inv_2
XFILLER_0_213_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27244_ _12022_ net1648 _12030_ _12035_ VGND VGND VPWR VPWR _03498_ sky130_fd_sc_hd__a31o_1
XFILLER_0_191_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_97_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24456_ _10416_ _10406_ VGND VGND VPWR VPWR _10417_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21668_ _08672_ _08907_ _08911_ _08915_ VGND VGND VPWR VPWR _08916_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_97_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20619_ datamem.data_ram\[12\]\[13\] datamem.data_ram\[13\]\[13\] _07874_ VGND VGND
+ VPWR VPWR _07910_ sky130_fd_sc_hd__mux2_1
X_27175_ _07028_ _11109_ _11839_ VGND VGND VPWR VPWR _11994_ sky130_fd_sc_hd__or3_1
XFILLER_0_151_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24387_ _10372_ VGND VGND VPWR VPWR _02304_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_10_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21599_ rvcpu.dp.rf.reg_file_arr\[28\]\[11\] rvcpu.dp.rf.reg_file_arr\[30\]\[11\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[11\] rvcpu.dp.rf.reg_file_arr\[31\]\[11\] _08559_
+ _08636_ VGND VGND VPWR VPWR _08850_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_10_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26126_ net1765 _11397_ VGND VGND VPWR VPWR _11399_ sky130_fd_sc_hd__and2_1
XFILLER_0_132_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26057_ _11353_ net1525 _11350_ _11357_ VGND VGND VPWR VPWR _02989_ sky130_fd_sc_hd__a31o_1
X_23269_ clknet_1_0__leaf__10108_ VGND VGND VPWR VPWR _10129_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_56_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25008_ _10724_ net3184 net100 VGND VGND VPWR VPWR _10726_ sky130_fd_sc_hd__mux2_1
X_17830_ _05214_ VGND VGND VPWR VPWR rvcpu.dp.SrcBFW_Mux.y\[23\] sky130_fd_sc_hd__clkbuf_2
X_29816_ net194 _01551_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[1\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_210_Right_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_206_438 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17761_ _13174_ rvcpu.dp.plde.Rs2E\[2\] VGND VGND VPWR VPWR _05159_ sky130_fd_sc_hd__xnor2_1
X_29747_ net1093 _01482_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[21\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_23978__514 clknet_1_1__leaf__10238_ VGND VGND VPWR VPWR net640 sky130_fd_sc_hd__inv_2
X_26959_ _11849_ net1354 _11853_ _11861_ VGND VGND VPWR VPWR _03387_ sky130_fd_sc_hd__a31o_1
X_14973_ _13502_ _13516_ _13520_ _13521_ VGND VGND VPWR VPWR _13522_ sky130_fd_sc_hd__a31o_1
XFILLER_0_215_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19500_ rvcpu.dp.plem.ALUResultM\[7\] _06750_ VGND VGND VPWR VPWR _06796_ sky130_fd_sc_hd__nor2_8
XFILLER_0_215_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16712_ _04600_ VGND VGND VPWR VPWR _01686_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17692_ _05120_ VGND VGND VPWR VPWR _01194_ sky130_fd_sc_hd__clkbuf_1
X_29678_ net1024 _01413_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[23\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_214_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_1079 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19431_ datamem.data_ram\[39\]\[16\] _06726_ _06699_ datamem.data_ram\[33\]\[16\]
+ VGND VGND VPWR VPWR _06727_ sky130_fd_sc_hd__o22a_1
XFILLER_0_187_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28629_ _12762_ net3069 _12805_ VGND VGND VPWR VPWR _12811_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16643_ _14175_ net4057 _04562_ VGND VGND VPWR VPWR _04564_ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31640_ clknet_leaf_45_clk net1165 VGND VGND VPWR VPWR rvcpu.dp.plmw.lAuiPCW\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_19362_ _06657_ VGND VGND VPWR VPWR _06658_ sky130_fd_sc_hd__buf_8
X_16574_ _14175_ net4135 _04525_ VGND VGND VPWR VPWR _04527_ sky130_fd_sc_hd__mux2_1
X_23796__381 clknet_1_1__leaf__10205_ VGND VGND VPWR VPWR net507 sky130_fd_sc_hd__inv_2
XFILLER_0_70_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_191_5072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_191_5083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18313_ _05672_ _05673_ _05677_ VGND VGND VPWR VPWR _05678_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15525_ _13413_ _14042_ _14045_ _14051_ VGND VGND VPWR VPWR _14052_ sky130_fd_sc_hd__a211o_1
XFILLER_0_31_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31571_ clknet_leaf_62_clk datamem.rd_data_mem\[21\] VGND VGND VPWR VPWR rvcpu.dp.plmw.ReadDataW\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_19293_ _06586_ _06588_ VGND VGND VPWR VPWR _06589_ sky130_fd_sc_hd__and2_1
XFILLER_0_57_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30522_ clknet_leaf_138_clk _02257_ VGND VGND VPWR VPWR datamem.data_ram\[56\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_18244_ _05410_ _05418_ _05605_ _05608_ VGND VGND VPWR VPWR _05609_ sky130_fd_sc_hd__o31a_1
XFILLER_0_155_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15456_ _13823_ _13747_ _13929_ VGND VGND VPWR VPWR _13986_ sky130_fd_sc_hd__or3_1
XFILLER_0_143_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18175_ rvcpu.dp.plde.ImmExtE\[27\] rvcpu.dp.SrcBFW_Mux.y\[27\] _05279_ VGND VGND
+ VPWR VPWR _05540_ sky130_fd_sc_hd__mux2_1
X_30453_ net131 _02188_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[19\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_15387_ _13309_ _13581_ _13451_ VGND VGND VPWR VPWR _13920_ sky130_fd_sc_hd__or3b_1
XFILLER_0_136_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17126_ _14181_ net2652 _04815_ VGND VGND VPWR VPWR _04820_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_4090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold506 datamem.data_ram\[57\]\[7\] VGND VGND VPWR VPWR net1656 sky130_fd_sc_hd__dlygate4sd3_1
X_30384_ clknet_leaf_268_clk _02119_ VGND VGND VPWR VPWR datamem.data_ram\[58\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold517 datamem.data_ram\[6\]\[1\] VGND VGND VPWR VPWR net1667 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold528 datamem.data_ram\[16\]\[2\] VGND VGND VPWR VPWR net1678 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32123_ clknet_leaf_211_clk _03545_ VGND VGND VPWR VPWR datamem.data_ram\[7\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold539 datamem.data_ram\[15\]\[3\] VGND VGND VPWR VPWR net1689 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17057_ _04783_ VGND VGND VPWR VPWR _01508_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_208_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16008_ net1906 _13269_ _14333_ VGND VGND VPWR VPWR _14342_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_206_5436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32054_ clknet_leaf_121_clk _03476_ VGND VGND VPWR VPWR datamem.data_ram\[30\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_206_5447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31005_ clknet_leaf_162_clk _02740_ VGND VGND VPWR VPWR datamem.data_ram\[11\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_198_5237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1206 datamem.data_ram\[16\]\[31\] VGND VGND VPWR VPWR net2356 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_198_5248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1217 rvcpu.dp.rf.reg_file_arr\[13\]\[16\] VGND VGND VPWR VPWR net2367 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_198_5259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17959_ rvcpu.dp.plde.ImmExtE\[12\] rvcpu.dp.SrcBFW_Mux.y\[12\] _05277_ VGND VGND
+ VPWR VPWR _05330_ sky130_fd_sc_hd__mux2_1
Xhold1228 rvcpu.dp.rf.reg_file_arr\[18\]\[19\] VGND VGND VPWR VPWR net2378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1239 rvcpu.dp.rf.reg_file_arr\[18\]\[10\] VGND VGND VPWR VPWR net2389 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_213_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32956_ clknet_leaf_99_clk _04378_ VGND VGND VPWR VPWR datamem.data_ram\[6\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_20970_ datamem.data_ram\[34\]\[15\] _07911_ _08258_ _06607_ VGND VGND VPWR VPWR
+ _08259_ sky130_fd_sc_hd__o211a_1
XFILLER_0_212_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31907_ _04418_ net119 VGND VGND VPWR VPWR datamem.rd_data_mem\[12\] sky130_fd_sc_hd__dlxtn_1
X_19629_ _06924_ VGND VGND VPWR VPWR _06925_ sky130_fd_sc_hd__buf_4
XFILLER_0_189_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32887_ clknet_leaf_279_clk _04309_ VGND VGND VPWR VPWR datamem.data_ram\[10\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_23504__149 clknet_1_0__leaf__10161_ VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__inv_2
X_22640_ _09387_ VGND VGND VPWR VPWR _09789_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_157_4255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31838_ clknet_leaf_209_clk _03292_ VGND VGND VPWR VPWR datamem.data_ram\[3\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_211_1029 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_4266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23371__1006 clknet_1_0__leaf__10139_ VGND VGND VPWR VPWR net1132 sky130_fd_sc_hd__inv_2
XFILLER_0_177_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23046__746 clknet_1_0__leaf__10090_ VGND VGND VPWR VPWR net872 sky130_fd_sc_hd__inv_2
X_22571_ _09627_ _09720_ _09723_ _09438_ VGND VGND VPWR VPWR _09724_ sky130_fd_sc_hd__a211o_1
XFILLER_0_8_610 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31769_ clknet_leaf_210_clk _03223_ VGND VGND VPWR VPWR datamem.data_ram\[1\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_60_clk clknet_5_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_60_clk sky130_fd_sc_hd__clkbuf_8
X_24310_ _10330_ VGND VGND VPWR VPWR _02269_ sky130_fd_sc_hd__clkbuf_1
X_21522_ _08768_ _08772_ _08776_ _08625_ VGND VGND VPWR VPWR _01035_ sky130_fd_sc_hd__o31a_1
XFILLER_0_180_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25290_ _10751_ net2701 _10887_ VGND VGND VPWR VPWR _10888_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24241_ _09279_ net2715 _10288_ VGND VGND VPWR VPWR _10292_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21453_ _08627_ _08706_ _08708_ _08710_ VGND VGND VPWR VPWR _08711_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_17_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_3284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20404_ datamem.data_ram\[35\]\[12\] _06737_ _06782_ datamem.data_ram\[33\]\[12\]
+ _07695_ VGND VGND VPWR VPWR _07696_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_92_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21384_ rvcpu.dp.rf.reg_file_arr\[0\]\[1\] rvcpu.dp.rf.reg_file_arr\[1\]\[1\] rvcpu.dp.rf.reg_file_arr\[2\]\[1\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[1\] _08550_ _08554_ VGND VGND VPWR VPWR _08645_ sky130_fd_sc_hd__mux4_1
XFILLER_0_43_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20335_ datamem.data_ram\[34\]\[4\] _06930_ _06941_ datamem.data_ram\[35\]\[4\] VGND
+ VGND VPWR VPWR _07627_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_187_4974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_187_4985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28980_ _10141_ _10997_ _12977_ VGND VGND VPWR VPWR _12999_ sky130_fd_sc_hd__a21oi_4
Xoutput15 net15 VGND VGND VPWR VPWR Instr[21] sky130_fd_sc_hd__buf_2
Xoutput26 net26 VGND VGND VPWR VPWR Instr[31] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_129_3601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27931_ _12417_ VGND VGND VPWR VPWR _03803_ sky130_fd_sc_hd__clkbuf_1
X_20266_ datamem.data_ram\[58\]\[19\] _06691_ _06768_ datamem.data_ram\[61\]\[19\]
+ VGND VGND VPWR VPWR _07559_ sky130_fd_sc_hd__o22a_1
XFILLER_0_12_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold3120 datamem.data_ram\[18\]\[12\] VGND VGND VPWR VPWR net4270 sky130_fd_sc_hd__dlygate4sd3_1
X_22005_ rvcpu.dp.plem.WriteDataM\[17\] _09221_ VGND VGND VPWR VPWR _09234_ sky130_fd_sc_hd__and2_1
Xhold3131 rvcpu.dp.rf.reg_file_arr\[0\]\[16\] VGND VGND VPWR VPWR net4281 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3142 datamem.data_ram\[39\]\[20\] VGND VGND VPWR VPWR net4292 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3153 rvcpu.dp.plem.ALUResultM\[4\] VGND VGND VPWR VPWR net4303 sky130_fd_sc_hd__dlygate4sd3_1
X_27862_ _12379_ VGND VGND VPWR VPWR _03772_ sky130_fd_sc_hd__clkbuf_1
X_20197_ datamem.data_ram\[32\]\[11\] _06778_ _06737_ datamem.data_ram\[35\]\[11\]
+ _06769_ VGND VGND VPWR VPWR _07490_ sky130_fd_sc_hd__o221a_1
Xhold3164 rvcpu.dp.rf.reg_file_arr\[16\]\[29\] VGND VGND VPWR VPWR net4314 sky130_fd_sc_hd__dlygate4sd3_1
X_29601_ net955 _01336_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[25\]\[4\] sky130_fd_sc_hd__dfxtp_1
Xhold2430 datamem.data_ram\[48\]\[9\] VGND VGND VPWR VPWR net3580 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3175 datamem.data_ram\[19\]\[10\] VGND VGND VPWR VPWR net4325 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26813_ _11672_ _11762_ VGND VGND VPWR VPWR _11771_ sky130_fd_sc_hd__and2_1
Xhold3186 datamem.data_ram\[62\]\[17\] VGND VGND VPWR VPWR net4336 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2441 datamem.data_ram\[0\]\[19\] VGND VGND VPWR VPWR net3591 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3197 datamem.data_ram\[20\]\[23\] VGND VGND VPWR VPWR net4347 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2452 rvcpu.dp.rf.reg_file_arr\[14\]\[17\] VGND VGND VPWR VPWR net3602 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27793_ _12338_ VGND VGND VPWR VPWR _03744_ sky130_fd_sc_hd__clkbuf_1
Xhold2463 datamem.data_ram\[8\]\[15\] VGND VGND VPWR VPWR net3613 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_146_3992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2474 datamem.data_ram\[51\]\[31\] VGND VGND VPWR VPWR net3624 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29532_ clknet_leaf_173_clk _01267_ VGND VGND VPWR VPWR datamem.data_ram\[5\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1740 datamem.data_ram\[22\]\[28\] VGND VGND VPWR VPWR net2890 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2485 datamem.data_ram\[33\]\[8\] VGND VGND VPWR VPWR net3635 sky130_fd_sc_hd__dlygate4sd3_1
X_26744_ _11684_ _11726_ VGND VGND VPWR VPWR _11730_ sky130_fd_sc_hd__and2_1
Xhold2496 datamem.data_ram\[42\]\[16\] VGND VGND VPWR VPWR net3646 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1751 datamem.data_ram\[47\]\[31\] VGND VGND VPWR VPWR net2901 sky130_fd_sc_hd__dlygate4sd3_1
X_23956_ _09240_ net4374 _10229_ VGND VGND VPWR VPWR _10232_ sky130_fd_sc_hd__mux2_1
Xhold1762 datamem.data_ram\[40\]\[25\] VGND VGND VPWR VPWR net2912 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_86_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1773 rvcpu.dp.rf.reg_file_arr\[27\]\[21\] VGND VGND VPWR VPWR net2923 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1784 rvcpu.dp.rf.reg_file_arr\[27\]\[20\] VGND VGND VPWR VPWR net2934 sky130_fd_sc_hd__dlygate4sd3_1
X_22907_ _06587_ VGND VGND VPWR VPWR _10041_ sky130_fd_sc_hd__buf_4
X_29463_ net825 _01198_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[2\]\[2\] sky130_fd_sc_hd__dfxtp_1
Xhold1795 rvcpu.dp.rf.reg_file_arr\[8\]\[27\] VGND VGND VPWR VPWR net2945 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f__10244_ clknet_0__10244_ VGND VGND VPWR VPWR clknet_1_1__leaf__10244_
+ sky130_fd_sc_hd__clkbuf_16
X_26675_ _11689_ _11677_ VGND VGND VPWR VPWR _11690_ sky130_fd_sc_hd__and2_1
XFILLER_0_54_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_211_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28414_ _12458_ net3940 _12678_ VGND VGND VPWR VPWR _12684_ sky130_fd_sc_hd__mux2_1
X_25626_ _11078_ _11079_ VGND VGND VPWR VPWR _11080_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29394_ clknet_leaf_1_clk _01129_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD2E\[5\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__10175_ clknet_0__10175_ VGND VGND VPWR VPWR clknet_1_1__leaf__10175_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_49_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22838_ _09495_ _09975_ _09472_ VGND VGND VPWR VPWR _09976_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_196_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23479__126 clknet_1_0__leaf__10159_ VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__inv_2
XFILLER_0_6_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28345_ _12441_ net4007 _12641_ VGND VGND VPWR VPWR _12647_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25557_ _10764_ net4101 _11030_ VGND VGND VPWR VPWR _11037_ sky130_fd_sc_hd__mux2_1
X_22769_ rvcpu.dp.rf.reg_file_arr\[4\]\[24\] rvcpu.dp.rf.reg_file_arr\[5\]\[24\] rvcpu.dp.rf.reg_file_arr\[6\]\[24\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[24\] _09416_ _09716_ VGND VGND VPWR VPWR _09911_
+ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_51_clk clknet_5_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_51_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_45_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15310_ _13414_ _13562_ VGND VGND VPWR VPWR _13847_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24508_ _10446_ datamem.data_ram\[52\]\[19\] _10440_ VGND VGND VPWR VPWR _10447_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28276_ _12609_ VGND VGND VPWR VPWR _03956_ sky130_fd_sc_hd__clkbuf_1
X_23559__183 clknet_1_1__leaf__10174_ VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__inv_2
X_16290_ _14507_ VGND VGND VPWR VPWR _01891_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25488_ _10500_ VGND VGND VPWR VPWR _10998_ sky130_fd_sc_hd__buf_8
XFILLER_0_93_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15241_ _13721_ _13780_ VGND VGND VPWR VPWR _13781_ sky130_fd_sc_hd__nand2_1
X_27227_ _12022_ net1606 _12018_ _12025_ VGND VGND VPWR VPWR _03491_ sky130_fd_sc_hd__a31o_1
XFILLER_0_191_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24439_ _10047_ VGND VGND VPWR VPWR _10405_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_124_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15172_ _13509_ _13294_ _13607_ VGND VGND VPWR VPWR _13715_ sky130_fd_sc_hd__a21o_1
X_27158_ _11965_ _11984_ VGND VGND VPWR VPWR _11985_ sky130_fd_sc_hd__and2_1
XFILLER_0_205_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26109_ net1376 _11386_ VGND VGND VPWR VPWR _11390_ sky130_fd_sc_hd__and2_1
XFILLER_0_133_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19980_ _06752_ _07268_ _07273_ VGND VGND VPWR VPWR _07274_ sky130_fd_sc_hd__or3_1
XFILLER_0_120_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_205_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27089_ _11939_ VGND VGND VPWR VPWR _11940_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_619 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18931_ _05456_ _05463_ _05665_ VGND VGND VPWR VPWR _06270_ sky130_fd_sc_hd__mux2_1
X_24045__574 clknet_1_1__leaf__10245_ VGND VGND VPWR VPWR net700 sky130_fd_sc_hd__inv_2
XFILLER_0_197_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_219_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18862_ _06200_ _06204_ _06205_ VGND VGND VPWR VPWR _06206_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_1186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_201_5311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17813_ _13189_ rvcpu.dp.plde.RD2E\[28\] _05196_ VGND VGND VPWR VPWR _05203_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_201_5322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18793_ _05313_ _05320_ _05506_ _05334_ _05670_ _05769_ VGND VGND VPWR VPWR _06141_
+ sky130_fd_sc_hd__mux4_1
X_32810_ clknet_leaf_285_clk _04232_ VGND VGND VPWR VPWR datamem.data_ram\[13\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_17744_ _05147_ VGND VGND VPWR VPWR _01169_ sky130_fd_sc_hd__clkbuf_1
X_14956_ _13284_ _13300_ VGND VGND VPWR VPWR _13505_ sky130_fd_sc_hd__nor2_4
XFILLER_0_221_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_178_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_193_5123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_193_5134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32741_ clknet_leaf_287_clk _04163_ VGND VGND VPWR VPWR datamem.data_ram\[16\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_17675_ net2677 _13262_ _05104_ VGND VGND VPWR VPWR _05111_ sky130_fd_sc_hd__mux2_1
X_14887_ _13438_ VGND VGND VPWR VPWR _13439_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19414_ _06681_ _06694_ _06709_ VGND VGND VPWR VPWR _06710_ sky130_fd_sc_hd__and3_1
XFILLER_0_202_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16626_ _14158_ net2422 _04551_ VGND VGND VPWR VPWR _04555_ sky130_fd_sc_hd__mux2_1
X_32672_ clknet_leaf_284_clk _04094_ VGND VGND VPWR VPWR datamem.data_ram\[19\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_31623_ clknet_leaf_65_clk net1206 VGND VGND VPWR VPWR rvcpu.dp.plmw.lAuiPCW\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_19345_ _06591_ _06622_ VGND VGND VPWR VPWR _06641_ sky130_fd_sc_hd__nor2_8
XFILLER_0_175_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16557_ _14158_ net2536 _04514_ VGND VGND VPWR VPWR _04518_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_42_clk clknet_5_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_42_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_223_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15508_ _13542_ _13372_ _13510_ _14033_ _14034_ VGND VGND VPWR VPWR _14035_ sky130_fd_sc_hd__o311a_1
X_31554_ clknet_leaf_62_clk datamem.rd_data_mem\[4\] VGND VGND VPWR VPWR rvcpu.dp.plmw.ReadDataW\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_19276_ rvcpu.dp.plfd.InstrD\[14\] rvcpu.c.ad.opb5 VGND VGND VPWR VPWR _06575_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_152_4141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16488_ _04481_ VGND VGND VPWR VPWR _01799_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_152_4152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18227_ _05587_ _05359_ VGND VGND VPWR VPWR _05592_ sky130_fd_sc_hd__nor2_1
XFILLER_0_155_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30505_ clknet_leaf_267_clk _02240_ VGND VGND VPWR VPWR datamem.data_ram\[57\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_15439_ _13692_ _13389_ _13465_ VGND VGND VPWR VPWR _13970_ sky130_fd_sc_hd__a21oi_1
X_31485_ clknet_leaf_48_clk rvcpu.dp.lAuiPCE\[11\] VGND VGND VPWR VPWR rvcpu.dp.plem.lAuiPCM\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18158_ _05461_ _05467_ _05521_ _05522_ VGND VGND VPWR VPWR _05523_ sky130_fd_sc_hd__a31o_1
X_30436_ net774 _02171_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[29\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold303 datamem.data_ram\[56\]\[5\] VGND VGND VPWR VPWR net1453 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__10264_ clknet_0__10264_ VGND VGND VPWR VPWR clknet_1_0__leaf__10264_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_41_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_390 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold314 datamem.data_ram\[39\]\[7\] VGND VGND VPWR VPWR net1464 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17109_ _14164_ net3031 _04804_ VGND VGND VPWR VPWR _04811_ sky130_fd_sc_hd__mux2_1
Xhold325 datamem.data_ram\[23\]\[4\] VGND VGND VPWR VPWR net1475 sky130_fd_sc_hd__dlygate4sd3_1
X_18089_ rvcpu.dp.plde.ImmExtE\[23\] rvcpu.dp.SrcBFW_Mux.y\[23\] _05278_ VGND VGND
+ VPWR VPWR _05457_ sky130_fd_sc_hd__mux2_1
X_30367_ net713 _02102_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[3\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_229_5981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold336 datamem.data_ram\[50\]\[1\] VGND VGND VPWR VPWR net1486 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_229_5992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold347 datamem.data_ram\[28\]\[1\] VGND VGND VPWR VPWR net1497 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__10195_ clknet_0__10195_ VGND VGND VPWR VPWR clknet_1_0__leaf__10195_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_1_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32106_ clknet_leaf_116_clk _03528_ VGND VGND VPWR VPWR datamem.data_ram\[58\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold358 datamem.data_ram\[49\]\[7\] VGND VGND VPWR VPWR net1508 sky130_fd_sc_hd__dlygate4sd3_1
X_20120_ _05391_ _06586_ _07368_ _07413_ _07120_ VGND VGND VPWR VPWR _07414_ sky130_fd_sc_hd__o32a_1
Xhold369 datamem.data_ram\[7\]\[1\] VGND VGND VPWR VPWR net1519 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_111_3170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30298_ net644 _02033_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[5\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_225_5889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32037_ clknet_leaf_132_clk _03459_ VGND VGND VPWR VPWR datamem.data_ram\[50\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_182_4860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20051_ datamem.data_ram\[37\]\[26\] _06721_ _06668_ datamem.data_ram\[39\]\[26\]
+ _07344_ VGND VGND VPWR VPWR _07345_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_182_4871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1003 rvcpu.dp.rf.reg_file_arr\[13\]\[4\] VGND VGND VPWR VPWR net2153 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1014 rvcpu.dp.rf.reg_file_arr\[1\]\[9\] VGND VGND VPWR VPWR net2164 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1025 rvcpu.dp.rf.reg_file_arr\[3\]\[17\] VGND VGND VPWR VPWR net2175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1036 rvcpu.dp.rf.reg_file_arr\[10\]\[16\] VGND VGND VPWR VPWR net2186 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1047 rvcpu.dp.rf.reg_file_arr\[6\]\[20\] VGND VGND VPWR VPWR net2197 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1058 rvcpu.dp.rf.reg_file_arr\[3\]\[5\] VGND VGND VPWR VPWR net2208 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_159_4306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24790_ _10607_ VGND VGND VPWR VPWR _02472_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_213_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1069 datamem.data_ram\[37\]\[30\] VGND VGND VPWR VPWR net2219 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_4317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20953_ datamem.data_ram\[54\]\[15\] _06625_ _06667_ datamem.data_ram\[55\]\[15\]
+ _06676_ VGND VGND VPWR VPWR _08242_ sky130_fd_sc_hd__o221a_1
XANTENNA_209 _09560_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32939_ clknet_leaf_153_clk _04361_ VGND VGND VPWR VPWR datamem.data_ram\[6\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_178_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26460_ _11535_ rvcpu.ALUResultE\[25\] _11288_ VGND VGND VPWR VPWR _11585_ sky130_fd_sc_hd__a21o_1
XFILLER_0_138_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20884_ datamem.data_ram\[60\]\[14\] datamem.data_ram\[61\]\[14\] _07826_ VGND VGND
+ VPWR VPWR _08174_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_282 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25411_ _10741_ _10960_ _10828_ VGND VGND VPWR VPWR _10961_ sky130_fd_sc_hd__a21oi_4
X_22623_ rvcpu.dp.rf.reg_file_arr\[8\]\[16\] rvcpu.dp.rf.reg_file_arr\[10\]\[16\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[16\] rvcpu.dp.rf.reg_file_arr\[11\]\[16\] _09608_
+ _09532_ VGND VGND VPWR VPWR _09773_ sky130_fd_sc_hd__mux4_1
X_26391_ _11535_ rvcpu.ALUResultE\[5\] VGND VGND VPWR VPWR _11536_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_33_clk clknet_5_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_33_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_192_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28130_ _12435_ net3705 _12528_ VGND VGND VPWR VPWR _12531_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_118_3324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25342_ _10766_ net2143 _10909_ VGND VGND VPWR VPWR _10917_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_118_3335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22554_ rvcpu.dp.rf.reg_file_arr\[20\]\[13\] rvcpu.dp.rf.reg_file_arr\[21\]\[13\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[13\] rvcpu.dp.rf.reg_file_arr\[23\]\[13\] _09401_
+ _09430_ VGND VGND VPWR VPWR _09707_ sky130_fd_sc_hd__mux4_1
XFILLER_0_63_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21505_ rvcpu.dp.rf.reg_file_arr\[16\]\[7\] rvcpu.dp.rf.reg_file_arr\[17\]\[7\] rvcpu.dp.rf.reg_file_arr\[18\]\[7\]
+ rvcpu.dp.rf.reg_file_arr\[19\]\[7\] _08703_ _08721_ VGND VGND VPWR VPWR _08760_
+ sky130_fd_sc_hd__mux4_1
X_28061_ _12494_ VGND VGND VPWR VPWR _03856_ sky130_fd_sc_hd__clkbuf_1
X_25273_ _10724_ net2436 _10878_ VGND VGND VPWR VPWR _10879_ sky130_fd_sc_hd__mux2_1
X_22485_ _09442_ _09635_ _09639_ _09641_ VGND VGND VPWR VPWR _09642_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_133_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27012_ _11889_ net1493 _11885_ _11892_ VGND VGND VPWR VPWR _03409_ sky130_fd_sc_hd__a31o_1
XFILLER_0_17_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24224_ _09244_ net3554 _10279_ VGND VGND VPWR VPWR _10283_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21436_ _08540_ VGND VGND VPWR VPWR _08695_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_79_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_15_Left_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21367_ _08535_ VGND VGND VPWR VPWR _08628_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_130_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20318_ _06916_ _07604_ _07609_ VGND VGND VPWR VPWR _07610_ sky130_fd_sc_hd__and3_1
X_23106_ clknet_1_1__leaf__10087_ VGND VGND VPWR VPWR _10104_ sky130_fd_sc_hd__buf_1
X_28963_ _10047_ _12989_ VGND VGND VPWR VPWR _12990_ sky130_fd_sc_hd__and2_1
X_24086_ _09285_ net2888 _10249_ VGND VGND VPWR VPWR _10255_ sky130_fd_sc_hd__mux2_1
Xhold870 datamem.data_ram\[40\]\[23\] VGND VGND VPWR VPWR net2020 sky130_fd_sc_hd__dlygate4sd3_1
X_21298_ _08559_ VGND VGND VPWR VPWR _08560_ sky130_fd_sc_hd__buf_4
Xhold881 rvcpu.dp.rf.reg_file_arr\[9\]\[7\] VGND VGND VPWR VPWR net2031 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22957__666 clknet_1_0__leaf__10081_ VGND VGND VPWR VPWR net792 sky130_fd_sc_hd__inv_2
X_27914_ _12408_ VGND VGND VPWR VPWR _03795_ sky130_fd_sc_hd__clkbuf_1
Xhold892 rvcpu.dp.rf.reg_file_arr\[0\]\[21\] VGND VGND VPWR VPWR net2042 sky130_fd_sc_hd__dlygate4sd3_1
X_20249_ datamem.data_ram\[37\]\[3\] _06919_ _06954_ datamem.data_ram\[36\]\[3\] VGND
+ VGND VPWR VPWR _07542_ sky130_fd_sc_hd__a22o_1
XFILLER_0_219_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28894_ _12737_ net4278 net68 VGND VGND VPWR VPWR _12952_ sky130_fd_sc_hd__mux2_1
XFILLER_0_229_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_216_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27845_ _12369_ net3010 _12357_ VGND VGND VPWR VPWR _12370_ sky130_fd_sc_hd__mux2_1
Xhold2260 datamem.data_ram\[43\]\[23\] VGND VGND VPWR VPWR net3410 sky130_fd_sc_hd__dlygate4sd3_1
X_14810_ _13303_ _13308_ VGND VGND VPWR VPWR _13363_ sky130_fd_sc_hd__nand2_2
Xhold2271 datamem.data_ram\[6\]\[19\] VGND VGND VPWR VPWR net3421 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2282 rvcpu.dp.rf.reg_file_arr\[19\]\[19\] VGND VGND VPWR VPWR net3432 sky130_fd_sc_hd__dlygate4sd3_1
X_27776_ _12085_ net3812 _12326_ VGND VGND VPWR VPWR _12329_ sky130_fd_sc_hd__mux2_1
Xhold2293 datamem.data_ram\[7\]\[25\] VGND VGND VPWR VPWR net3443 sky130_fd_sc_hd__dlygate4sd3_1
X_15790_ _14179_ net2910 _14221_ VGND VGND VPWR VPWR _14225_ sky130_fd_sc_hd__mux2_1
XFILLER_0_188_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24988_ _10714_ VGND VGND VPWR VPWR _02563_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_24_Left_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29515_ net877 _01250_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[28\]\[22\] sky130_fd_sc_hd__dfxtp_1
Xhold1570 datamem.data_ram\[9\]\[14\] VGND VGND VPWR VPWR net2720 sky130_fd_sc_hd__dlygate4sd3_1
X_14741_ _13293_ VGND VGND VPWR VPWR _13294_ sky130_fd_sc_hd__clkbuf_4
X_26727_ _11719_ VGND VGND VPWR VPWR _03297_ sky130_fd_sc_hd__clkbuf_1
Xhold1581 datamem.data_ram\[34\]\[29\] VGND VGND VPWR VPWR net2731 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1592 datamem.data_ram\[22\]\[15\] VGND VGND VPWR VPWR net2742 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24191__31 clknet_1_0__leaf__10266_ VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__inv_2
XFILLER_0_54_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17460_ _04997_ VGND VGND VPWR VPWR _01311_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_47_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__10227_ clknet_0__10227_ VGND VGND VPWR VPWR clknet_1_1__leaf__10227_
+ sky130_fd_sc_hd__clkbuf_16
X_29446_ net808 _01181_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[30\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_26658_ _11665_ net1834 _11675_ _11678_ VGND VGND VPWR VPWR _03269_ sky130_fd_sc_hd__a31o_1
XFILLER_0_196_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14672_ net2079 _13238_ _13214_ VGND VGND VPWR VPWR _13239_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16411_ _14571_ VGND VGND VPWR VPWR _01834_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_103_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_3_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_3_0_clk sky130_fd_sc_hd__clkbuf_8
X_25609_ _10729_ net3921 net53 VGND VGND VPWR VPWR _11069_ sky130_fd_sc_hd__mux2_1
Xclkbuf_0__10258_ _10258_ VGND VGND VPWR VPWR clknet_0__10258_ sky130_fd_sc_hd__clkbuf_16
X_29377_ clknet_leaf_197_clk _01112_ VGND VGND VPWR VPWR datamem.data_ram\[60\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_17391_ _14172_ net3582 _04960_ VGND VGND VPWR VPWR _04961_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1__f__10158_ clknet_0__10158_ VGND VGND VPWR VPWR clknet_1_1__leaf__10158_
+ sky130_fd_sc_hd__clkbuf_16
X_26589_ _11618_ net1793 _11639_ _11641_ VGND VGND VPWR VPWR _03237_ sky130_fd_sc_hd__a31o_1
XFILLER_0_168_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_24_clk clknet_5_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_24_clk sky130_fd_sc_hd__clkbuf_8
X_19130_ _06448_ VGND VGND VPWR VPWR rvcpu.dp.lAuiPCE\[14\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28328_ _12367_ net3416 _12632_ VGND VGND VPWR VPWR _12638_ sky130_fd_sc_hd__mux2_1
X_16342_ net2182 _14440_ _14525_ VGND VGND VPWR VPWR _14535_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23715__308 clknet_1_0__leaf__10197_ VGND VGND VPWR VPWR net434 sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__10089_ clknet_0__10089_ VGND VGND VPWR VPWR clknet_1_1__leaf__10089_
+ sky130_fd_sc_hd__clkbuf_16
X_19061_ _06386_ _06387_ VGND VGND VPWR VPWR _06388_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_180_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16273_ _14498_ VGND VGND VPWR VPWR _01899_ sky130_fd_sc_hd__clkbuf_1
X_28259_ _12599_ VGND VGND VPWR VPWR _03949_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18012_ rvcpu.dp.plde.RD1E\[2\] _05266_ _05381_ VGND VGND VPWR VPWR _05382_ sky130_fd_sc_hd__a21oi_4
XPHY_EDGE_ROW_33_Left_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15224_ _13298_ _13717_ _13764_ _13315_ VGND VGND VPWR VPWR _13765_ sky130_fd_sc_hd__a211oi_1
X_31270_ clknet_5_0__leaf_clk _02973_ VGND VGND VPWR VPWR rvcpu.dp.plfd.InstrD\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30221_ net575 _01956_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[7\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15155_ _13599_ _13659_ _13696_ _13697_ _13698_ VGND VGND VPWR VPWR _13699_ sky130_fd_sc_hd__o32a_1
XFILLER_0_23_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30152_ net514 _01887_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[0\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_15086_ _13376_ _13383_ _13631_ _13319_ VGND VGND VPWR VPWR _13632_ sky130_fd_sc_hd__o31a_1
X_19963_ datamem.data_ram\[3\]\[18\] _06635_ _06783_ datamem.data_ram\[1\]\[18\] _07256_
+ VGND VGND VPWR VPWR _07257_ sky130_fd_sc_hd__o221a_1
XFILLER_0_10_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23370__1005 clknet_1_0__leaf__10139_ VGND VGND VPWR VPWR net1131 sky130_fd_sc_hd__inv_2
X_18914_ _05537_ _06251_ _06055_ _06253_ VGND VGND VPWR VPWR _06254_ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30083_ net445 _01818_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[11\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_19894_ _06681_ _07186_ _07188_ VGND VGND VPWR VPWR _07189_ sky130_fd_sc_hd__and3_1
XFILLER_0_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18845_ _05889_ _05907_ _06189_ VGND VGND VPWR VPWR _06190_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_220_5764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Left_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_1035 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_220_5775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_220_5786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_588 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18776_ _05315_ _05732_ _05730_ _05316_ VGND VGND VPWR VPWR _06125_ sky130_fd_sc_hd__a2bb2o_1
X_15988_ _14331_ VGND VGND VPWR VPWR _02033_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_222_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_32 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17727_ _05138_ VGND VGND VPWR VPWR _01177_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14939_ _13487_ VGND VGND VPWR VPWR _13488_ sky130_fd_sc_hd__clkbuf_4
X_30985_ clknet_leaf_117_clk _02720_ VGND VGND VPWR VPWR datamem.data_ram\[39\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_222_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23876__437 clknet_1_0__leaf__10221_ VGND VGND VPWR VPWR net563 sky130_fd_sc_hd__inv_2
XFILLER_0_188_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32724_ clknet_leaf_244_clk _04146_ VGND VGND VPWR VPWR datamem.data_ram\[16\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_17658_ net2157 _13237_ _05093_ VGND VGND VPWR VPWR _05102_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_4203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16609_ _14141_ net3685 _04540_ VGND VGND VPWR VPWR _04546_ sky130_fd_sc_hd__mux2_1
XFILLER_0_212_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32655_ clknet_leaf_184_clk _04077_ VGND VGND VPWR VPWR datamem.data_ram\[19\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17589_ _05065_ VGND VGND VPWR VPWR _01242_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_15_clk clknet_5_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_161_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31606_ clknet_leaf_28_clk net1158 VGND VGND VPWR VPWR rvcpu.dp.plmw.PCPlus4W\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_359 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19328_ _06605_ _06623_ VGND VGND VPWR VPWR _06624_ sky130_fd_sc_hd__nand2_4
X_32586_ clknet_leaf_87_clk _04008_ VGND VGND VPWR VPWR datamem.data_ram\[21\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_51_Left_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19259_ rvcpu.dp.plde.ImmExtE\[31\] rvcpu.dp.plde.PCE\[31\] VGND VGND VPWR VPWR _06561_
+ sky130_fd_sc_hd__xnor2_1
X_31537_ clknet_leaf_26_clk net1175 VGND VGND VPWR VPWR rvcpu.dp.plem.PCPlus4M\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_171_4594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22270_ _09433_ _09435_ VGND VGND VPWR VPWR _09436_ sky130_fd_sc_hd__and2_1
X_31468_ clknet_leaf_5_clk rvcpu.dp.SrcBFW_Mux.y\[26\] VGND VGND VPWR VPWR rvcpu.dp.plem.WriteDataM\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_182_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold100 rvcpu.dp.plde.PCPlus4E\[6\] VGND VGND VPWR VPWR net1250 sky130_fd_sc_hd__dlygate4sd3_1
X_21221_ _08487_ _07070_ _08490_ VGND VGND VPWR VPWR _04432_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_103_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_184_4900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30419_ net757 _02154_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[31\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_184_4911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold111 rvcpu.dp.plde.funct3E\[2\] VGND VGND VPWR VPWR net1261 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31399_ clknet_leaf_46_clk _03102_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCE\[16\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_184_4922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold122 rvcpu.dp.plem.ALUResultM\[24\] VGND VGND VPWR VPWR net1272 sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 rvcpu.dp.plde.RdE\[0\] VGND VGND VPWR VPWR net1283 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__10247_ clknet_0__10247_ VGND VGND VPWR VPWR clknet_1_0__leaf__10247_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_229_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold144 datamem.data_ram\[40\]\[7\] VGND VGND VPWR VPWR net1294 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21152_ datamem.data_ram\[21\]\[23\] _06721_ _08439_ _08440_ VGND VGND VPWR VPWR
+ _08441_ sky130_fd_sc_hd__o211a_1
Xhold155 datamem.data_ram\[0\]\[4\] VGND VGND VPWR VPWR net1305 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold166 datamem.data_ram\[46\]\[0\] VGND VGND VPWR VPWR net1316 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold177 datamem.data_ram\[43\]\[3\] VGND VGND VPWR VPWR net1327 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_180_4808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold188 datamem.data_ram\[46\]\[2\] VGND VGND VPWR VPWR net1338 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_180_4819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__10178_ clknet_0__10178_ VGND VGND VPWR VPWR clknet_1_0__leaf__10178_
+ sky130_fd_sc_hd__clkbuf_16
X_20103_ datamem.data_ram\[14\]\[10\] _06717_ _06730_ datamem.data_ram\[11\]\[10\]
+ VGND VGND VPWR VPWR _07397_ sky130_fd_sc_hd__o22a_1
Xhold199 datamem.data_ram\[46\]\[4\] VGND VGND VPWR VPWR net1349 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_186_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21083_ _08370_ _08371_ _07820_ VGND VGND VPWR VPWR _08372_ sky130_fd_sc_hd__o21a_1
X_25960_ net24 _11289_ VGND VGND VPWR VPWR _11303_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20034_ datamem.data_ram\[31\]\[26\] _06761_ _07324_ _07327_ VGND VGND VPWR VPWR
+ _07328_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_60_Left_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24911_ _10673_ VGND VGND VPWR VPWR _02527_ sky130_fd_sc_hd__clkbuf_1
X_25891_ _11142_ VGND VGND VPWR VPWR _11263_ sky130_fd_sc_hd__buf_2
X_23820__403 clknet_1_1__leaf__10207_ VGND VGND VPWR VPWR net529 sky130_fd_sc_hd__inv_2
X_27630_ _12095_ net2010 net80 VGND VGND VPWR VPWR _12250_ sky130_fd_sc_hd__mux2_1
X_24842_ _10448_ net3365 _10631_ VGND VGND VPWR VPWR _10636_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_107_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_198_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27561_ _12213_ VGND VGND VPWR VPWR _03637_ sky130_fd_sc_hd__clkbuf_1
X_24773_ _10596_ VGND VGND VPWR VPWR _02466_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_201_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_178_4759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21985_ _09214_ VGND VGND VPWR VPWR _09215_ sky130_fd_sc_hd__buf_4
XFILLER_0_205_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_248 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29300_ clknet_leaf_1_clk _01035_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD1E\[7\] sky130_fd_sc_hd__dfxtp_1
X_27492_ _12176_ VGND VGND VPWR VPWR _03605_ sky130_fd_sc_hd__clkbuf_1
X_20936_ datamem.data_ram\[54\]\[22\] _06630_ _06665_ datamem.data_ram\[53\]\[22\]
+ _06777_ VGND VGND VPWR VPWR _08226_ sky130_fd_sc_hd__o221a_1
XFILLER_0_7_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0__10112_ _10112_ VGND VGND VPWR VPWR clknet_0__10112_ sky130_fd_sc_hd__clkbuf_16
X_29231_ _13135_ VGND VGND VPWR VPWR _04385_ sky130_fd_sc_hd__clkbuf_1
X_26443_ _11143_ VGND VGND VPWR VPWR _11573_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23655_ clknet_1_1__leaf__10172_ VGND VGND VPWR VPWR _10191_ sky130_fd_sc_hd__buf_1
XFILLER_0_77_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20867_ datamem.data_ram\[39\]\[14\] _07859_ _07862_ datamem.data_ram\[37\]\[14\]
+ _08156_ VGND VGND VPWR VPWR _08157_ sky130_fd_sc_hd__o221a_1
XFILLER_0_83_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29162_ _09243_ net3041 _13094_ VGND VGND VPWR VPWR _13098_ sky130_fd_sc_hd__mux2_1
X_22606_ _09534_ _09756_ VGND VGND VPWR VPWR _09757_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26374_ _11521_ VGND VGND VPWR VPWR _11522_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_42_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20798_ datamem.data_ram\[33\]\[30\] _06949_ _08087_ rvcpu.dp.plem.ALUResultM\[4\]
+ VGND VGND VPWR VPWR _08088_ sky130_fd_sc_hd__a22o_1
XFILLER_0_193_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_3777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28113_ _12361_ net3036 net74 VGND VGND VPWR VPWR _12522_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_666 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25325_ _10907_ VGND VGND VPWR VPWR _02707_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_137_3788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22537_ rvcpu.dp.rf.reg_file_arr\[24\]\[12\] rvcpu.dp.rf.reg_file_arr\[25\]\[12\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[12\] rvcpu.dp.rf.reg_file_arr\[27\]\[12\] _09393_
+ _09465_ VGND VGND VPWR VPWR _09691_ sky130_fd_sc_hd__mux4_1
X_29093_ _13061_ VGND VGND VPWR VPWR _04321_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_146_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28044_ _12485_ VGND VGND VPWR VPWR _03848_ sky130_fd_sc_hd__clkbuf_1
X_25256_ _10538_ net1403 _10867_ _10869_ VGND VGND VPWR VPWR _02676_ sky130_fd_sc_hd__a31o_1
XFILLER_0_162_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22468_ _09622_ _09623_ _09625_ VGND VGND VPWR VPWR _09626_ sky130_fd_sc_hd__a21o_1
XFILLER_0_228_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24207_ _09314_ net3366 _10270_ VGND VGND VPWR VPWR _10274_ sky130_fd_sc_hd__mux2_1
X_21419_ rvcpu.dp.rf.reg_file_arr\[16\]\[3\] rvcpu.dp.rf.reg_file_arr\[17\]\[3\] rvcpu.dp.rf.reg_file_arr\[18\]\[3\]
+ rvcpu.dp.rf.reg_file_arr\[19\]\[3\] _08524_ _08527_ VGND VGND VPWR VPWR _08678_
+ sky130_fd_sc_hd__mux4_1
X_25187_ _10831_ VGND VGND VPWR VPWR _02645_ sky130_fd_sc_hd__clkbuf_1
X_22399_ _09557_ _09559_ _09449_ VGND VGND VPWR VPWR _09560_ sky130_fd_sc_hd__mux2_2
XFILLER_0_20_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29995_ net365 _01730_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[14\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16960_ net3053 _14442_ _04731_ VGND VGND VPWR VPWR _04732_ sky130_fd_sc_hd__mux2_1
XFILLER_0_202_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_1270 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28946_ _12737_ net3948 net67 VGND VGND VPWR VPWR _12980_ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15911_ net2445 _13226_ _14286_ VGND VGND VPWR VPWR _14291_ sky130_fd_sc_hd__mux2_1
X_28877_ _12754_ net2968 _12941_ VGND VGND VPWR VPWR _12943_ sky130_fd_sc_hd__mux2_1
X_16891_ _04683_ VGND VGND VPWR VPWR _04695_ sky130_fd_sc_hd__buf_4
XFILLER_0_216_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_188_Right_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18630_ _05741_ _05375_ _05719_ VGND VGND VPWR VPWR _05987_ sky130_fd_sc_hd__or3_1
XFILLER_0_21_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27828_ _12358_ VGND VGND VPWR VPWR _03759_ sky130_fd_sc_hd__clkbuf_1
X_15842_ net2417 _13229_ _14247_ VGND VGND VPWR VPWR _14253_ sky130_fd_sc_hd__mux2_1
Xhold2090 datamem.data_ram\[23\]\[17\] VGND VGND VPWR VPWR net3240 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18561_ _05675_ _05778_ _05920_ _05776_ VGND VGND VPWR VPWR _05921_ sky130_fd_sc_hd__a211o_1
X_27759_ _12319_ VGND VGND VPWR VPWR _03729_ sky130_fd_sc_hd__clkbuf_1
X_15773_ _14162_ net4260 _14210_ VGND VGND VPWR VPWR _14216_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17512_ _13223_ net2914 _05021_ VGND VGND VPWR VPWR _05025_ sky130_fd_sc_hd__mux2_1
X_14724_ _13277_ VGND VGND VPWR VPWR _13278_ sky130_fd_sc_hd__buf_4
X_18492_ _05850_ _05853_ _05799_ VGND VGND VPWR VPWR _05854_ sky130_fd_sc_hd__mux2_1
X_30770_ clknet_leaf_181_clk _02505_ VGND VGND VPWR VPWR datamem.data_ram\[47\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_540 _06610_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_551 _07177_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_562 _11970_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17443_ _04988_ VGND VGND VPWR VPWR _01319_ sky130_fd_sc_hd__clkbuf_1
X_29429_ net791 _01164_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[30\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_573 _07839_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14655_ _13225_ VGND VGND VPWR VPWR _13226_ sky130_fd_sc_hd__buf_4
XFILLER_0_129_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32440_ clknet_leaf_183_clk _03862_ VGND VGND VPWR VPWR datamem.data_ram\[27\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_931 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17374_ _14156_ net2112 _04949_ VGND VGND VPWR VPWR _04952_ sky130_fd_sc_hd__mux2_1
X_14586_ _13170_ VGND VGND VPWR VPWR _13171_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_188_5000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19113_ _06433_ VGND VGND VPWR VPWR rvcpu.dp.lAuiPCE\[12\] sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_188_5011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16325_ _14526_ VGND VGND VPWR VPWR _01875_ sky130_fd_sc_hd__clkbuf_1
X_32371_ clknet_leaf_241_clk _03793_ VGND VGND VPWR VPWR datamem.data_ram\[2\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19044_ rvcpu.dp.plde.ImmExtE\[4\] rvcpu.dp.plde.PCE\[4\] VGND VGND VPWR VPWR _06373_
+ sky130_fd_sc_hd__and2_1
X_31322_ clknet_leaf_24_clk _03025_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCPlus4E\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16256_ net2582 _14420_ _14489_ VGND VGND VPWR VPWR _14490_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15207_ _13364_ _13353_ _13746_ _13748_ _13646_ VGND VGND VPWR VPWR _13749_ sky130_fd_sc_hd__a32o_1
X_31253_ clknet_leaf_21_clk _02956_ VGND VGND VPWR VPWR rvcpu.dp.plfd.InstrD\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_16187_ _14421_ VGND VGND VPWR VPWR _14443_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_872 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30204_ net558 _01939_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[8\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_15138_ _13304_ VGND VGND VPWR VPWR _13682_ sky130_fd_sc_hd__clkbuf_4
X_31184_ clknet_leaf_37_clk _02887_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCPlus4D\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_227_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_222_5815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30135_ net497 _01870_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[10\]\[26\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_222_5826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15069_ _13397_ _13282_ VGND VGND VPWR VPWR _13615_ sky130_fd_sc_hd__or2_1
X_19946_ datamem.data_ram\[53\]\[18\] _06702_ _06706_ datamem.data_ram\[55\]\[18\]
+ VGND VGND VPWR VPWR _07240_ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_4_clk clknet_5_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_177_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30066_ net428 _01801_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[12\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_19877_ datamem.data_ram\[18\]\[1\] _06931_ _06942_ datamem.data_ram\[19\]\[1\] VGND
+ VGND VPWR VPWR _07172_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_155_Right_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18828_ _06173_ VGND VGND VPWR VPWR _06174_ sky130_fd_sc_hd__inv_2
XFILLER_0_207_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18759_ _05720_ VGND VGND VPWR VPWR _06109_ sky130_fd_sc_hd__buf_2
XFILLER_0_179_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_222_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21770_ _08626_ _09005_ _09007_ _09011_ _08808_ VGND VGND VPWR VPWR _09012_ sky130_fd_sc_hd__a311o_1
X_30968_ clknet_leaf_227_clk _02703_ VGND VGND VPWR VPWR datamem.data_ram\[39\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24170__12 clknet_1_0__leaf__10264_ VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__inv_2
X_20721_ _06583_ _06588_ _07965_ _08011_ VGND VGND VPWR VPWR _08012_ sky130_fd_sc_hd__o31a_1
X_32707_ clknet_leaf_171_clk _04129_ VGND VGND VPWR VPWR datamem.data_ram\[17\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_23125__802 clknet_1_1__leaf__10105_ VGND VGND VPWR VPWR net928 sky130_fd_sc_hd__inv_2
XFILLER_0_37_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_4645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30899_ clknet_leaf_137_clk _02634_ VGND VGND VPWR VPWR datamem.data_ram\[41\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_173_4656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20652_ datamem.data_ram\[38\]\[29\] _06626_ _06812_ datamem.data_ram\[35\]\[29\]
+ VGND VGND VPWR VPWR _07943_ sky130_fd_sc_hd__o22a_1
XFILLER_0_74_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_176_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_175_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32638_ clknet_leaf_283_clk _04060_ VGND VGND VPWR VPWR datamem.data_ram\[1\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20583_ _07824_ VGND VGND VPWR VPWR _07874_ sky130_fd_sc_hd__buf_8
XFILLER_0_184_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32569_ clknet_leaf_252_clk _03991_ VGND VGND VPWR VPWR datamem.data_ram\[22\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_5_18__f_clk clknet_2_2_0_clk VGND VGND VPWR VPWR clknet_5_18__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_2_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25110_ _10786_ VGND VGND VPWR VPWR _02613_ sky130_fd_sc_hd__clkbuf_1
X_22322_ _09482_ _09486_ VGND VGND VPWR VPWR _09487_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_76_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26090_ net1597 _11372_ VGND VGND VPWR VPWR _11380_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_76_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_3652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_3663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22253_ _09418_ VGND VGND VPWR VPWR _09419_ sky130_fd_sc_hd__clkbuf_8
X_25041_ _10474_ net3283 net90 VGND VGND VPWR VPWR _10747_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_3674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21204_ _08471_ _08484_ VGND VGND VPWR VPWR _08485_ sky130_fd_sc_hd__or2_1
X_22184_ _09364_ VGND VGND VPWR VPWR _01109_ sky130_fd_sc_hd__clkbuf_1
X_21135_ datamem.data_ram\[49\]\[23\] _06944_ VGND VGND VPWR VPWR _08424_ sky130_fd_sc_hd__or2_1
X_28800_ _12745_ net4188 _12896_ VGND VGND VPWR VPWR _12902_ sky130_fd_sc_hd__mux2_1
X_29780_ net1126 _01515_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[20\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_26992_ _11880_ VGND VGND VPWR VPWR _03401_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28731_ _12762_ net2789 _12859_ VGND VGND VPWR VPWR _12865_ sky130_fd_sc_hd__mux2_1
X_25943_ net1900 _11290_ _11286_ _11293_ VGND VGND VPWR VPWR _02939_ sky130_fd_sc_hd__o211a_1
X_21066_ _05347_ _06860_ VGND VGND VPWR VPWR _08355_ sky130_fd_sc_hd__nor2_4
XFILLER_0_219_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20017_ datamem.data_ram\[35\]\[2\] _06941_ _06924_ datamem.data_ram\[39\]\[2\] VGND
+ VGND VPWR VPWR _07311_ sky130_fd_sc_hd__a22o_1
X_23212__863 clknet_1_1__leaf__10112_ VGND VGND VPWR VPWR net989 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_122_Right_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28662_ _12828_ VGND VGND VPWR VPWR _04123_ sky130_fd_sc_hd__clkbuf_1
X_25874_ _11251_ VGND VGND VPWR VPWR _02912_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_31_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_213_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27613_ _12157_ net2082 net81 VGND VGND VPWR VPWR _12241_ sky130_fd_sc_hd__mux2_1
XFILLER_0_225_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24825_ _10626_ VGND VGND VPWR VPWR _02488_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_214_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28593_ _12791_ VGND VGND VPWR VPWR _04091_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27544_ _12204_ VGND VGND VPWR VPWR _03629_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_185_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24756_ _10587_ VGND VGND VPWR VPWR _02458_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21968_ rvcpu.dp.rf.reg_file_arr\[16\]\[31\] rvcpu.dp.rf.reg_file_arr\[17\]\[31\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[31\] rvcpu.dp.rf.reg_file_arr\[19\]\[31\] _08548_
+ _08552_ VGND VGND VPWR VPWR _09199_ sky130_fd_sc_hd__mux4_1
XFILLER_0_154_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_3828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20919_ datamem.data_ram\[24\]\[22\] _07191_ _06659_ datamem.data_ram\[25\]\[22\]
+ _08208_ VGND VGND VPWR VPWR _08209_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_139_3839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27475_ _12095_ net2058 _12159_ VGND VGND VPWR VPWR _12167_ sky130_fd_sc_hd__mux2_1
X_24687_ _10550_ VGND VGND VPWR VPWR _02426_ sky130_fd_sc_hd__clkbuf_1
X_21899_ _08626_ _09127_ _09129_ _09133_ _08509_ VGND VGND VPWR VPWR _09134_ sky130_fd_sc_hd__a311o_1
X_29214_ _11533_ net1622 _13122_ _13126_ VGND VGND VPWR VPWR _04377_ sky130_fd_sc_hd__a31o_1
X_26426_ net4453 _11542_ _11561_ _11534_ VGND VGND VPWR VPWR _03154_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_29_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23638_ _10185_ VGND VGND VPWR VPWR _01742_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29145_ _09278_ net3594 net39 VGND VGND VPWR VPWR _13089_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26357_ _11501_ net1741 _11510_ _11512_ VGND VGND VPWR VPWR _03134_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_61_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16110_ _14397_ VGND VGND VPWR VPWR _01969_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25308_ _09300_ _10897_ VGND VGND VPWR VPWR _10898_ sky130_fd_sc_hd__nor2_4
X_29076_ _13052_ VGND VGND VPWR VPWR _04313_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17090_ _14145_ rvcpu.dp.rf.reg_file_arr\[21\]\[24\] _04793_ VGND VGND VPWR VPWR
+ _04801_ sky130_fd_sc_hd__mux2_1
X_26288_ _11476_ VGND VGND VPWR VPWR _03101_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23293__935 clknet_1_0__leaf__10132_ VGND VGND VPWR VPWR net1061 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_21_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28027_ _12435_ net2777 _12473_ VGND VGND VPWR VPWR _12476_ sky130_fd_sc_hd__mux2_1
X_16041_ net1968 _13213_ _14360_ VGND VGND VPWR VPWR _14361_ sky130_fd_sc_hd__mux2_1
X_25239_ _10859_ VGND VGND VPWR VPWR _02669_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_1223 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24124__630 clknet_1_0__leaf__10260_ VGND VGND VPWR VPWR net756 sky130_fd_sc_hd__inv_2
XFILLER_0_209_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19800_ _06753_ _07089_ _07094_ _06713_ VGND VGND VPWR VPWR _07095_ sky130_fd_sc_hd__o31a_1
X_17992_ _05277_ rvcpu.dp.plde.ImmExtE\[4\] VGND VGND VPWR VPWR _05362_ sky130_fd_sc_hd__or2_1
X_29978_ net348 _01713_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[14\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_208_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16943_ net1891 _14426_ _04720_ VGND VGND VPWR VPWR _04723_ sky130_fd_sc_hd__mux2_1
X_19731_ datamem.data_ram\[14\]\[25\] _06683_ _07023_ datamem.data_ram\[10\]\[25\]
+ _07025_ VGND VGND VPWR VPWR _07026_ sky130_fd_sc_hd__o221a_1
X_28929_ _12970_ VGND VGND VPWR VPWR _04248_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_198_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31940_ clknet_leaf_111_clk _03362_ VGND VGND VPWR VPWR datamem.data_ram\[59\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_19662_ _06947_ VGND VGND VPWR VPWR _06958_ sky130_fd_sc_hd__buf_4
X_16874_ _04686_ VGND VGND VPWR VPWR _01602_ sky130_fd_sc_hd__clkbuf_1
X_18613_ _05799_ _05838_ _05970_ VGND VGND VPWR VPWR _05971_ sky130_fd_sc_hd__o21ai_2
X_15825_ net2421 _13204_ _14236_ VGND VGND VPWR VPWR _14244_ sky130_fd_sc_hd__mux2_1
X_31871_ clknet_leaf_125_clk _03325_ VGND VGND VPWR VPWR datamem.data_ram\[56\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19593_ datamem.data_ram\[62\]\[8\] _06743_ _06617_ datamem.data_ram\[60\]\[8\] _06888_
+ VGND VGND VPWR VPWR _06889_ sky130_fd_sc_hd__o221a_1
XFILLER_0_99_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30822_ clknet_leaf_227_clk _02557_ VGND VGND VPWR VPWR datamem.data_ram\[44\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_18544_ _05704_ _05711_ VGND VGND VPWR VPWR _05905_ sky130_fd_sc_hd__nor2_1
X_15756_ _14145_ net4137 _14199_ VGND VGND VPWR VPWR _14207_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14707_ rvcpu.dp.plmw.ALUResultW\[4\] rvcpu.dp.plmw.ReadDataW\[4\] rvcpu.dp.plmw.PCPlus4W\[4\]
+ rvcpu.dp.plmw.lAuiPCW\[4\] _13168_ _13170_ VGND VGND VPWR VPWR _13265_ sky130_fd_sc_hd__mux4_2
XFILLER_0_213_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18475_ _05750_ VGND VGND VPWR VPWR _05837_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30753_ clknet_leaf_179_clk _02488_ VGND VGND VPWR VPWR datamem.data_ram\[48\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_15687_ _13228_ VGND VGND VPWR VPWR _14162_ sky130_fd_sc_hd__buf_4
XFILLER_0_213_1263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_370 rvcpu.dp.plem.ALUResultM\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_381 net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_215_5652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17426_ _04979_ VGND VGND VPWR VPWR _01327_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_392 clknet_1_1__leaf__10079_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_215_5663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14638_ _13212_ VGND VGND VPWR VPWR _13213_ sky130_fd_sc_hd__clkbuf_8
X_30684_ clknet_leaf_85_clk _02419_ VGND VGND VPWR VPWR datamem.data_ram\[4\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32423_ clknet_leaf_74_clk _03845_ VGND VGND VPWR VPWR datamem.data_ram\[28\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17357_ _14139_ net4366 _04938_ VGND VGND VPWR VPWR _04943_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_211_5549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16308_ net3473 _14474_ _14511_ VGND VGND VPWR VPWR _14517_ sky130_fd_sc_hd__mux2_1
X_32354_ clknet_leaf_258_clk _03776_ VGND VGND VPWR VPWR datamem.data_ram\[30\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_17288_ _04906_ VGND VGND VPWR VPWR _01400_ sky130_fd_sc_hd__clkbuf_1
Xclkload301 clknet_1_1__leaf__10204_ VGND VGND VPWR VPWR clkload301/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_153_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload312 clknet_1_0__leaf__10181_ VGND VGND VPWR VPWR clkload312/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload20 clknet_5_24__leaf_clk VGND VGND VPWR VPWR clkload20/Y sky130_fd_sc_hd__inv_8
X_31305_ clknet_leaf_51_clk _03008_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCPlus4E\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_19027_ _06358_ rvcpu.dp.plde.ImmExtE\[1\] _06355_ VGND VGND VPWR VPWR _06359_ sky130_fd_sc_hd__mux2_1
Xclkload323 clknet_1_1__leaf__10153_ VGND VGND VPWR VPWR clkload323/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload31 clknet_leaf_21_clk VGND VGND VPWR VPWR clkload31/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_0_140_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16239_ _13265_ VGND VGND VPWR VPWR _14478_ sky130_fd_sc_hd__buf_4
Xclkload334 clknet_1_1__leaf__10134_ VGND VGND VPWR VPWR clkload334/Y sky130_fd_sc_hd__clkinvlp_4
XPHY_EDGE_ROW_224_Right_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload42 clknet_leaf_30_clk VGND VGND VPWR VPWR clkload42/Y sky130_fd_sc_hd__inv_6
Xclkload345 clknet_1_0__leaf__10112_ VGND VGND VPWR VPWR clkload345/Y sky130_fd_sc_hd__clkinvlp_4
X_32285_ clknet_leaf_242_clk _03707_ VGND VGND VPWR VPWR datamem.data_ram\[33\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload53 clknet_leaf_2_clk VGND VGND VPWR VPWR clkload53/Y sky130_fd_sc_hd__inv_8
Xclkload356 clknet_1_0__leaf__10084_ VGND VGND VPWR VPWR clkload356/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_23_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload64 clknet_leaf_169_clk VGND VGND VPWR VPWR clkload64/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_23_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload75 clknet_leaf_58_clk VGND VGND VPWR VPWR clkload75/X sky130_fd_sc_hd__clkbuf_4
X_31236_ clknet_leaf_31_clk _02939_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCD\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23155__828 clknet_1_0__leaf__10109_ VGND VGND VPWR VPWR net954 sky130_fd_sc_hd__inv_2
Xclkload86 clknet_leaf_50_clk VGND VGND VPWR VPWR clkload86/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload97 clknet_leaf_84_clk VGND VGND VPWR VPWR clkload97/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_80_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_166_4471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31167_ clknet_leaf_9_clk rvcpu.ALUResultE\[26\] VGND VGND VPWR VPWR rvcpu.dp.plem.ALUResultM\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_166_4482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2804 datamem.data_ram\[54\]\[9\] VGND VGND VPWR VPWR net3954 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2815 datamem.data_ram\[60\]\[20\] VGND VGND VPWR VPWR net3965 sky130_fd_sc_hd__dlygate4sd3_1
X_30118_ net480 _01853_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[10\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_19929_ _06753_ _07218_ _07223_ _06713_ VGND VGND VPWR VPWR _07224_ sky130_fd_sc_hd__o31a_1
Xhold2826 rvcpu.dp.rf.reg_file_arr\[19\]\[5\] VGND VGND VPWR VPWR net3976 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2837 rvcpu.dp.rf.reg_file_arr\[18\]\[30\] VGND VGND VPWR VPWR net3987 sky130_fd_sc_hd__dlygate4sd3_1
X_31098_ clknet_leaf_279_clk _02833_ VGND VGND VPWR VPWR datamem.data_ram\[9\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2848 rvcpu.dp.rf.reg_file_arr\[0\]\[23\] VGND VGND VPWR VPWR net3998 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_162_4379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2859 rvcpu.dp.rf.reg_file_arr\[31\]\[20\] VGND VGND VPWR VPWR net4009 sky130_fd_sc_hd__dlygate4sd3_1
X_22940_ rvcpu.dp.plem.WriteDataM\[5\] VGND VGND VPWR VPWR _10069_ sky130_fd_sc_hd__buf_4
XFILLER_0_138_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30049_ net411 _01784_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[12\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_207_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_1300 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_223_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22871_ rvcpu.dp.rf.reg_file_arr\[20\]\[30\] rvcpu.dp.rf.reg_file_arr\[21\]\[30\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[30\] rvcpu.dp.rf.reg_file_arr\[23\]\[30\] _09384_
+ _09577_ VGND VGND VPWR VPWR _10007_ sky130_fd_sc_hd__mux4_1
XFILLER_0_222_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_175_4707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_719 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24610_ _10507_ VGND VGND VPWR VPWR _02392_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21822_ _08515_ _09060_ VGND VGND VPWR VPWR _09061_ sky130_fd_sc_hd__nor2_1
XFILLER_0_223_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25590_ _11057_ net1460 _11053_ _11058_ VGND VGND VPWR VPWR _02821_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_65_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_3397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24541_ _10465_ net3859 net60 VGND VGND VPWR VPWR _10467_ sky130_fd_sc_hd__mux2_1
X_21753_ rvcpu.dp.rf.reg_file_arr\[4\]\[19\] rvcpu.dp.rf.reg_file_arr\[5\]\[19\] rvcpu.dp.rf.reg_file_arr\[6\]\[19\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[19\] _08687_ _08856_ VGND VGND VPWR VPWR _08996_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_59_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20704_ datamem.data_ram\[8\]\[5\] _06937_ _06925_ datamem.data_ram\[15\]\[5\] _06679_
+ VGND VGND VPWR VPWR _07995_ sky130_fd_sc_hd__a221o_1
X_27260_ _10782_ net52 _12042_ net1370 VGND VGND VPWR VPWR _03507_ sky130_fd_sc_hd__a22o_1
XFILLER_0_164_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24472_ _09318_ net3846 _10421_ VGND VGND VPWR VPWR _10426_ sky130_fd_sc_hd__mux2_1
X_21684_ rvcpu.dp.rf.reg_file_arr\[12\]\[15\] rvcpu.dp.rf.reg_file_arr\[13\]\[15\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[15\] rvcpu.dp.rf.reg_file_arr\[15\]\[15\] _08696_
+ _08568_ VGND VGND VPWR VPWR _08931_ sky130_fd_sc_hd__mux4_1
XFILLER_0_65_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_188_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26211_ net1762 _11442_ _03040_ _11443_ VGND VGND VPWR VPWR _03057_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_134_3703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_3714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27191_ _11991_ net1353 _11995_ _12003_ VGND VGND VPWR VPWR _03477_ sky130_fd_sc_hd__a31o_1
XFILLER_0_163_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20635_ datamem.data_ram\[13\]\[29\] _06702_ _06706_ datamem.data_ram\[15\]\[29\]
+ _07925_ VGND VGND VPWR VPWR _07926_ sky130_fd_sc_hd__o221a_1
XFILLER_0_46_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_202_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload3 clknet_5_4__leaf_clk VGND VGND VPWR VPWR clkload3/Y sky130_fd_sc_hd__clkinv_8
XTAP_TAPCELL_ROW_24_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26142_ net1777 _11397_ VGND VGND VPWR VPWR _11407_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_24_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20566_ _06985_ _07807_ _07856_ VGND VGND VPWR VPWR _07857_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_11_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_466 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22305_ rvcpu.dp.rf.reg_file_arr\[0\]\[1\] rvcpu.dp.rf.reg_file_arr\[1\]\[1\] rvcpu.dp.rf.reg_file_arr\[2\]\[1\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[1\] _09463_ _09466_ VGND VGND VPWR VPWR _09470_ sky130_fd_sc_hd__mux4_1
XFILLER_0_225_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26073_ rvcpu.dp.plfd.InstrD\[3\] rvcpu.dp.plfd.InstrD\[2\] rvcpu.dp.plfd.InstrD\[0\]
+ _11366_ VGND VGND VPWR VPWR _11367_ sky130_fd_sc_hd__and4b_1
X_20497_ datamem.data_ram\[38\]\[21\] _06630_ _06688_ datamem.data_ram\[36\]\[21\]
+ VGND VGND VPWR VPWR _07788_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_95_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29901_ clknet_leaf_141_clk _01636_ VGND VGND VPWR VPWR datamem.data_ram\[59\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_25024_ _10736_ VGND VGND VPWR VPWR _02577_ sky130_fd_sc_hd__clkbuf_1
X_22236_ _09401_ VGND VGND VPWR VPWR _09402_ sky130_fd_sc_hd__buf_4
XFILLER_0_30_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29832_ net210 _01567_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[1\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_22167_ _09310_ net3341 _09352_ VGND VGND VPWR VPWR _09355_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23668__265 clknet_1_0__leaf__10193_ VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__inv_2
XFILLER_0_218_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21118_ _06796_ _08394_ _08406_ _06751_ VGND VGND VPWR VPWR _08407_ sky130_fd_sc_hd__o22a_1
X_26975_ _11863_ net1562 _11865_ _11871_ VGND VGND VPWR VPWR _03393_ sky130_fd_sc_hd__a31o_1
X_22098_ _09309_ VGND VGND VPWR VPWR _09310_ sky130_fd_sc_hd__clkbuf_2
X_29763_ net1109 _01498_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[21\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_54_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25926_ net1720 _11279_ VGND VGND VPWR VPWR _11283_ sky130_fd_sc_hd__or2_1
X_28714_ _12698_ net2684 _12850_ VGND VGND VPWR VPWR _12856_ sky130_fd_sc_hd__mux2_1
X_21049_ _07859_ _08332_ _08337_ _06732_ VGND VGND VPWR VPWR _08338_ sky130_fd_sc_hd__o211a_1
XFILLER_0_227_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29694_ net1040 _01429_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[23\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28645_ _12819_ VGND VGND VPWR VPWR _04115_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25857_ _11206_ _11207_ _11237_ VGND VGND VPWR VPWR _11238_ sky130_fd_sc_hd__and3_1
XFILLER_0_202_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15610_ net2415 _13241_ _14103_ VGND VGND VPWR VPWR _14113_ sky130_fd_sc_hd__mux2_1
X_24808_ _10617_ VGND VGND VPWR VPWR _02480_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_213_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28576_ _12782_ VGND VGND VPWR VPWR _04083_ sky130_fd_sc_hd__clkbuf_1
X_16590_ _14191_ net3351 _04525_ VGND VGND VPWR VPWR _04535_ sky130_fd_sc_hd__mux2_1
X_25788_ rvcpu.dp.pcreg.q\[13\] _11178_ VGND VGND VPWR VPWR _11183_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15541_ _13341_ _13510_ _13744_ VGND VGND VPWR VPWR _14067_ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27527_ _12195_ VGND VGND VPWR VPWR _03621_ sky130_fd_sc_hd__clkbuf_1
X_24739_ _10578_ VGND VGND VPWR VPWR _02450_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18260_ rvcpu.dp.plde.RD1E\[23\] _05564_ _05455_ VGND VGND VPWR VPWR _05625_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_194_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15472_ _13572_ _13984_ _13987_ _13993_ _14001_ VGND VGND VPWR VPWR _14002_ sky130_fd_sc_hd__o311a_1
X_27458_ _12157_ net2056 _12143_ VGND VGND VPWR VPWR _12158_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_964 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17211_ _04864_ VGND VGND VPWR VPWR _04865_ sky130_fd_sc_hd__buf_4
X_26409_ _11170_ _11526_ VGND VGND VPWR VPWR _11550_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18191_ _05296_ _05297_ VGND VGND VPWR VPWR _05556_ sky130_fd_sc_hd__and2_1
XFILLER_0_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27389_ _10737_ net3862 net86 VGND VGND VPWR VPWR _12114_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_7_Left_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29128_ _09243_ net3591 _13076_ VGND VGND VPWR VPWR _13080_ sky130_fd_sc_hd__mux2_1
X_17142_ _04538_ _04755_ VGND VGND VPWR VPWR _04828_ sky130_fd_sc_hd__nand2_2
XFILLER_0_80_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23913__470 clknet_1_0__leaf__10225_ VGND VGND VPWR VPWR net596 sky130_fd_sc_hd__inv_2
XFILLER_0_53_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29059_ _13043_ VGND VGND VPWR VPWR _04305_ sky130_fd_sc_hd__clkbuf_1
X_17073_ _04791_ VGND VGND VPWR VPWR _01500_ sky130_fd_sc_hd__clkbuf_1
X_23612__231 clknet_1_0__leaf__10179_ VGND VGND VPWR VPWR net357 sky130_fd_sc_hd__inv_2
XFILLER_0_165_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16024_ net1934 _13187_ _14349_ VGND VGND VPWR VPWR _14352_ sky130_fd_sc_hd__mux2_1
X_32070_ clknet_leaf_121_clk _03492_ VGND VGND VPWR VPWR datamem.data_ram\[29\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_23219__869 clknet_1_0__leaf__10124_ VGND VGND VPWR VPWR net995 sky130_fd_sc_hd__inv_2
XFILLER_0_21_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31021_ clknet_leaf_59_clk _02756_ VGND VGND VPWR VPWR datamem.data_ram\[40\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17975_ _05344_ _05345_ VGND VGND VPWR VPWR _05346_ sky130_fd_sc_hd__nor2_2
XFILLER_0_218_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19714_ datamem.data_ram\[31\]\[0\] _06925_ _06958_ datamem.data_ram\[25\]\[0\] VGND
+ VGND VPWR VPWR _07010_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_204_5386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16926_ _04713_ VGND VGND VPWR VPWR _01577_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_204_5397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32972_ clknet_leaf_143_clk _04394_ VGND VGND VPWR VPWR datamem.data_ram\[63\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19645_ _06605_ _06940_ VGND VGND VPWR VPWR _06941_ sky130_fd_sc_hd__nor2_8
X_31923_ _04435_ net118 VGND VGND VPWR VPWR datamem.rd_data_mem\[28\] sky130_fd_sc_hd__dlxtn_1
XFILLER_0_204_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16857_ net1992 _14476_ _04670_ VGND VGND VPWR VPWR _04677_ sky130_fd_sc_hd__mux2_1
XFILLER_0_189_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_220_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_217_5703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_196_5198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15808_ _13174_ rvcpu.dp.plmw.RdW\[3\] _13176_ VGND VGND VPWR VPWR _14234_ sky130_fd_sc_hd__or3_4
XTAP_TAPCELL_ROW_217_5714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31854_ clknet_leaf_90_clk _03308_ VGND VGND VPWR VPWR datamem.data_ram\[61\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_16788_ _04640_ VGND VGND VPWR VPWR _01650_ sky130_fd_sc_hd__clkbuf_1
X_19576_ datamem.data_ram\[11\]\[8\] _06731_ _06726_ datamem.data_ram\[15\]\[8\] _06741_
+ VGND VGND VPWR VPWR _06872_ sky130_fd_sc_hd__o221a_1
XFILLER_0_220_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18527_ _05378_ _05400_ _05887_ VGND VGND VPWR VPWR _05888_ sky130_fd_sc_hd__o21a_1
X_30805_ clknet_leaf_154_clk _02540_ VGND VGND VPWR VPWR datamem.data_ram\[45\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15739_ rvcpu.dp.plmw.RegWriteW rvcpu.dp.plmw.RdW\[0\] rvcpu.dp.plmw.RdW\[1\] VGND
+ VGND VPWR VPWR _14197_ sky130_fd_sc_hd__and3_4
X_31785_ clknet_leaf_53_clk _03239_ VGND VGND VPWR VPWR datamem.data_ram\[8\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_213_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18458_ _05370_ _05674_ _05820_ VGND VGND VPWR VPWR _05821_ sky130_fd_sc_hd__and3_1
X_30736_ clknet_leaf_224_clk _02471_ VGND VGND VPWR VPWR datamem.data_ram\[47\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17409_ _14191_ net3794 _04960_ VGND VGND VPWR VPWR _04970_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30667_ clknet_leaf_139_clk _02402_ VGND VGND VPWR VPWR datamem.data_ram\[50\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18389_ _05752_ VGND VGND VPWR VPWR _05753_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20420_ datamem.data_ram\[50\]\[12\] _06691_ _07708_ _07711_ VGND VGND VPWR VPWR
+ _07712_ sky130_fd_sc_hd__o211a_1
X_32406_ clknet_leaf_250_clk _03828_ VGND VGND VPWR VPWR datamem.data_ram\[29\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30598_ clknet_leaf_217_clk _02333_ VGND VGND VPWR VPWR datamem.data_ram\[53\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload120 clknet_leaf_105_clk VGND VGND VPWR VPWR clkload120/Y sky130_fd_sc_hd__clkinvlp_4
X_20351_ datamem.data_ram\[53\]\[4\] _06970_ _07639_ _07642_ VGND VGND VPWR VPWR _07643_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_31_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_168_4522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32337_ clknet_leaf_231_clk _03759_ VGND VGND VPWR VPWR datamem.data_ram\[30\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload131 clknet_leaf_262_clk VGND VGND VPWR VPWR clkload131/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_168_4533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload142 clknet_leaf_247_clk VGND VGND VPWR VPWR clkload142/Y sky130_fd_sc_hd__clkinv_4
Xclkload153 clknet_leaf_276_clk VGND VGND VPWR VPWR clkload153/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload164 clknet_leaf_265_clk VGND VGND VPWR VPWR clkload164/Y sky130_fd_sc_hd__inv_6
X_23070_ _09279_ datamem.data_ram\[5\]\[11\] _10093_ VGND VGND VPWR VPWR _10097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20282_ datamem.data_ram\[29\]\[19\] _06865_ _06672_ datamem.data_ram\[31\]\[19\]
+ VGND VGND VPWR VPWR _07575_ sky130_fd_sc_hd__o22a_1
Xclkload175 clknet_leaf_230_clk VGND VGND VPWR VPWR clkload175/Y sky130_fd_sc_hd__clkinv_4
X_32268_ clknet_leaf_225_clk _03690_ VGND VGND VPWR VPWR datamem.data_ram\[33\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_222_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload186 clknet_leaf_220_clk VGND VGND VPWR VPWR clkload186/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_87_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22021_ rvcpu.dp.plem.WriteDataM\[4\] _09215_ _09219_ _09246_ VGND VGND VPWR VPWR
+ _09247_ sky130_fd_sc_hd__a31o_4
XFILLER_0_11_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload197 clknet_leaf_187_clk VGND VGND VPWR VPWR clkload197/Y sky130_fd_sc_hd__inv_6
X_31219_ clknet_leaf_37_clk _02922_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCD\[8\] sky130_fd_sc_hd__dfxtp_1
Xhold3302 rvcpu.dp.pcreg.q\[29\] VGND VGND VPWR VPWR net4452 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32199_ clknet_leaf_193_clk _03621_ VGND VGND VPWR VPWR datamem.data_ram\[36\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2601 datamem.data_ram\[60\]\[22\] VGND VGND VPWR VPWR net3751 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2612 rvcpu.dp.rf.reg_file_arr\[13\]\[29\] VGND VGND VPWR VPWR net3762 sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 rvcpu.dp.plem.lAuiPCM\[20\] VGND VGND VPWR VPWR net1165 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2623 datamem.data_ram\[57\]\[15\] VGND VGND VPWR VPWR net3773 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 rvcpu.dp.plfd.InstrD\[28\] VGND VGND VPWR VPWR net1176 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_127_3540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2634 datamem.data_ram\[33\]\[27\] VGND VGND VPWR VPWR net3784 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 rvcpu.dp.plem.PCPlus4M\[6\] VGND VGND VPWR VPWR net1187 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_127_3551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1900 datamem.data_ram\[41\]\[25\] VGND VGND VPWR VPWR net3050 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2645 datamem.data_ram\[45\]\[28\] VGND VGND VPWR VPWR net3795 sky130_fd_sc_hd__dlygate4sd3_1
X_26760_ _11679_ _11738_ VGND VGND VPWR VPWR _11740_ sky130_fd_sc_hd__and2_1
Xhold1911 datamem.data_ram\[27\]\[29\] VGND VGND VPWR VPWR net3061 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2656 datamem.data_ram\[50\]\[27\] VGND VGND VPWR VPWR net3806 sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 rvcpu.dp.plem.lAuiPCM\[1\] VGND VGND VPWR VPWR net1198 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2667 datamem.data_ram\[29\]\[16\] VGND VGND VPWR VPWR net3817 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1922 datamem.data_ram\[18\]\[29\] VGND VGND VPWR VPWR net3072 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold59 rvcpu.dp.plem.lAuiPCM\[14\] VGND VGND VPWR VPWR net1209 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1933 datamem.data_ram\[53\]\[17\] VGND VGND VPWR VPWR net3083 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2678 datamem.data_ram\[9\]\[24\] VGND VGND VPWR VPWR net3828 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_67_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1944 datamem.data_ram\[32\]\[28\] VGND VGND VPWR VPWR net3094 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2689 datamem.data_ram\[44\]\[24\] VGND VGND VPWR VPWR net3839 sky130_fd_sc_hd__dlygate4sd3_1
X_25711_ _10820_ net2495 _11124_ VGND VGND VPWR VPWR _11129_ sky130_fd_sc_hd__mux2_1
XFILLER_0_194_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22923_ _10055_ VGND VGND VPWR VPWR _10056_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_123_3437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1955 rvcpu.dp.rf.reg_file_arr\[26\]\[8\] VGND VGND VPWR VPWR net3105 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__10260_ clknet_0__10260_ VGND VGND VPWR VPWR clknet_1_1__leaf__10260_
+ sky130_fd_sc_hd__clkbuf_16
X_26691_ _11683_ net1839 _11693_ _11699_ VGND VGND VPWR VPWR _03281_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_123_3448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1966 datamem.data_ram\[44\]\[30\] VGND VGND VPWR VPWR net3116 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1977 datamem.data_ram\[23\]\[22\] VGND VGND VPWR VPWR net3127 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_123_3459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1988 datamem.data_ram\[61\]\[29\] VGND VGND VPWR VPWR net3138 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28430_ _09313_ VGND VGND VPWR VPWR _12694_ sky130_fd_sc_hd__clkbuf_2
X_25642_ _11085_ net1781 _11077_ _11090_ VGND VGND VPWR VPWR _02841_ sky130_fd_sc_hd__a31o_1
Xhold1999 datamem.data_ram\[51\]\[13\] VGND VGND VPWR VPWR net3149 sky130_fd_sc_hd__dlygate4sd3_1
X_22854_ rvcpu.dp.rf.reg_file_arr\[28\]\[29\] rvcpu.dp.rf.reg_file_arr\[30\]\[29\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[29\] rvcpu.dp.rf.reg_file_arr\[31\]\[29\] _09381_
+ _09423_ VGND VGND VPWR VPWR _09991_ sky130_fd_sc_hd__mux4_1
Xclkbuf_1_1__f__10191_ clknet_0__10191_ VGND VGND VPWR VPWR clknet_1_1__leaf__10191_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_78_330 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28361_ _12655_ VGND VGND VPWR VPWR _03995_ sky130_fd_sc_hd__clkbuf_1
X_21805_ _08742_ _09044_ VGND VGND VPWR VPWR _09045_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25573_ _10066_ VGND VGND VPWR VPWR _11047_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_196_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22785_ _09442_ _09921_ _09923_ _09925_ VGND VGND VPWR VPWR _09926_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_213_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27312_ _11946_ _12066_ VGND VGND VPWR VPWR _12071_ sky130_fd_sc_hd__and2_1
XFILLER_0_210_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23324__964 clknet_1_0__leaf__10134_ VGND VGND VPWR VPWR net1090 sky130_fd_sc_hd__inv_2
X_24524_ _10457_ VGND VGND VPWR VPWR _02356_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28292_ _12618_ VGND VGND VPWR VPWR _03963_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_26_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21736_ _08835_ _08979_ VGND VGND VPWR VPWR _08980_ sky130_fd_sc_hd__or2_1
XFILLER_0_164_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27243_ _11972_ _12031_ VGND VGND VPWR VPWR _12035_ sky130_fd_sc_hd__and2_1
XFILLER_0_148_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24455_ _10069_ VGND VGND VPWR VPWR _10416_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_97_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21667_ _08817_ _08912_ _08914_ _08700_ VGND VGND VPWR VPWR _08915_ sky130_fd_sc_hd__a211o_1
X_23023__725 clknet_1_0__leaf__10088_ VGND VGND VPWR VPWR net851 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_97_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27174_ _11991_ net1508 _11983_ _11993_ VGND VGND VPWR VPWR _03470_ sky130_fd_sc_hd__a31o_1
X_20618_ _07906_ _07908_ VGND VGND VPWR VPWR _07909_ sky130_fd_sc_hd__and2_1
X_24386_ _09248_ net3361 _10367_ VGND VGND VPWR VPWR _10372_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21598_ _08798_ _08848_ VGND VGND VPWR VPWR _08849_ sky130_fd_sc_hd__or2_1
XFILLER_0_163_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26125_ _11398_ VGND VGND VPWR VPWR _03015_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_286_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_286_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_149_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23103__782 clknet_1_1__leaf__10103_ VGND VGND VPWR VPWR net908 sky130_fd_sc_hd__inv_2
X_20549_ _07839_ VGND VGND VPWR VPWR _07840_ sky130_fd_sc_hd__buf_6
XFILLER_0_120_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26056_ _11047_ _11351_ VGND VGND VPWR VPWR _11357_ sky130_fd_sc_hd__and2_1
XFILLER_0_104_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25007_ _10542_ _10640_ _10705_ VGND VGND VPWR VPWR _10725_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_56_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22219_ _09384_ VGND VGND VPWR VPWR _09385_ sky130_fd_sc_hd__buf_8
X_23199_ _10120_ VGND VGND VPWR VPWR _01368_ sky130_fd_sc_hd__clkbuf_1
X_29815_ net193 _01550_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[1\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_14972_ rvcpu.dp.pcreg.q\[9\] VGND VGND VPWR VPWR _13521_ sky130_fd_sc_hd__clkbuf_4
X_17760_ rvcpu.dp.plde.Rs2E\[3\] _05157_ VGND VGND VPWR VPWR _05158_ sky130_fd_sc_hd__nor2_1
X_29746_ net1092 _01481_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[21\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_26958_ _11835_ _11854_ VGND VGND VPWR VPWR _11861_ sky130_fd_sc_hd__and2_1
X_16711_ _14175_ net3417 _04598_ VGND VGND VPWR VPWR _04600_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25909_ _11146_ VGND VGND VPWR VPWR _11273_ sky130_fd_sc_hd__buf_2
X_17691_ _13184_ net3900 _05118_ VGND VGND VPWR VPWR _05120_ sky130_fd_sc_hd__mux2_1
X_26889_ _11687_ _11810_ VGND VGND VPWR VPWR _11817_ sky130_fd_sc_hd__and2_1
X_29677_ net1023 _01412_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[23\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_214_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_210_clk clknet_5_22__leaf_clk VGND VGND VPWR VPWR clknet_leaf_210_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_159_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19430_ _06725_ VGND VGND VPWR VPWR _06726_ sky130_fd_sc_hd__buf_6
X_16642_ _04563_ VGND VGND VPWR VPWR _01719_ sky130_fd_sc_hd__clkbuf_1
X_28628_ _12810_ VGND VGND VPWR VPWR _04107_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_202_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19361_ _06656_ VGND VGND VPWR VPWR _06657_ sky130_fd_sc_hd__buf_6
X_16573_ _04526_ VGND VGND VPWR VPWR _01759_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28559_ _12773_ VGND VGND VPWR VPWR _04075_ sky130_fd_sc_hd__clkbuf_1
X_26501__54 clknet_1_0__leaf__11601_ VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__inv_2
XFILLER_0_123_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_694 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15524_ _13514_ _13796_ _14046_ _14047_ _14050_ VGND VGND VPWR VPWR _14051_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_191_5073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18312_ _05676_ VGND VGND VPWR VPWR _05677_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_191_5084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31570_ clknet_leaf_71_clk datamem.rd_data_mem\[20\] VGND VGND VPWR VPWR rvcpu.dp.plmw.ReadDataW\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_19292_ _06587_ rvcpu.dp.plem.ALUResultM\[0\] VGND VGND VPWR VPWR _06588_ sky130_fd_sc_hd__nand2_2
XFILLER_0_167_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18243_ net103 _05409_ _05410_ _05607_ VGND VGND VPWR VPWR _05608_ sky130_fd_sc_hd__o22a_1
XFILLER_0_132_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30521_ clknet_leaf_197_clk _02256_ VGND VGND VPWR VPWR datamem.data_ram\[56\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_23299__941 clknet_1_1__leaf__10132_ VGND VGND VPWR VPWR net1067 sky130_fd_sc_hd__inv_2
X_15455_ _13402_ _13505_ _13294_ _13292_ VGND VGND VPWR VPWR _13985_ sky130_fd_sc_hd__a211o_1
XFILLER_0_182_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23456__105 clknet_1_0__leaf__10157_ VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__inv_2
XFILLER_0_167_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18174_ rvcpu.dp.plde.RD1E\[27\] _05291_ _05538_ VGND VGND VPWR VPWR _05539_ sky130_fd_sc_hd__o21a_1
X_30452_ net790 _02187_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[29\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_15386_ _13706_ _13339_ _13918_ _13439_ VGND VGND VPWR VPWR _13919_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_5_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17125_ _04819_ VGND VGND VPWR VPWR _01476_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_338 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_277_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_277_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_13_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_4091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30383_ clknet_leaf_266_clk _02118_ VGND VGND VPWR VPWR datamem.data_ram\[58\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold507 rvcpu.dp.pcreg.q\[11\] VGND VGND VPWR VPWR net1657 sky130_fd_sc_hd__dlygate4sd3_1
Xhold518 rvcpu.dp.pcreg.q\[22\] VGND VGND VPWR VPWR net1668 sky130_fd_sc_hd__dlygate4sd3_1
X_32122_ clknet_leaf_214_clk _03544_ VGND VGND VPWR VPWR datamem.data_ram\[7\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold529 rvcpu.dp.pcreg.q\[0\] VGND VGND VPWR VPWR net1679 sky130_fd_sc_hd__dlygate4sd3_1
X_17056_ net2769 _14470_ _04779_ VGND VGND VPWR VPWR _04783_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_650 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16007_ _14341_ VGND VGND VPWR VPWR _02024_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32053_ clknet_leaf_127_clk _03475_ VGND VGND VPWR VPWR datamem.data_ram\[30\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_206_5437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_206_5448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31004_ clknet_leaf_100_clk _02739_ VGND VGND VPWR VPWR datamem.data_ram\[22\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_198_5238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1207 datamem.data_ram\[30\]\[15\] VGND VGND VPWR VPWR net2357 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_198_5249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17958_ _05329_ VGND VGND VPWR VPWR rvcpu.dp.SrcBFW_Mux.y\[12\] sky130_fd_sc_hd__buf_1
Xhold1218 datamem.data_ram\[63\]\[29\] VGND VGND VPWR VPWR net2368 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1229 rvcpu.dp.rf.reg_file_arr\[6\]\[0\] VGND VGND VPWR VPWR net2379 sky130_fd_sc_hd__dlygate4sd3_1
X_16909_ _04704_ VGND VGND VPWR VPWR _01585_ sky130_fd_sc_hd__clkbuf_1
X_32955_ clknet_leaf_97_clk _04377_ VGND VGND VPWR VPWR datamem.data_ram\[6\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17889_ rvcpu.dp.plde.Rs1E\[3\] _05242_ _05259_ _05260_ _05261_ VGND VGND VPWR VPWR
+ _05262_ sky130_fd_sc_hd__o2111a_1
X_23805__389 clknet_1_1__leaf__10206_ VGND VGND VPWR VPWR net515 sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_201_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_201_clk
+ sky130_fd_sc_hd__clkbuf_8
X_19628_ _06923_ VGND VGND VPWR VPWR _06924_ sky130_fd_sc_hd__buf_4
X_31906_ _04417_ net120 VGND VGND VPWR VPWR datamem.rd_data_mem\[11\] sky130_fd_sc_hd__dlxtn_1
XFILLER_0_73_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32886_ clknet_leaf_283_clk _04308_ VGND VGND VPWR VPWR datamem.data_ram\[10\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_195 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19559_ datamem.data_ram\[0\]\[24\] _06811_ _06669_ datamem.data_ram\[7\]\[24\] VGND
+ VGND VPWR VPWR _06855_ sky130_fd_sc_hd__o22a_1
X_31837_ clknet_leaf_209_clk _03291_ VGND VGND VPWR VPWR datamem.data_ram\[3\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_157_4256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_157_4267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22570_ _09534_ _09722_ VGND VGND VPWR VPWR _09723_ sky130_fd_sc_hd__and2_1
XFILLER_0_119_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31768_ clknet_leaf_213_clk _03222_ VGND VGND VPWR VPWR datamem.data_ram\[1\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_622 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21521_ _08565_ _08773_ _08775_ _08652_ VGND VGND VPWR VPWR _08776_ sky130_fd_sc_hd__o211a_1
XFILLER_0_146_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23619__237 clknet_1_0__leaf__10180_ VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__inv_2
X_30719_ clknet_leaf_179_clk _02454_ VGND VGND VPWR VPWR datamem.data_ram\[49\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31699_ clknet_leaf_46_clk _03157_ VGND VGND VPWR VPWR rvcpu.dp.pcreg.q\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24240_ _10291_ VGND VGND VPWR VPWR _02238_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_161_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21452_ _08515_ _08709_ _08513_ VGND VGND VPWR VPWR _08710_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_8_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_268_clk clknet_5_19__leaf_clk VGND VGND VPWR VPWR clknet_leaf_268_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_181_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_3274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20403_ datamem.data_ram\[38\]\[12\] _07085_ _06618_ datamem.data_ram\[36\]\[12\]
+ VGND VGND VPWR VPWR _07695_ sky130_fd_sc_hd__o22a_1
XFILLER_0_71_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_3285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21383_ rvcpu.dp.rf.reg_file_arr\[4\]\[1\] rvcpu.dp.rf.reg_file_arr\[5\]\[1\] rvcpu.dp.rf.reg_file_arr\[6\]\[1\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[1\] _08551_ _08555_ VGND VGND VPWR VPWR _08644_ sky130_fd_sc_hd__mux4_1
XFILLER_0_4_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20334_ datamem.data_ram\[37\]\[4\] _06921_ _06993_ datamem.data_ram\[39\]\[4\] VGND
+ VGND VPWR VPWR _07626_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_187_4975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_187_4986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput16 net16 VGND VGND VPWR VPWR Instr[22] sky130_fd_sc_hd__buf_2
Xoutput27 net27 VGND VGND VPWR VPWR Instr[3] sky130_fd_sc_hd__buf_2
XFILLER_0_3_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20265_ datamem.data_ram\[56\]\[19\] _06697_ _06657_ datamem.data_ram\[57\]\[19\]
+ _07557_ VGND VGND VPWR VPWR _07558_ sky130_fd_sc_hd__o221a_1
X_27930_ _12134_ net4415 _12412_ VGND VGND VPWR VPWR _12417_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_129_3602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_79_Left_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold3110 rvcpu.dp.rf.reg_file_arr\[31\]\[16\] VGND VGND VPWR VPWR net4260 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3121 datamem.data_ram\[27\]\[27\] VGND VGND VPWR VPWR net4271 sky130_fd_sc_hd__dlygate4sd3_1
X_22004_ _09233_ VGND VGND VPWR VPWR _01060_ sky130_fd_sc_hd__clkbuf_1
X_27861_ _12136_ net3525 _12373_ VGND VGND VPWR VPWR _12379_ sky130_fd_sc_hd__mux2_1
Xhold3132 rvcpu.dp.rf.reg_file_arr\[5\]\[7\] VGND VGND VPWR VPWR net4282 sky130_fd_sc_hd__dlygate4sd3_1
X_20196_ datamem.data_ram\[39\]\[11\] _06760_ _06699_ datamem.data_ram\[33\]\[11\]
+ VGND VGND VPWR VPWR _07489_ sky130_fd_sc_hd__o22a_1
Xhold3143 datamem.data_ram\[55\]\[8\] VGND VGND VPWR VPWR net4293 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3154 datamem.data_ram\[14\]\[31\] VGND VGND VPWR VPWR net4304 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3165 rvcpu.dp.rf.reg_file_arr\[28\]\[30\] VGND VGND VPWR VPWR net4315 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2420 rvcpu.dp.rf.reg_file_arr\[28\]\[0\] VGND VGND VPWR VPWR net3570 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29600_ net954 _01335_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[25\]\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_51_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2431 datamem.data_ram\[23\]\[9\] VGND VGND VPWR VPWR net3581 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3176 rvcpu.dp.rf.reg_file_arr\[0\]\[11\] VGND VGND VPWR VPWR net4326 sky130_fd_sc_hd__dlygate4sd3_1
X_26812_ _11767_ net1440 _11761_ _11770_ VGND VGND VPWR VPWR _03331_ sky130_fd_sc_hd__a31o_1
X_27792_ _12128_ net3232 _12336_ VGND VGND VPWR VPWR _12338_ sky130_fd_sc_hd__mux2_1
Xhold2442 datamem.data_ram\[35\]\[19\] VGND VGND VPWR VPWR net3592 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3187 datamem.data_ram\[59\]\[18\] VGND VGND VPWR VPWR net4337 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3198 rvcpu.dp.rf.reg_file_arr\[21\]\[4\] VGND VGND VPWR VPWR net4348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2453 datamem.data_ram\[22\]\[13\] VGND VGND VPWR VPWR net3603 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_3993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2464 datamem.data_ram\[63\]\[23\] VGND VGND VPWR VPWR net3614 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1730 datamem.data_ram\[21\]\[24\] VGND VGND VPWR VPWR net2880 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2475 datamem.data_ram\[63\]\[11\] VGND VGND VPWR VPWR net3625 sky130_fd_sc_hd__dlygate4sd3_1
X_26743_ _11700_ net1753 _11724_ _11729_ VGND VGND VPWR VPWR _03303_ sky130_fd_sc_hd__a31o_1
Xhold1741 datamem.data_ram\[17\]\[17\] VGND VGND VPWR VPWR net2891 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2486 datamem.data_ram\[22\]\[18\] VGND VGND VPWR VPWR net3636 sky130_fd_sc_hd__dlygate4sd3_1
X_29531_ clknet_leaf_174_clk _01266_ VGND VGND VPWR VPWR datamem.data_ram\[5\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_23955_ _10231_ VGND VGND VPWR VPWR _02013_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1752 datamem.data_ram\[3\]\[13\] VGND VGND VPWR VPWR net2902 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2497 datamem.data_ram\[46\]\[17\] VGND VGND VPWR VPWR net3647 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1763 rvcpu.dp.rf.reg_file_arr\[11\]\[13\] VGND VGND VPWR VPWR net2913 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1774 datamem.data_ram\[6\]\[12\] VGND VGND VPWR VPWR net2924 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22906_ _10040_ VGND VGND VPWR VPWR _01155_ sky130_fd_sc_hd__clkbuf_1
X_29462_ net824 _01197_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[2\]\[1\] sky130_fd_sc_hd__dfxtp_1
Xhold1785 datamem.data_ram\[49\]\[12\] VGND VGND VPWR VPWR net2935 sky130_fd_sc_hd__dlygate4sd3_1
X_26674_ _10072_ VGND VGND VPWR VPWR _11689_ sky130_fd_sc_hd__buf_2
XFILLER_0_212_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1796 datamem.data_ram\[61\]\[24\] VGND VGND VPWR VPWR net2946 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f__10243_ clknet_0__10243_ VGND VGND VPWR VPWR clknet_1_1__leaf__10243_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_169_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25625_ _10946_ _11075_ VGND VGND VPWR VPWR _11079_ sky130_fd_sc_hd__nor2_2
XFILLER_0_212_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28413_ _12683_ VGND VGND VPWR VPWR _04019_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_88_Left_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_211_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29393_ clknet_leaf_2_clk _01128_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD2E\[4\] sky130_fd_sc_hd__dfxtp_1
X_23248__895 clknet_1_1__leaf__10127_ VGND VGND VPWR VPWR net1021 sky130_fd_sc_hd__inv_2
X_22837_ rvcpu.dp.rf.reg_file_arr\[28\]\[28\] rvcpu.dp.rf.reg_file_arr\[30\]\[28\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[28\] rvcpu.dp.rf.reg_file_arr\[31\]\[28\] _09382_
+ _09417_ VGND VGND VPWR VPWR _09975_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_49_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__10174_ clknet_0__10174_ VGND VGND VPWR VPWR clknet_1_1__leaf__10174_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_156_508 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28344_ _12646_ VGND VGND VPWR VPWR _03987_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25556_ _11036_ VGND VGND VPWR VPWR _02809_ sky130_fd_sc_hd__clkbuf_1
X_22768_ rvcpu.dp.rf.reg_file_arr\[0\]\[24\] rvcpu.dp.rf.reg_file_arr\[1\]\[24\] rvcpu.dp.rf.reg_file_arr\[2\]\[24\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[24\] _09714_ _09383_ VGND VGND VPWR VPWR _09910_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_67_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24507_ _09243_ VGND VGND VPWR VPWR _10446_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_45_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28275_ _12367_ net3394 _12603_ VGND VGND VPWR VPWR _12609_ sky130_fd_sc_hd__mux2_1
X_21719_ _08663_ _08961_ _08963_ _08575_ VGND VGND VPWR VPWR _08964_ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25487_ _08151_ net110 VGND VGND VPWR VPWR _10997_ sky130_fd_sc_hd__nor2_8
X_22699_ rvcpu.dp.rf.reg_file_arr\[8\]\[20\] rvcpu.dp.rf.reg_file_arr\[10\]\[20\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[20\] rvcpu.dp.rf.reg_file_arr\[11\]\[20\] _09608_
+ _09656_ VGND VGND VPWR VPWR _09845_ sky130_fd_sc_hd__mux4_1
XFILLER_0_82_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15240_ _13305_ _13346_ VGND VGND VPWR VPWR _13780_ sky130_fd_sc_hd__nand2_4
X_27226_ _11946_ _12019_ VGND VGND VPWR VPWR _12025_ sky130_fd_sc_hd__and2_1
XFILLER_0_192_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24438_ _10403_ VGND VGND VPWR VPWR _10404_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_191_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_259_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_259_clk
+ sky130_fd_sc_hd__clkbuf_8
X_15171_ _13307_ _13317_ _13707_ VGND VGND VPWR VPWR _13714_ sky130_fd_sc_hd__a21o_1
X_27157_ _10268_ _08059_ _11898_ VGND VGND VPWR VPWR _11984_ sky130_fd_sc_hd__and3_1
X_24369_ _10362_ VGND VGND VPWR VPWR _02296_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26108_ _11389_ VGND VGND VPWR VPWR _03007_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_205_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_97_Left_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27088_ _10402_ _11075_ VGND VGND VPWR VPWR _11939_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26039_ _11121_ net1528 _11339_ _11346_ VGND VGND VPWR VPWR _02982_ sky130_fd_sc_hd__a31o_1
X_18930_ _05551_ _05730_ _06108_ _05529_ _06259_ VGND VGND VPWR VPWR _06269_ sky130_fd_sc_hd__a221o_1
XFILLER_0_31_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_219_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18861_ _05693_ _05917_ _05866_ VGND VGND VPWR VPWR _06205_ sky130_fd_sc_hd__o21a_1
XFILLER_0_120_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_201_5312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17812_ _05202_ VGND VGND VPWR VPWR rvcpu.dp.SrcBFW_Mux.y\[29\] sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_24_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_219_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_201_5323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18792_ _06137_ _06139_ VGND VGND VPWR VPWR _06140_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_175_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14955_ _13503_ VGND VGND VPWR VPWR _13504_ sky130_fd_sc_hd__clkbuf_4
X_29729_ net1075 _01464_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[22\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_17743_ _13263_ net3346 _05140_ VGND VGND VPWR VPWR _05147_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_1309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_193_5124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32740_ clknet_leaf_253_clk _04162_ VGND VGND VPWR VPWR datamem.data_ram\[16\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14886_ rvcpu.dp.pcreg.q\[8\] VGND VGND VPWR VPWR _13438_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_193_5135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17674_ _05110_ VGND VGND VPWR VPWR _01202_ sky130_fd_sc_hd__clkbuf_1
X_19413_ datamem.data_ram\[0\]\[16\] _06698_ _06701_ datamem.data_ram\[1\]\[16\] _06708_
+ VGND VGND VPWR VPWR _06709_ sky130_fd_sc_hd__o221a_1
X_16625_ _04554_ VGND VGND VPWR VPWR _01727_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_212_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32671_ clknet_leaf_284_clk _04093_ VGND VGND VPWR VPWR datamem.data_ram\[19\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap80 _12242_ VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__buf_4
XFILLER_0_174_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31622_ clknet_leaf_65_clk net1202 VGND VGND VPWR VPWR rvcpu.dp.plmw.lAuiPCW\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_175_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19344_ net1 _05371_ VGND VGND VPWR VPWR _06640_ sky130_fd_sc_hd__nor2_8
X_16556_ _04517_ VGND VGND VPWR VPWR _01767_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15507_ _13322_ _13492_ _13394_ VGND VGND VPWR VPWR _14034_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_14_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31553_ clknet_leaf_63_clk datamem.rd_data_mem\[3\] VGND VGND VPWR VPWR rvcpu.dp.plmw.ReadDataW\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_19275_ rvcpu.dp.plfd.InstrD\[13\] rvcpu.dp.plfd.InstrD\[12\] VGND VGND VPWR VPWR
+ _06574_ sky130_fd_sc_hd__and2b_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_16487_ net2734 _14447_ _04478_ VGND VGND VPWR VPWR _04481_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_152_4142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_4153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15438_ _13533_ _13359_ _13829_ VGND VGND VPWR VPWR _13969_ sky130_fd_sc_hd__or3b_1
X_18226_ _05590_ _05365_ VGND VGND VPWR VPWR _05591_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30504_ clknet_leaf_271_clk _02239_ VGND VGND VPWR VPWR datamem.data_ram\[57\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_31484_ clknet_leaf_48_clk rvcpu.dp.lAuiPCE\[10\] VGND VGND VPWR VPWR rvcpu.dp.plem.lAuiPCM\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_980 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22980__687 clknet_1_0__leaf__10083_ VGND VGND VPWR VPWR net813 sky130_fd_sc_hd__inv_2
XFILLER_0_53_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30435_ net773 _02170_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[29\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_15369_ _13903_ VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__inv_2
X_18157_ _05458_ _05466_ _05459_ VGND VGND VPWR VPWR _05522_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_26_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__10263_ clknet_0__10263_ VGND VGND VPWR VPWR clknet_1_0__leaf__10263_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_4_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold304 datamem.data_ram\[23\]\[0\] VGND VGND VPWR VPWR net1454 sky130_fd_sc_hd__dlygate4sd3_1
X_17108_ _04810_ VGND VGND VPWR VPWR _01484_ sky130_fd_sc_hd__clkbuf_1
Xhold315 datamem.data_ram\[58\]\[6\] VGND VGND VPWR VPWR net1465 sky130_fd_sc_hd__dlygate4sd3_1
X_18088_ rvcpu.dp.plde.RD1E\[23\] _05292_ _05455_ VGND VGND VPWR VPWR _05456_ sky130_fd_sc_hd__o21a_2
X_30366_ net712 _02101_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[3\]\[17\] sky130_fd_sc_hd__dfxtp_1
Xhold326 datamem.data_ram\[11\]\[7\] VGND VGND VPWR VPWR net1476 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_229_5982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold337 datamem.data_ram\[28\]\[3\] VGND VGND VPWR VPWR net1487 sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 datamem.data_ram\[1\]\[5\] VGND VGND VPWR VPWR net1498 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__10194_ clknet_0__10194_ VGND VGND VPWR VPWR clknet_1_0__leaf__10194_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_229_5993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32105_ clknet_leaf_120_clk _03527_ VGND VGND VPWR VPWR datamem.data_ram\[58\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17039_ net3626 _14453_ _04768_ VGND VGND VPWR VPWR _04774_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold359 datamem.data_ram\[5\]\[6\] VGND VGND VPWR VPWR net1509 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_111_3171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30297_ net643 _02032_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[5\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_23353__990 clknet_1_0__leaf__10137_ VGND VGND VPWR VPWR net1116 sky130_fd_sc_hd__inv_2
X_32036_ clknet_leaf_131_clk _03458_ VGND VGND VPWR VPWR datamem.data_ram\[50\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20050_ datamem.data_ram\[34\]\[26\] _06608_ _06644_ datamem.data_ram\[32\]\[26\]
+ VGND VGND VPWR VPWR _07344_ sky130_fd_sc_hd__o22a_1
XFILLER_0_102_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_182_4861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_4872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24177__18 clknet_1_0__leaf__10265_ VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__inv_2
XFILLER_0_175_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1004 rvcpu.dp.rf.reg_file_arr\[6\]\[2\] VGND VGND VPWR VPWR net2154 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1015 rvcpu.dp.rf.reg_file_arr\[23\]\[21\] VGND VGND VPWR VPWR net2165 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1026 rvcpu.dp.rf.reg_file_arr\[7\]\[17\] VGND VGND VPWR VPWR net2176 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1037 rvcpu.dp.rf.reg_file_arr\[22\]\[2\] VGND VGND VPWR VPWR net2187 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1048 rvcpu.dp.rf.reg_file_arr\[3\]\[7\] VGND VGND VPWR VPWR net2198 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_213_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1059 datamem.data_ram\[36\]\[15\] VGND VGND VPWR VPWR net2209 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_206_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_159_4307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_4318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20952_ _06988_ _08069_ _08241_ VGND VGND VPWR VPWR _04443_ sky130_fd_sc_hd__a21bo_1
X_32938_ clknet_leaf_156_clk _04360_ VGND VGND VPWR VPWR datamem.data_ram\[6\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_3890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32869_ clknet_leaf_286_clk _04291_ VGND VGND VPWR VPWR datamem.data_ram\[11\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_81_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20883_ datamem.data_ram\[56\]\[14\] _06837_ _06829_ datamem.data_ram\[59\]\[14\]
+ _06714_ VGND VGND VPWR VPWR _08173_ sky130_fd_sc_hd__o221a_1
XFILLER_0_221_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25410_ _10932_ net104 VGND VGND VPWR VPWR _10960_ sky130_fd_sc_hd__nor2_8
XTAP_TAPCELL_ROW_81_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22622_ _09622_ _09769_ _09771_ VGND VGND VPWR VPWR _09772_ sky130_fd_sc_hd__a21o_1
XFILLER_0_192_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26390_ rvcpu.dp.plde.JalrE VGND VGND VPWR VPWR _11535_ sky130_fd_sc_hd__buf_2
X_23853__416 clknet_1_0__leaf__10219_ VGND VGND VPWR VPWR net542 sky130_fd_sc_hd__inv_2
XFILLER_0_220_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25341_ _10916_ VGND VGND VPWR VPWR _02714_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22553_ rvcpu.dp.rf.reg_file_arr\[16\]\[13\] rvcpu.dp.rf.reg_file_arr\[17\]\[13\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[13\] rvcpu.dp.rf.reg_file_arr\[19\]\[13\] _09384_
+ _09577_ VGND VGND VPWR VPWR _09706_ sky130_fd_sc_hd__mux4_1
XFILLER_0_1_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26492__45 clknet_1_1__leaf__11601_ VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_118_3336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28060_ _12359_ net3652 _12492_ VGND VGND VPWR VPWR _12494_ sky130_fd_sc_hd__mux2_1
X_21504_ _08751_ _08755_ _08759_ _08625_ VGND VGND VPWR VPWR _01034_ sky130_fd_sc_hd__o31a_1
XFILLER_0_1_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25272_ _10741_ _10092_ _10828_ VGND VGND VPWR VPWR _10878_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_17_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22484_ _09495_ _09640_ _09457_ VGND VGND VPWR VPWR _09641_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_106_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27011_ _11803_ _11886_ VGND VGND VPWR VPWR _11892_ sky130_fd_sc_hd__and2_1
XFILLER_0_173_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24223_ _10282_ VGND VGND VPWR VPWR _02230_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21435_ rvcpu.dp.rf.reg_file_arr\[8\]\[3\] rvcpu.dp.rf.reg_file_arr\[10\]\[3\] rvcpu.dp.rf.reg_file_arr\[9\]\[3\]
+ rvcpu.dp.rf.reg_file_arr\[11\]\[3\] _08693_ _08578_ VGND VGND VPWR VPWR _08694_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_146_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21366_ _08626_ VGND VGND VPWR VPWR _08627_ sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_169_Right_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20317_ datamem.data_ram\[14\]\[4\] _07159_ _07605_ _07608_ VGND VGND VPWR VPWR _07609_
+ sky130_fd_sc_hd__a211o_1
X_28962_ _10325_ _10049_ _11898_ VGND VGND VPWR VPWR _12989_ sky130_fd_sc_hd__and3_2
X_24085_ _10254_ VGND VGND VPWR VPWR _02120_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21297_ rvcpu.dp.plfd.InstrD\[16\] VGND VGND VPWR VPWR _08559_ sky130_fd_sc_hd__clkbuf_8
Xhold860 datamem.data_ram\[34\]\[31\] VGND VGND VPWR VPWR net2010 sky130_fd_sc_hd__dlygate4sd3_1
Xhold871 rvcpu.dp.rf.reg_file_arr\[7\]\[14\] VGND VGND VPWR VPWR net2021 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold882 datamem.data_ram\[10\]\[23\] VGND VGND VPWR VPWR net2032 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold893 rvcpu.dp.rf.reg_file_arr\[20\]\[14\] VGND VGND VPWR VPWR net2043 sky130_fd_sc_hd__dlygate4sd3_1
X_27913_ _12151_ net2976 net47 VGND VGND VPWR VPWR _12408_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20248_ datamem.data_ram\[38\]\[3\] _06952_ _06958_ datamem.data_ram\[33\]\[3\] _07540_
+ VGND VGND VPWR VPWR _07541_ sky130_fd_sc_hd__a221o_1
XFILLER_0_200_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28893_ _12951_ VGND VGND VPWR VPWR _04231_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_194_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20179_ datamem.data_ram\[15\]\[11\] _06761_ _07024_ datamem.data_ram\[12\]\[11\]
+ VGND VGND VPWR VPWR _07472_ sky130_fd_sc_hd__o22a_1
X_27844_ _09325_ VGND VGND VPWR VPWR _12369_ sky130_fd_sc_hd__clkbuf_2
Xhold2250 datamem.data_ram\[40\]\[9\] VGND VGND VPWR VPWR net3400 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2261 datamem.data_ram\[50\]\[12\] VGND VGND VPWR VPWR net3411 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2272 datamem.data_ram\[10\]\[22\] VGND VGND VPWR VPWR net3422 sky130_fd_sc_hd__dlygate4sd3_1
X_27775_ _12328_ VGND VGND VPWR VPWR _03736_ sky130_fd_sc_hd__clkbuf_1
Xhold2283 datamem.data_ram\[60\]\[8\] VGND VGND VPWR VPWR net3433 sky130_fd_sc_hd__dlygate4sd3_1
X_24987_ _10480_ net2089 net101 VGND VGND VPWR VPWR _10714_ sky130_fd_sc_hd__mux2_1
XFILLER_0_216_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2294 datamem.data_ram\[40\]\[18\] VGND VGND VPWR VPWR net3444 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1560 datamem.data_ram\[45\]\[8\] VGND VGND VPWR VPWR net2710 sky130_fd_sc_hd__dlygate4sd3_1
X_14740_ rvcpu.dp.pcreg.q\[5\] _13281_ VGND VGND VPWR VPWR _13293_ sky130_fd_sc_hd__and2_1
Xhold1571 datamem.data_ram\[46\]\[28\] VGND VGND VPWR VPWR net2721 sky130_fd_sc_hd__dlygate4sd3_1
X_29514_ net876 _01249_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[28\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_26726_ _10760_ net2319 _11714_ VGND VGND VPWR VPWR _11719_ sky130_fd_sc_hd__mux2_1
Xhold1582 datamem.data_ram\[60\]\[28\] VGND VGND VPWR VPWR net2732 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1593 rvcpu.dp.rf.reg_file_arr\[30\]\[1\] VGND VGND VPWR VPWR net2743 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26657_ _11676_ _11677_ VGND VGND VPWR VPWR _11678_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_47_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14671_ _13237_ VGND VGND VPWR VPWR _13238_ sky130_fd_sc_hd__buf_4
X_29445_ net807 _01180_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[30\]\[16\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__10226_ clknet_0__10226_ VGND VGND VPWR VPWR clknet_1_1__leaf__10226_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_200_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16410_ net1984 _14440_ _14561_ VGND VGND VPWR VPWR _14571_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23029__731 clknet_1_1__leaf__10088_ VGND VGND VPWR VPWR net857 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_103_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25608_ _11068_ VGND VGND VPWR VPWR _02829_ sky130_fd_sc_hd__clkbuf_1
X_17390_ _04937_ VGND VGND VPWR VPWR _04960_ sky130_fd_sc_hd__clkbuf_4
X_26588_ _11078_ _11640_ VGND VGND VPWR VPWR _11641_ sky130_fd_sc_hd__and2_1
XFILLER_0_156_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29376_ clknet_leaf_144_clk _01111_ VGND VGND VPWR VPWR datamem.data_ram\[60\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__10157_ clknet_0__10157_ VGND VGND VPWR VPWR clknet_1_1__leaf__10157_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_200_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_530 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16341_ _14534_ VGND VGND VPWR VPWR _01867_ sky130_fd_sc_hd__clkbuf_1
X_28327_ _12637_ VGND VGND VPWR VPWR _03979_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25539_ _11027_ VGND VGND VPWR VPWR _02801_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__10088_ clknet_0__10088_ VGND VGND VPWR VPWR clknet_1_1__leaf__10088_
+ sky130_fd_sc_hd__clkbuf_16
X_19060_ rvcpu.dp.plde.ImmExtE\[6\] rvcpu.dp.plde.PCE\[6\] VGND VGND VPWR VPWR _06387_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_164_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16272_ net3998 _14438_ _14489_ VGND VGND VPWR VPWR _14498_ sky130_fd_sc_hd__mux2_1
X_28258_ _12460_ net4344 net44 VGND VGND VPWR VPWR _12599_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15223_ _13332_ _13763_ _13721_ VGND VGND VPWR VPWR _13764_ sky130_fd_sc_hd__or3_2
X_27209_ _12005_ net1572 _12007_ _12014_ VGND VGND VPWR VPWR _03484_ sky130_fd_sc_hd__a31o_1
XFILLER_0_180_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18011_ net122 _05268_ _05269_ _13271_ VGND VGND VPWR VPWR _05381_ sky130_fd_sc_hd__a22o_1
XFILLER_0_168_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28189_ _12443_ net4397 _12555_ VGND VGND VPWR VPWR _12562_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30220_ net574 _01955_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[7\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15154_ _13506_ _13472_ VGND VGND VPWR VPWR _13698_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_205_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_136_Right_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30151_ net513 _01886_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[0\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15085_ _13447_ _13630_ VGND VGND VPWR VPWR _13631_ sky130_fd_sc_hd__nor2_1
X_19962_ datamem.data_ram\[6\]\[18\] _06628_ _06806_ datamem.data_ram\[4\]\[18\] VGND
+ VGND VPWR VPWR _07256_ sky130_fd_sc_hd__o22a_1
X_18913_ _05619_ _05620_ _05629_ _06252_ VGND VGND VPWR VPWR _06253_ sky130_fd_sc_hd__a211o_1
XFILLER_0_226_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30082_ net444 _01817_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[11\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_19893_ datamem.data_ram\[19\]\[17\] _06739_ _06621_ datamem.data_ram\[20\]\[17\]
+ _07187_ VGND VGND VPWR VPWR _07188_ sky130_fd_sc_hd__o221a_1
XFILLER_0_219_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18844_ _05488_ _05728_ _06180_ _06187_ _06188_ VGND VGND VPWR VPWR _06189_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_8_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_220_5765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_220_5776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18775_ _05318_ _06123_ VGND VGND VPWR VPWR _06124_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24093__602 clknet_1_0__leaf__10248_ VGND VGND VPWR VPWR net728 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_220_5787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15987_ net1964 _13238_ _14322_ VGND VGND VPWR VPWR _14331_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17726_ _13238_ net2845 _05129_ VGND VGND VPWR VPWR _05138_ sky130_fd_sc_hd__mux2_1
X_14938_ _13287_ _13281_ VGND VGND VPWR VPWR _13487_ sky130_fd_sc_hd__and2_1
XFILLER_0_145_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30984_ clknet_leaf_115_clk _02719_ VGND VGND VPWR VPWR datamem.data_ram\[39\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_216_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_203_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_19_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32723_ clknet_leaf_239_clk _04145_ VGND VGND VPWR VPWR datamem.data_ram\[16\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17657_ _05101_ VGND VGND VPWR VPWR _01210_ sky130_fd_sc_hd__clkbuf_1
X_14869_ _13358_ _13420_ VGND VGND VPWR VPWR _13421_ sky130_fd_sc_hd__nand2_1
XFILLER_0_159_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16608_ _04545_ VGND VGND VPWR VPWR _01735_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32654_ clknet_leaf_243_clk _04076_ VGND VGND VPWR VPWR datamem.data_ram\[19\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_17588_ _13235_ net3694 _05057_ VGND VGND VPWR VPWR _05065_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31605_ clknet_leaf_28_clk net1197 VGND VGND VPWR VPWR rvcpu.dp.plmw.PCPlus4W\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19327_ _06622_ _06606_ VGND VGND VPWR VPWR _06623_ sky130_fd_sc_hd__nor2_8
XFILLER_0_9_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16539_ _04508_ VGND VGND VPWR VPWR _01775_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32585_ clknet_leaf_75_clk _04007_ VGND VGND VPWR VPWR datamem.data_ram\[21\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19258_ _06548_ _06555_ _06556_ _06553_ VGND VGND VPWR VPWR _06560_ sky130_fd_sc_hd__a31o_1
X_31536_ clknet_leaf_18_clk net1218 VGND VGND VPWR VPWR rvcpu.dp.plem.PCPlus4M\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_171_4595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18209_ rvcpu.dp.plde.RD1E\[19\] _05564_ _05483_ VGND VGND VPWR VPWR _05574_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_113_3200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_3211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19189_ _06500_ VGND VGND VPWR VPWR rvcpu.dp.lAuiPCE\[21\] sky130_fd_sc_hd__clkbuf_1
X_31467_ clknet_leaf_2_clk rvcpu.dp.SrcBFW_Mux.y\[25\] VGND VGND VPWR VPWR rvcpu.dp.plem.WriteDataM\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21220_ _06862_ _08487_ _08490_ VGND VGND VPWR VPWR _04431_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_184_4901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold101 rvcpu.dp.plem.RdM\[0\] VGND VGND VPWR VPWR net1251 sky130_fd_sc_hd__dlygate4sd3_1
X_30418_ net756 _02153_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[31\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_223_1210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31398_ clknet_leaf_49_clk _03101_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCE\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_184_4912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold112 rvcpu.dp.plem.RdM\[3\] VGND VGND VPWR VPWR net1262 sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 rvcpu.dp.plde.RdE\[1\] VGND VGND VPWR VPWR net1273 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__10246_ clknet_0__10246_ VGND VGND VPWR VPWR clknet_1_0__leaf__10246_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_184_4923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold134 rvcpu.dp.plfd.PCD\[3\] VGND VGND VPWR VPWR net1284 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_103_Right_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold145 rvcpu.dp.plfd.PCD\[20\] VGND VGND VPWR VPWR net1295 sky130_fd_sc_hd__dlygate4sd3_1
X_21151_ datamem.data_ram\[18\]\[23\] _06608_ _06631_ datamem.data_ram\[19\]\[23\]
+ _06676_ VGND VGND VPWR VPWR _08440_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_74_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold156 rvcpu.dp.plfd.InstrD\[27\] VGND VGND VPWR VPWR net1306 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30349_ net695 _02084_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[3\]\[0\] sky130_fd_sc_hd__dfxtp_1
Xhold167 datamem.data_ram\[42\]\[2\] VGND VGND VPWR VPWR net1317 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__10177_ clknet_0__10177_ VGND VGND VPWR VPWR clknet_1_0__leaf__10177_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_223_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold178 datamem.data_ram\[41\]\[0\] VGND VGND VPWR VPWR net1328 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_180_4809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20102_ datamem.data_ram\[13\]\[10\] _06724_ _06697_ datamem.data_ram\[8\]\[10\]
+ VGND VGND VPWR VPWR _07396_ sky130_fd_sc_hd__o22a_1
X_21082_ _07823_ datamem.data_ram\[39\]\[7\] _07825_ datamem.data_ram\[38\]\[7\] _07866_
+ VGND VGND VPWR VPWR _08371_ sky130_fd_sc_hd__o221a_1
Xhold189 datamem.data_ram\[46\]\[7\] VGND VGND VPWR VPWR net1339 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20033_ datamem.data_ram\[29\]\[26\] _06702_ _06741_ _07326_ VGND VGND VPWR VPWR
+ _07327_ sky130_fd_sc_hd__o211a_1
X_24910_ _10392_ net3112 _10669_ VGND VGND VPWR VPWR _10673_ sky130_fd_sc_hd__mux2_1
X_32019_ clknet_leaf_129_clk _03441_ VGND VGND VPWR VPWR datamem.data_ram\[51\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_6_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25890_ _13665_ _11256_ _11258_ _11262_ VGND VGND VPWR VPWR _02917_ sky130_fd_sc_hd__o211a_1
XFILLER_0_226_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_143_3930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24841_ _10635_ VGND VGND VPWR VPWR _02495_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_107_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27560_ _12155_ net3358 _12206_ VGND VGND VPWR VPWR _12213_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24772_ _10478_ net3420 _10589_ VGND VGND VPWR VPWR _10596_ sky130_fd_sc_hd__mux2_1
X_21984_ _06582_ _09213_ VGND VGND VPWR VPWR _09214_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_205_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20935_ _06681_ _08217_ _08224_ VGND VGND VPWR VPWR _08225_ sky130_fd_sc_hd__o21a_1
X_27491_ _12138_ net2325 _12169_ VGND VGND VPWR VPWR _12176_ sky130_fd_sc_hd__mux2_1
Xclkbuf_0__10111_ _10111_ VGND VGND VPWR VPWR clknet_0__10111_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_178_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26442_ net2078 _11542_ _11572_ _11570_ VGND VGND VPWR VPWR _03159_ sky130_fd_sc_hd__o211a_1
XFILLER_0_166_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29230_ _09309_ net2206 _13132_ VGND VGND VPWR VPWR _13135_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20866_ datamem.data_ram\[33\]\[14\] _06934_ VGND VGND VPWR VPWR _08156_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29161_ _13097_ VGND VGND VPWR VPWR _04353_ sky130_fd_sc_hd__clkbuf_1
X_22605_ rvcpu.dp.rf.reg_file_arr\[12\]\[15\] rvcpu.dp.rf.reg_file_arr\[13\]\[15\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[15\] rvcpu.dp.rf.reg_file_arr\[15\]\[15\] _09552_
+ _09721_ VGND VGND VPWR VPWR _09756_ sky130_fd_sc_hd__mux4_1
XFILLER_0_7_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26373_ _08620_ _08621_ rvcpu.dp.plde.JalrE VGND VGND VPWR VPWR _11521_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_166_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20797_ _08085_ _08086_ _07822_ VGND VGND VPWR VPWR _08087_ sky130_fd_sc_hd__mux2_1
XFILLER_0_221_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28112_ _12521_ VGND VGND VPWR VPWR _03880_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25324_ _10826_ net1948 _10899_ VGND VGND VPWR VPWR _10907_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_3778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22536_ _09688_ _09689_ _09421_ VGND VGND VPWR VPWR _09690_ sky130_fd_sc_hd__mux2_2
XFILLER_0_9_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29092_ _09309_ net2898 _13058_ VGND VGND VPWR VPWR _13061_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_137_3789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28043_ _12450_ net2790 net96 VGND VGND VPWR VPWR _12485_ sky130_fd_sc_hd__mux2_1
X_25255_ _10405_ _10868_ VGND VGND VPWR VPWR _10869_ sky130_fd_sc_hd__and2_1
XFILLER_0_134_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22467_ _09528_ _09624_ _09426_ VGND VGND VPWR VPWR _09625_ sky130_fd_sc_hd__a21o_1
XFILLER_0_161_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24206_ _10273_ VGND VGND VPWR VPWR _02222_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21418_ _08531_ _08676_ _08512_ VGND VGND VPWR VPWR _08677_ sky130_fd_sc_hd__o21a_1
X_25186_ _10727_ net4086 _10829_ VGND VGND VPWR VPWR _10831_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22398_ rvcpu.dp.rf.reg_file_arr\[20\]\[5\] rvcpu.dp.rf.reg_file_arr\[21\]\[5\] rvcpu.dp.rf.reg_file_arr\[22\]\[5\]
+ rvcpu.dp.rf.reg_file_arr\[23\]\[5\] _09434_ _09558_ VGND VGND VPWR VPWR _09559_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_103_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21349_ rvcpu.ALUResultE\[31\] rvcpu.ALUResultE\[30\] _08599_ _08610_ VGND VGND VPWR
+ VPWR _08611_ sky130_fd_sc_hd__or4_1
XFILLER_0_20_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29994_ net364 _01729_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[14\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28945_ _12979_ VGND VGND VPWR VPWR _04255_ sky130_fd_sc_hd__clkbuf_1
X_24068_ clknet_1_1__leaf__10244_ VGND VGND VPWR VPWR _10248_ sky130_fd_sc_hd__buf_1
Xhold690 rvcpu.dp.plfd.PCD\[11\] VGND VGND VPWR VPWR net1840 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15910_ _14290_ VGND VGND VPWR VPWR _02070_ sky130_fd_sc_hd__clkbuf_1
X_28876_ _12942_ VGND VGND VPWR VPWR _04223_ sky130_fd_sc_hd__clkbuf_1
X_16890_ _04694_ VGND VGND VPWR VPWR _01594_ sky130_fd_sc_hd__clkbuf_1
X_27827_ _12355_ net2338 _12357_ VGND VGND VPWR VPWR _12358_ sky130_fd_sc_hd__mux2_1
X_15841_ _14252_ VGND VGND VPWR VPWR _02101_ sky130_fd_sc_hd__clkbuf_1
Xhold2080 datamem.data_ram\[14\]\[29\] VGND VGND VPWR VPWR net3230 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2091 datamem.data_ram\[20\]\[31\] VGND VGND VPWR VPWR net3241 sky130_fd_sc_hd__dlygate4sd3_1
X_18560_ _05674_ _05766_ VGND VGND VPWR VPWR _05920_ sky130_fd_sc_hd__nor2_1
XFILLER_0_188_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27758_ _12147_ net2771 net48 VGND VGND VPWR VPWR _12319_ sky130_fd_sc_hd__mux2_1
X_15772_ _14215_ VGND VGND VPWR VPWR _02141_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_188_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1390 datamem.data_ram\[58\]\[12\] VGND VGND VPWR VPWR net2540 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17511_ _05024_ VGND VGND VPWR VPWR _01287_ sky130_fd_sc_hd__clkbuf_1
X_14723_ rvcpu.dp.plmw.ALUResultW\[0\] rvcpu.dp.plmw.ReadDataW\[0\] rvcpu.dp.plmw.PCPlus4W\[0\]
+ rvcpu.dp.plmw.lAuiPCW\[0\] rvcpu.dp.plmw.ResultSrcW\[0\] rvcpu.dp.plmw.ResultSrcW\[1\]
+ VGND VGND VPWR VPWR _13277_ sky130_fd_sc_hd__mux4_2
XFILLER_0_8_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26709_ _11709_ VGND VGND VPWR VPWR _03289_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18491_ _05852_ _05770_ _05768_ VGND VGND VPWR VPWR _05853_ sky130_fd_sc_hd__mux2_1
X_27689_ _12282_ VGND VGND VPWR VPWR _03696_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_530 _14432_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_197_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_541 _06706_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_552 _07635_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_200_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14654_ rvcpu.dp.plmw.ALUResultW\[17\] rvcpu.dp.plmw.ReadDataW\[17\] rvcpu.dp.plmw.PCPlus4W\[17\]
+ rvcpu.dp.plmw.lAuiPCW\[17\] _13169_ _13171_ VGND VGND VPWR VPWR _13225_ sky130_fd_sc_hd__mux4_2
X_29428_ clknet_leaf_85_clk _01163_ VGND VGND VPWR VPWR datamem.data_ram\[5\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17442_ _14156_ net4237 _04985_ VGND VGND VPWR VPWR _04988_ sky130_fd_sc_hd__mux2_1
XANTENNA_563 _11970_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_205_Right_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_185_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14585_ rvcpu.dp.plmw.ResultSrcW\[1\] VGND VGND VPWR VPWR _13170_ sky130_fd_sc_hd__buf_4
X_29359_ clknet_leaf_266_clk _01094_ VGND VGND VPWR VPWR datamem.data_ram\[61\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_17373_ _04951_ VGND VGND VPWR VPWR _01352_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_184_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19112_ _06432_ rvcpu.dp.plde.ImmExtE\[12\] _06419_ VGND VGND VPWR VPWR _06433_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_188_5001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_188_5012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16324_ net1917 _14420_ _14525_ VGND VGND VPWR VPWR _14526_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32370_ clknet_leaf_260_clk _03792_ VGND VGND VPWR VPWR datamem.data_ram\[2\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19043_ _06372_ VGND VGND VPWR VPWR rvcpu.dp.lAuiPCE\[3\] sky130_fd_sc_hd__clkbuf_1
X_31321_ clknet_leaf_25_clk _03024_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCPlus4E\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16255_ _14488_ VGND VGND VPWR VPWR _14489_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_152_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15206_ _13391_ _13523_ _13747_ VGND VGND VPWR VPWR _13748_ sky130_fd_sc_hd__a21o_1
XFILLER_0_125_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31252_ clknet_leaf_21_clk _02955_ VGND VGND VPWR VPWR rvcpu.dp.plfd.InstrD\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16186_ _13212_ VGND VGND VPWR VPWR _14442_ sky130_fd_sc_hd__buf_4
XFILLER_0_207_1249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_226_5930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15137_ _13546_ VGND VGND VPWR VPWR _13681_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30203_ net557 _01938_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[8\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31183_ clknet_leaf_32_clk _02886_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCPlus4D\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_147_4030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30134_ net496 _01869_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[10\]\[25\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_222_5816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15068_ _13331_ _13562_ _13613_ VGND VGND VPWR VPWR _13614_ sky130_fd_sc_hd__or3_1
X_19945_ datamem.data_ram\[43\]\[18\] _06636_ _07235_ _07238_ VGND VGND VPWR VPWR
+ _07239_ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_227_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_222_5827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30065_ net427 _01800_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[12\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19876_ datamem.data_ram\[21\]\[1\] _06970_ _06977_ datamem.data_ram\[20\]\[1\] VGND
+ VGND VPWR VPWR _07171_ sky130_fd_sc_hd__a22o_1
XFILLER_0_177_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23581__203 clknet_1_1__leaf__10176_ VGND VGND VPWR VPWR net329 sky130_fd_sc_hd__inv_2
X_18827_ _06112_ _06172_ _05706_ VGND VGND VPWR VPWR _06173_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_222_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18758_ _05974_ VGND VGND VPWR VPWR _06108_ sky130_fd_sc_hd__buf_2
X_23661__260 clknet_1_1__leaf__10191_ VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__inv_2
XFILLER_0_222_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24058__585 clknet_1_0__leaf__10247_ VGND VGND VPWR VPWR net711 sky130_fd_sc_hd__inv_2
XFILLER_0_76_1180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17709_ _05117_ VGND VGND VPWR VPWR _05129_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_222_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18689_ _05781_ _05841_ _05857_ _05775_ VGND VGND VPWR VPWR _06043_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30967_ clknet_leaf_207_clk _02702_ VGND VGND VPWR VPWR datamem.data_ram\[39\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20720_ _06985_ _07987_ _08010_ VGND VGND VPWR VPWR _08011_ sky130_fd_sc_hd__o21ai_2
X_32706_ clknet_leaf_87_clk _04128_ VGND VGND VPWR VPWR datamem.data_ram\[17\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_173_4646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30898_ clknet_leaf_137_clk _02633_ VGND VGND VPWR VPWR datamem.data_ram\[41\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_22986__693 clknet_1_1__leaf__10083_ VGND VGND VPWR VPWR net819 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_173_4657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32637_ clknet_leaf_286_clk _04059_ VGND VGND VPWR VPWR datamem.data_ram\[1\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_20651_ datamem.data_ram\[37\]\[29\] _07037_ _06784_ datamem.data_ram\[39\]\[29\]
+ VGND VGND VPWR VPWR _07942_ sky130_fd_sc_hd__o22a_1
XFILLER_0_163_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32568_ clknet_leaf_171_clk _03990_ VGND VGND VPWR VPWR datamem.data_ram\[22\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_20582_ _07635_ datamem.data_ram\[51\]\[13\] _07831_ datamem.data_ram\[50\]\[13\]
+ VGND VGND VPWR VPWR _07873_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22321_ rvcpu.dp.rf.reg_file_arr\[8\]\[1\] rvcpu.dp.rf.reg_file_arr\[10\]\[1\] rvcpu.dp.rf.reg_file_arr\[9\]\[1\]
+ rvcpu.dp.rf.reg_file_arr\[11\]\[1\] _09483_ _09485_ VGND VGND VPWR VPWR _09486_
+ sky130_fd_sc_hd__mux4_1
X_31519_ clknet_leaf_48_clk net1160 VGND VGND VPWR VPWR rvcpu.dp.plem.PCPlus4M\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32499_ clknet_leaf_248_clk _03921_ VGND VGND VPWR VPWR datamem.data_ram\[25\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_76_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_3653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25040_ _10746_ VGND VGND VPWR VPWR _02583_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_3664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22252_ _09400_ VGND VGND VPWR VPWR _09418_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_132_3675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21203_ _06915_ _08123_ _08182_ _07277_ VGND VGND VPWR VPWR _08484_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_44_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22183_ _09236_ net3752 _09362_ VGND VGND VPWR VPWR _09364_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_223_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21134_ datamem.data_ram\[54\]\[23\] _06717_ _06725_ datamem.data_ram\[55\]\[23\]
+ _06732_ VGND VGND VPWR VPWR _08423_ sky130_fd_sc_hd__o221a_1
XFILLER_0_44_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26991_ _10760_ net4214 _11875_ VGND VGND VPWR VPWR _11880_ sky130_fd_sc_hd__mux2_1
Xclkbuf_2_2_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_2_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_35_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28730_ _12864_ VGND VGND VPWR VPWR _04155_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25942_ net1847 _11279_ VGND VGND VPWR VPWR _11293_ sky130_fd_sc_hd__or2_1
X_21065_ _08299_ _08353_ _06911_ VGND VGND VPWR VPWR _08354_ sky130_fd_sc_hd__mux2_1
X_20016_ datamem.data_ram\[37\]\[2\] _06919_ _06947_ datamem.data_ram\[33\]\[2\] VGND
+ VGND VPWR VPWR _07310_ sky130_fd_sc_hd__a22o_1
X_25873_ _11206_ _11207_ _11250_ VGND VGND VPWR VPWR _11251_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_31_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28661_ _12696_ net2383 _12823_ VGND VGND VPWR VPWR _12828_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_31_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27612_ _12240_ VGND VGND VPWR VPWR _03661_ sky130_fd_sc_hd__clkbuf_1
X_24824_ _10394_ net3293 _10621_ VGND VGND VPWR VPWR _10626_ sky130_fd_sc_hd__mux2_1
XFILLER_0_216_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_213_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28592_ _12743_ net2905 _12786_ VGND VGND VPWR VPWR _12791_ sky130_fd_sc_hd__mux2_1
XFILLER_0_216_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_213_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23859__422 clknet_1_0__leaf__10219_ VGND VGND VPWR VPWR net548 sky130_fd_sc_hd__inv_2
XFILLER_0_201_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27543_ _12138_ net1925 _12197_ VGND VGND VPWR VPWR _12204_ sky130_fd_sc_hd__mux2_1
X_24755_ _10398_ net3160 _10580_ VGND VGND VPWR VPWR _10587_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21967_ _08522_ _09197_ _08512_ VGND VGND VPWR VPWR _09198_ sky130_fd_sc_hd__o21a_1
XFILLER_0_185_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_179_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20918_ _07860_ _08204_ _08207_ _07081_ VGND VGND VPWR VPWR _08208_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_100_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27474_ _12166_ VGND VGND VPWR VPWR _03597_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_139_3829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24686_ _10398_ net1956 _10543_ VGND VGND VPWR VPWR _10550_ sky130_fd_sc_hd__mux2_1
X_21898_ _08798_ _09130_ _09132_ _08512_ VGND VGND VPWR VPWR _09133_ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_193_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29213_ _10060_ _13123_ VGND VGND VPWR VPWR _13126_ sky130_fd_sc_hd__and2_1
X_26425_ _06447_ _11539_ _11529_ _11187_ _11560_ VGND VGND VPWR VPWR _11561_ sky130_fd_sc_hd__a221o_1
X_23637_ _09276_ net2565 _10182_ VGND VGND VPWR VPWR _10185_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_202_Left_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20849_ datamem.data_ram\[0\]\[14\] _06648_ _08138_ _07863_ VGND VGND VPWR VPWR _08139_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_166_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26356_ _11078_ _11511_ VGND VGND VPWR VPWR _11512_ sky130_fd_sc_hd__and2_1
X_29144_ _13088_ VGND VGND VPWR VPWR _04345_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_61_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25307_ _10896_ VGND VGND VPWR VPWR _10897_ sky130_fd_sc_hd__clkbuf_8
X_22519_ rvcpu.dp.rf.reg_file_arr\[24\]\[11\] rvcpu.dp.rf.reg_file_arr\[25\]\[11\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[11\] rvcpu.dp.rf.reg_file_arr\[27\]\[11\] _09463_
+ _09637_ VGND VGND VPWR VPWR _09674_ sky130_fd_sc_hd__mux4_1
XFILLER_0_18_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26287_ net1803 _11467_ VGND VGND VPWR VPWR _11476_ sky130_fd_sc_hd__and2_1
X_29075_ _12756_ net2819 _13049_ VGND VGND VPWR VPWR _13052_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23499_ clknet_1_0__leaf__10152_ VGND VGND VPWR VPWR _10161_ sky130_fd_sc_hd__buf_1
XFILLER_0_190_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16040_ _14348_ VGND VGND VPWR VPWR _14360_ sky130_fd_sc_hd__clkbuf_4
X_28026_ _12475_ VGND VGND VPWR VPWR _03840_ sky130_fd_sc_hd__clkbuf_1
X_25238_ _10727_ net3400 _10857_ VGND VGND VPWR VPWR _10859_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_21_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25169_ _10819_ VGND VGND VPWR VPWR _02639_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23530__157 clknet_1_1__leaf__10171_ VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_211_Left_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_209_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17991_ _05360_ VGND VGND VPWR VPWR _05361_ sky130_fd_sc_hd__inv_2
X_29977_ net347 _01712_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[14\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19730_ datamem.data_ram\[11\]\[25\] _06738_ _07024_ datamem.data_ram\[12\]\[25\]
+ VGND VGND VPWR VPWR _07025_ sky130_fd_sc_hd__o22a_1
X_28928_ _12754_ net3253 _12968_ VGND VGND VPWR VPWR _12970_ sky130_fd_sc_hd__mux2_1
X_16942_ _04722_ VGND VGND VPWR VPWR _01570_ sky130_fd_sc_hd__clkbuf_1
X_19661_ datamem.data_ram\[35\]\[0\] _06943_ _06949_ datamem.data_ram\[33\]\[0\] _06956_
+ VGND VGND VPWR VPWR _06957_ sky130_fd_sc_hd__a221o_1
XFILLER_0_217_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28859_ _12933_ VGND VGND VPWR VPWR _04215_ sky130_fd_sc_hd__clkbuf_1
X_16873_ net3987 _14424_ _04684_ VGND VGND VPWR VPWR _04686_ sky130_fd_sc_hd__mux2_1
XFILLER_0_189_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_205_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18612_ _05675_ _05856_ VGND VGND VPWR VPWR _05970_ sky130_fd_sc_hd__or2_1
X_15824_ _14243_ VGND VGND VPWR VPWR _02109_ sky130_fd_sc_hd__clkbuf_1
X_31870_ clknet_leaf_113_clk _03324_ VGND VGND VPWR VPWR datamem.data_ram\[63\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19592_ datamem.data_ram\[61\]\[8\] _06721_ _06654_ datamem.data_ram\[57\]\[8\] VGND
+ VGND VPWR VPWR _06888_ sky130_fd_sc_hd__o22a_1
Xclkbuf_5_24__f_clk clknet_2_3_0_clk VGND VGND VPWR VPWR clknet_5_24__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_205_879 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18543_ _05648_ _05642_ _05643_ _05636_ _05683_ _05688_ VGND VGND VPWR VPWR _05904_
+ sky130_fd_sc_hd__mux4_2
X_30821_ clknet_leaf_222_clk _02556_ VGND VGND VPWR VPWR datamem.data_ram\[44\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_15755_ _14206_ VGND VGND VPWR VPWR _02149_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14706_ _13264_ VGND VGND VPWR VPWR _03177_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_206_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18474_ _05836_ VGND VGND VPWR VPWR rvcpu.ALUResultE\[1\] sky130_fd_sc_hd__buf_1
X_30752_ clknet_leaf_189_clk _02487_ VGND VGND VPWR VPWR datamem.data_ram\[48\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_220_Left_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_360 rvcpu.dp.SrcBFW_Mux.y\[22\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15686_ _14161_ VGND VGND VPWR VPWR _02173_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_169_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_184_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_371 rvcpu.dp.plem.ALUResultM\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_382 net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_215_5653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17425_ _14139_ net4231 _04974_ VGND VGND VPWR VPWR _04979_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_215_5664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14637_ rvcpu.dp.plmw.ALUResultW\[21\] rvcpu.dp.plmw.ReadDataW\[21\] rvcpu.dp.plmw.PCPlus4W\[21\]
+ rvcpu.dp.plmw.lAuiPCW\[21\] _13169_ _13171_ VGND VGND VPWR VPWR _13212_ sky130_fd_sc_hd__mux4_2
XFILLER_0_158_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_393 clknet_1_0__leaf__10108_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_30683_ clknet_leaf_84_clk _02418_ VGND VGND VPWR VPWR datamem.data_ram\[4\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32422_ clknet_leaf_74_clk _03844_ VGND VGND VPWR VPWR datamem.data_ram\[28\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17356_ _04942_ VGND VGND VPWR VPWR _01360_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16307_ _14516_ VGND VGND VPWR VPWR _01883_ sky130_fd_sc_hd__clkbuf_1
X_23691__286 clknet_1_1__leaf__10195_ VGND VGND VPWR VPWR net412 sky130_fd_sc_hd__inv_2
XFILLER_0_27_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32353_ clknet_leaf_248_clk _03775_ VGND VGND VPWR VPWR datamem.data_ram\[30\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_17287_ net4420 _13189_ _04902_ VGND VGND VPWR VPWR _04906_ sky130_fd_sc_hd__mux2_1
Xclkload302 clknet_1_1__leaf__10192_ VGND VGND VPWR VPWR clkload302/X sky130_fd_sc_hd__clkbuf_8
Xclkload10 clknet_5_11__leaf_clk VGND VGND VPWR VPWR clkload10/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_28_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload313 clknet_1_0__leaf__10180_ VGND VGND VPWR VPWR clkload313/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_71_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31304_ clknet_leaf_51_clk _03007_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCPlus4E\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_19026_ _06352_ _06357_ VGND VGND VPWR VPWR _06358_ sky130_fd_sc_hd__xnor2_1
Xclkload21 clknet_5_25__leaf_clk VGND VGND VPWR VPWR clkload21/Y sky130_fd_sc_hd__inv_12
Xclkload324 clknet_1_1__leaf__10079_ VGND VGND VPWR VPWR clkload324/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_207_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload32 clknet_leaf_12_clk VGND VGND VPWR VPWR clkload32/Y sky130_fd_sc_hd__clkinv_4
Xclkload335 clknet_1_1__leaf__10133_ VGND VGND VPWR VPWR clkload335/Y sky130_fd_sc_hd__clkinvlp_4
X_16238_ _14477_ VGND VGND VPWR VPWR _01921_ sky130_fd_sc_hd__clkbuf_1
X_32284_ clknet_leaf_257_clk _03706_ VGND VGND VPWR VPWR datamem.data_ram\[33\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload43 clknet_leaf_32_clk VGND VGND VPWR VPWR clkload43/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_140_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload346 clknet_1_1__leaf__10110_ VGND VGND VPWR VPWR clkload346/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload54 clknet_leaf_281_clk VGND VGND VPWR VPWR clkload54/Y sky130_fd_sc_hd__inv_8
Xclkload357 clknet_1_1__leaf__10083_ VGND VGND VPWR VPWR clkload357/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_141_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload65 clknet_leaf_170_clk VGND VGND VPWR VPWR clkload65/Y sky130_fd_sc_hd__clkinv_4
Xclkload76 clknet_leaf_33_clk VGND VGND VPWR VPWR clkload76/Y sky130_fd_sc_hd__inv_6
X_31235_ clknet_leaf_31_clk _02938_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCD\[24\] sky130_fd_sc_hd__dfxtp_1
Xclkload87 clknet_leaf_51_clk VGND VGND VPWR VPWR clkload87/Y sky130_fd_sc_hd__inv_6
XFILLER_0_207_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16169_ net2945 _14430_ _14422_ VGND VGND VPWR VPWR _14431_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_71_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload98 clknet_leaf_97_clk VGND VGND VPWR VPWR clkload98/Y sky130_fd_sc_hd__clkinv_1
XFILLER_0_100_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_220_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31166_ clknet_leaf_28_clk rvcpu.ALUResultE\[25\] VGND VGND VPWR VPWR rvcpu.dp.plem.ALUResultM\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_166_4472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_578 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_4483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_220_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2805 datamem.data_ram\[1\]\[17\] VGND VGND VPWR VPWR net3955 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19928_ datamem.data_ram\[50\]\[17\] _06613_ _07219_ _07222_ VGND VGND VPWR VPWR
+ _07223_ sky130_fd_sc_hd__o211a_1
X_30117_ net479 _01852_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[10\]\[8\] sky130_fd_sc_hd__dfxtp_1
Xhold2816 datamem.data_ram\[45\]\[12\] VGND VGND VPWR VPWR net3966 sky130_fd_sc_hd__dlygate4sd3_1
X_31097_ clknet_leaf_286_clk _02832_ VGND VGND VPWR VPWR datamem.data_ram\[9\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2827 datamem.data_ram\[59\]\[23\] VGND VGND VPWR VPWR net3977 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2838 datamem.data_ram\[36\]\[11\] VGND VGND VPWR VPWR net3988 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2849 datamem.data_ram\[41\]\[20\] VGND VGND VPWR VPWR net3999 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30048_ net410 _01783_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[12\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_19859_ _06750_ _06860_ VGND VGND VPWR VPWR _07154_ sky130_fd_sc_hd__nand2_8
XTAP_TAPCELL_ROW_179_4800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22870_ _09380_ _10005_ VGND VGND VPWR VPWR _10006_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_69_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_125_3490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21821_ rvcpu.dp.rf.reg_file_arr\[24\]\[23\] rvcpu.dp.rf.reg_file_arr\[25\]\[23\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[23\] rvcpu.dp.rf.reg_file_arr\[27\]\[23\] _08525_
+ _08528_ VGND VGND VPWR VPWR _09060_ sky130_fd_sc_hd__mux4_1
X_31999_ clknet_leaf_134_clk _03421_ VGND VGND VPWR VPWR datamem.data_ram\[52\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_65_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_222_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_65_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24540_ _10142_ _10327_ _10366_ VGND VGND VPWR VPWR _10466_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_188_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21752_ rvcpu.dp.rf.reg_file_arr\[0\]\[19\] rvcpu.dp.rf.reg_file_arr\[1\]\[19\] rvcpu.dp.rf.reg_file_arr\[2\]\[19\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[19\] _08810_ _08811_ VGND VGND VPWR VPWR _08995_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_121_3398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20703_ datamem.data_ram\[12\]\[5\] _06955_ _06958_ datamem.data_ram\[9\]\[5\] VGND
+ VGND VPWR VPWR _07994_ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24471_ _10425_ VGND VGND VPWR VPWR _02335_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_191_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21683_ rvcpu.dp.rf.reg_file_arr\[8\]\[15\] rvcpu.dp.rf.reg_file_arr\[10\]\[15\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[15\] rvcpu.dp.rf.reg_file_arr\[11\]\[15\] _08534_
+ _08818_ VGND VGND VPWR VPWR _08930_ sky130_fd_sc_hd__mux4_1
XFILLER_0_148_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26210_ net1785 _11442_ _03039_ _11443_ VGND VGND VPWR VPWR _03056_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23422_ clknet_1_1__leaf__10152_ VGND VGND VPWR VPWR _10154_ sky130_fd_sc_hd__buf_1
X_27190_ _11978_ _11996_ VGND VGND VPWR VPWR _12003_ sky130_fd_sc_hd__and2_1
XFILLER_0_190_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_3704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20634_ datamem.data_ram\[14\]\[29\] _06627_ _06781_ datamem.data_ram\[9\]\[29\]
+ VGND VGND VPWR VPWR _07925_ sky130_fd_sc_hd__o22a_1
XFILLER_0_110_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_134_3715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire108 net109 VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__buf_2
Xclkload4 clknet_5_5__leaf_clk VGND VGND VPWR VPWR clkload4/Y sky130_fd_sc_hd__inv_8
XFILLER_0_11_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26141_ _11406_ VGND VGND VPWR VPWR _03023_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20565_ _07177_ _07813_ _07818_ _07855_ VGND VGND VPWR VPWR _07856_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_24_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22304_ _09391_ VGND VGND VPWR VPWR _09469_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_190_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26072_ rvcpu.dp.plfd.InstrD\[4\] rvcpu.c.ad.opb5 rvcpu.dp.plfd.InstrD\[6\] VGND
+ VGND VPWR VPWR _11366_ sky130_fd_sc_hd__and3b_1
XFILLER_0_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20496_ datamem.data_ram\[37\]\[21\] _06665_ _07021_ datamem.data_ram\[39\]\[21\]
+ _07786_ VGND VGND VPWR VPWR _07787_ sky130_fd_sc_hd__o221a_1
X_24108__615 clknet_1_0__leaf__10259_ VGND VGND VPWR VPWR net741 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_95_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29900_ net278 _01635_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[17\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_25023_ _10735_ net3953 net100 VGND VGND VPWR VPWR _10736_ sky130_fd_sc_hd__mux2_1
X_23588__209 clknet_1_0__leaf__10177_ VGND VGND VPWR VPWR net335 sky130_fd_sc_hd__inv_2
X_22235_ _08592_ VGND VGND VPWR VPWR _09401_ sky130_fd_sc_hd__clkbuf_8
X_29831_ net209 _01566_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[1\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_22166_ _09354_ VGND VGND VPWR VPWR _01101_ sky130_fd_sc_hd__clkbuf_1
X_21117_ _06732_ _08400_ _08405_ _08124_ VGND VGND VPWR VPWR _08406_ sky130_fd_sc_hd__a22o_1
XFILLER_0_218_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29762_ net1108 _01497_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[21\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_26974_ _11803_ _11866_ VGND VGND VPWR VPWR _11871_ sky130_fd_sc_hd__and2_1
X_22097_ rvcpu.dp.plem.WriteDataM\[26\] _09221_ _09295_ rvcpu.dp.plem.WriteDataM\[10\]
+ _09308_ VGND VGND VPWR VPWR _09309_ sky130_fd_sc_hd__a221o_4
XFILLER_0_22_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28713_ _12855_ VGND VGND VPWR VPWR _04147_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_54_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25925_ net2375 _11275_ _11273_ _11282_ VGND VGND VPWR VPWR _02932_ sky130_fd_sc_hd__o211a_1
X_21048_ _07866_ _08335_ _08336_ _07862_ VGND VGND VPWR VPWR _08337_ sky130_fd_sc_hd__o22a_1
XFILLER_0_22_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29693_ net1039 _01428_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[23\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_227_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28644_ _12743_ net4270 net71 VGND VGND VPWR VPWR _12819_ sky130_fd_sc_hd__mux2_1
X_25856_ rvcpu.dp.plfd.PCPlus4D\[27\] _11236_ _08598_ VGND VGND VPWR VPWR _11237_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24807_ _10448_ net3947 _10612_ VGND VGND VPWR VPWR _10617_ sky130_fd_sc_hd__mux2_1
X_28575_ _12760_ net2990 _12777_ VGND VGND VPWR VPWR _12782_ sky130_fd_sc_hd__mux2_1
X_25787_ rvcpu.dp.pcreg.q\[13\] _11178_ VGND VGND VPWR VPWR _11182_ sky130_fd_sc_hd__and2_1
XFILLER_0_201_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22999_ clknet_1_1__leaf__10080_ VGND VGND VPWR VPWR _10085_ sky130_fd_sc_hd__buf_1
XFILLER_0_96_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24154__657 clknet_1_0__leaf__10263_ VGND VGND VPWR VPWR net783 sky130_fd_sc_hd__inv_2
XFILLER_0_9_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15540_ _13403_ _13689_ _13747_ VGND VGND VPWR VPWR _14066_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_57_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27526_ _12093_ net1993 _12188_ VGND VGND VPWR VPWR _12195_ sky130_fd_sc_hd__mux2_1
X_24738_ _10452_ net2100 _10571_ VGND VGND VPWR VPWR _10578_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15471_ _13997_ _13998_ _14000_ _13469_ VGND VGND VPWR VPWR _14001_ sky130_fd_sc_hd__a31o_1
XFILLER_0_166_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24669_ _10538_ net1355 _10531_ _10540_ VGND VGND VPWR VPWR _02418_ sky130_fd_sc_hd__a31o_1
X_27457_ _09290_ VGND VGND VPWR VPWR _12157_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_127_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17210_ _14197_ _04755_ VGND VGND VPWR VPWR _04864_ sky130_fd_sc_hd__nand2_2
X_26408_ _11524_ rvcpu.ALUResultE\[9\] VGND VGND VPWR VPWR _11549_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18190_ _05525_ _05550_ _05553_ _05554_ VGND VGND VPWR VPWR _05555_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_154_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27388_ _12113_ VGND VGND VPWR VPWR _03564_ sky130_fd_sc_hd__clkbuf_1
X_23301__943 clknet_1_1__leaf__10132_ VGND VGND VPWR VPWR net1069 sky130_fd_sc_hd__inv_2
X_29127_ _13079_ VGND VGND VPWR VPWR _04337_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17141_ _04827_ VGND VGND VPWR VPWR _01468_ sky130_fd_sc_hd__clkbuf_1
X_26339_ _11091_ _11497_ VGND VGND VPWR VPWR _11505_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17072_ net3986 _14486_ _04756_ VGND VGND VPWR VPWR _04791_ sky130_fd_sc_hd__mux2_1
X_29058_ _09275_ net3761 net65 VGND VGND VPWR VPWR _13043_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28009_ _12466_ VGND VGND VPWR VPWR _03832_ sky130_fd_sc_hd__clkbuf_1
X_16023_ _14351_ VGND VGND VPWR VPWR _02010_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31020_ clknet_leaf_153_clk _02755_ VGND VGND VPWR VPWR datamem.data_ram\[42\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_208_5490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17974_ _05342_ _05343_ VGND VGND VPWR VPWR _05345_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19713_ datamem.data_ram\[30\]\[0\] _06978_ _06976_ datamem.data_ram\[28\]\[0\] VGND
+ VGND VPWR VPWR _07009_ sky130_fd_sc_hd__a22o_1
X_16925_ net2040 _14476_ _04706_ VGND VGND VPWR VPWR _04713_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_204_5387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32971_ clknet_leaf_145_clk _04393_ VGND VGND VPWR VPWR datamem.data_ram\[63\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_204_5398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_108_Left_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_174_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19644_ _06928_ VGND VGND VPWR VPWR _06940_ sky130_fd_sc_hd__buf_6
X_31922_ _04434_ net118 VGND VGND VPWR VPWR datamem.rd_data_mem\[27\] sky130_fd_sc_hd__dlxtn_1
X_16856_ _04676_ VGND VGND VPWR VPWR _01610_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_205_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_196_5188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15807_ _14233_ VGND VGND VPWR VPWR _02124_ sky130_fd_sc_hd__clkbuf_1
X_31853_ clknet_leaf_124_clk _03307_ VGND VGND VPWR VPWR datamem.data_ram\[61\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_217_5704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_196_5199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19575_ datamem.data_ram\[12\]\[8\] _06686_ _06656_ datamem.data_ram\[9\]\[8\] VGND
+ VGND VPWR VPWR _06871_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_217_5715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16787_ net3174 _14474_ _04634_ VGND VGND VPWR VPWR _04640_ sky130_fd_sc_hd__mux2_1
XFILLER_0_204_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_204_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18526_ _05378_ _05400_ _05886_ VGND VGND VPWR VPWR _05887_ sky130_fd_sc_hd__a21oi_1
X_30804_ clknet_leaf_200_clk _02539_ VGND VGND VPWR VPWR datamem.data_ram\[45\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15738_ _14196_ VGND VGND VPWR VPWR _02156_ sky130_fd_sc_hd__clkbuf_1
X_31784_ clknet_leaf_104_clk _03238_ VGND VGND VPWR VPWR datamem.data_ram\[8\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_887 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18457_ _05274_ _05733_ _05819_ VGND VGND VPWR VPWR _05820_ sky130_fd_sc_hd__and3_2
XFILLER_0_146_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30735_ clknet_leaf_203_clk _02470_ VGND VGND VPWR VPWR datamem.data_ram\[47\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15669_ _14149_ net4141 _14131_ VGND VGND VPWR VPWR _14150_ sky130_fd_sc_hd__mux2_1
XANTENNA_190 _09226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17408_ _04969_ VGND VGND VPWR VPWR _01335_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_172_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23773__361 clknet_1_0__leaf__10202_ VGND VGND VPWR VPWR net487 sky130_fd_sc_hd__inv_2
XFILLER_0_44_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30666_ clknet_leaf_139_clk _02401_ VGND VGND VPWR VPWR datamem.data_ram\[50\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18388_ _05456_ _05463_ _05469_ _05475_ _05683_ _05688_ VGND VGND VPWR VPWR _05752_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_56_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_117_Left_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32405_ clknet_leaf_249_clk _03827_ VGND VGND VPWR VPWR datamem.data_ram\[29\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_209_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17339_ rvcpu.dp.rf.reg_file_arr\[24\]\[3\] _13268_ _04924_ VGND VGND VPWR VPWR _04933_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30597_ clknet_leaf_217_clk _02332_ VGND VGND VPWR VPWR datamem.data_ram\[53\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_20350_ datamem.data_ram\[55\]\[4\] _06993_ _07640_ _07641_ VGND VGND VPWR VPWR _07642_
+ sky130_fd_sc_hd__a211o_1
Xclkload110 clknet_leaf_60_clk VGND VGND VPWR VPWR clkload110/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_153_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32336_ clknet_leaf_275_clk _03758_ VGND VGND VPWR VPWR datamem.data_ram\[31\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload121 clknet_leaf_106_clk VGND VGND VPWR VPWR clkload121/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_4523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload132 clknet_leaf_286_clk VGND VGND VPWR VPWR clkload132/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_109_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_168_4534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload143 clknet_leaf_248_clk VGND VGND VPWR VPWR clkload143/Y sky130_fd_sc_hd__clkinv_4
X_19009_ _06335_ _05728_ _06137_ _06342_ VGND VGND VPWR VPWR _06343_ sky130_fd_sc_hd__a211o_1
Xclkload154 clknet_leaf_277_clk VGND VGND VPWR VPWR clkload154/Y sky130_fd_sc_hd__inv_6
XFILLER_0_140_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20281_ _06916_ _07562_ _07573_ _06713_ VGND VGND VPWR VPWR _07574_ sky130_fd_sc_hd__o211a_1
Xclkload165 clknet_leaf_266_clk VGND VGND VPWR VPWR clkload165/Y sky130_fd_sc_hd__clkinvlp_4
X_32267_ clknet_leaf_210_clk _03689_ VGND VGND VPWR VPWR datamem.data_ram\[33\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload176 clknet_leaf_231_clk VGND VGND VPWR VPWR clkload176/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_45_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload187 clknet_leaf_221_clk VGND VGND VPWR VPWR clkload187/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_178_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22020_ rvcpu.dp.plem.WriteDataM\[20\] _09221_ VGND VGND VPWR VPWR _09246_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload198 clknet_leaf_188_clk VGND VGND VPWR VPWR clkload198/Y sky130_fd_sc_hd__clkinv_4
X_31218_ clknet_leaf_37_clk _02921_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCD\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_228_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3303 rvcpu.dp.pcreg.q\[14\] VGND VGND VPWR VPWR net4453 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32198_ clknet_leaf_229_clk _03620_ VGND VGND VPWR VPWR datamem.data_ram\[36\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_90_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_227_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31149_ clknet_leaf_67_clk rvcpu.ALUResultE\[8\] VGND VGND VPWR VPWR rvcpu.dp.plem.ALUResultM\[8\]
+ sky130_fd_sc_hd__dfxtp_2
Xhold2602 datamem.data_ram\[60\]\[17\] VGND VGND VPWR VPWR net3752 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2613 datamem.data_ram\[51\]\[9\] VGND VGND VPWR VPWR net3763 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2624 datamem.data_ram\[16\]\[24\] VGND VGND VPWR VPWR net3774 sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 rvcpu.dp.plem.lAuiPCM\[21\] VGND VGND VPWR VPWR net1166 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2635 datamem.data_ram\[29\]\[20\] VGND VGND VPWR VPWR net3785 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_126_Left_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_89_Right_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold27 rvcpu.dp.plem.PCPlus4M\[29\] VGND VGND VPWR VPWR net1177 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_127_3541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1901 rvcpu.dp.rf.reg_file_arr\[11\]\[15\] VGND VGND VPWR VPWR net3051 sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 rvcpu.dp.plde.PCPlus4E\[7\] VGND VGND VPWR VPWR net1188 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_127_3552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2646 datamem.data_ram\[14\]\[27\] VGND VGND VPWR VPWR net3796 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 rvcpu.dp.plde.PCPlus4E\[23\] VGND VGND VPWR VPWR net1199 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1912 datamem.data_ram\[41\]\[18\] VGND VGND VPWR VPWR net3062 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2657 datamem.data_ram\[27\]\[10\] VGND VGND VPWR VPWR net3807 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2668 rvcpu.dp.rf.reg_file_arr\[20\]\[26\] VGND VGND VPWR VPWR net3818 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1923 datamem.data_ram\[50\]\[25\] VGND VGND VPWR VPWR net3073 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1934 datamem.data_ram\[24\]\[16\] VGND VGND VPWR VPWR net3084 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2679 datamem.data_ram\[10\]\[9\] VGND VGND VPWR VPWR net3829 sky130_fd_sc_hd__dlygate4sd3_1
X_22922_ _06587_ VGND VGND VPWR VPWR _10055_ sky130_fd_sc_hd__buf_2
Xhold1945 rvcpu.dp.rf.reg_file_arr\[12\]\[22\] VGND VGND VPWR VPWR net3095 sky130_fd_sc_hd__dlygate4sd3_1
X_25710_ _11128_ VGND VGND VPWR VPWR _02871_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_67_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26690_ _11645_ _11694_ VGND VGND VPWR VPWR _11699_ sky130_fd_sc_hd__and2_1
Xhold1956 datamem.data_ram\[1\]\[29\] VGND VGND VPWR VPWR net3106 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_123_3438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_123_3449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1967 datamem.data_ram\[42\]\[29\] VGND VGND VPWR VPWR net3117 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1978 rvcpu.dp.rf.reg_file_arr\[28\]\[15\] VGND VGND VPWR VPWR net3128 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1989 datamem.data_ram\[27\]\[31\] VGND VGND VPWR VPWR net3139 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25641_ _11089_ _11079_ VGND VGND VPWR VPWR _11090_ sky130_fd_sc_hd__and2_1
X_22853_ _09398_ _09989_ VGND VGND VPWR VPWR _09990_ sky130_fd_sc_hd__or2_1
XFILLER_0_155_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21804_ rvcpu.dp.rf.reg_file_arr\[24\]\[22\] rvcpu.dp.rf.reg_file_arr\[25\]\[22\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[22\] rvcpu.dp.rf.reg_file_arr\[27\]\[22\] rvcpu.dp.plfd.InstrD\[15\]
+ _08526_ VGND VGND VPWR VPWR _09044_ sky130_fd_sc_hd__mux4_1
XFILLER_0_211_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25572_ _11018_ net1405 _11041_ _11046_ VGND VGND VPWR VPWR _02815_ sky130_fd_sc_hd__a31o_1
X_28360_ _12456_ net2545 net95 VGND VGND VPWR VPWR _12655_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22784_ _09495_ _09924_ _09472_ VGND VGND VPWR VPWR _09925_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27311_ _12061_ net1617 _12065_ _12070_ VGND VGND VPWR VPWR _03530_ sky130_fd_sc_hd__a31o_1
X_24523_ _10385_ datamem.data_ram\[52\]\[8\] _10456_ VGND VGND VPWR VPWR _10457_ sky130_fd_sc_hd__mux2_1
XFILLER_0_213_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21735_ rvcpu.dp.rf.reg_file_arr\[8\]\[18\] rvcpu.dp.rf.reg_file_arr\[10\]\[18\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[18\] rvcpu.dp.rf.reg_file_arr\[11\]\[18\] _08560_
+ _08561_ VGND VGND VPWR VPWR _08979_ sky130_fd_sc_hd__mux4_1
XFILLER_0_52_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28291_ _12439_ net4156 _12613_ VGND VGND VPWR VPWR _12618_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_26_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_135_Left_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_98_Right_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24454_ _10412_ net1916 _10404_ _10415_ VGND VGND VPWR VPWR _02328_ sky130_fd_sc_hd__a31o_1
X_27242_ _12022_ net1630 _12030_ _12034_ VGND VGND VPWR VPWR _03497_ sky130_fd_sc_hd__a31o_1
XFILLER_0_108_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21666_ _08695_ _08913_ VGND VGND VPWR VPWR _08914_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27173_ _11980_ _11984_ VGND VGND VPWR VPWR _11993_ sky130_fd_sc_hd__and2_1
XFILLER_0_117_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20617_ datamem.data_ram\[30\]\[13\] _07085_ _06633_ datamem.data_ram\[27\]\[13\]
+ _07907_ VGND VGND VPWR VPWR _07908_ sky130_fd_sc_hd__o221a_1
X_24385_ _10371_ VGND VGND VPWR VPWR _02303_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21597_ rvcpu.dp.rf.reg_file_arr\[20\]\[11\] rvcpu.dp.rf.reg_file_arr\[21\]\[11\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[11\] rvcpu.dp.rf.reg_file_arr\[23\]\[11\] _08799_
+ _08800_ VGND VGND VPWR VPWR _08848_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_10_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26124_ net1775 _11397_ VGND VGND VPWR VPWR _11398_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_10_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23336_ clknet_1_1__leaf__10130_ VGND VGND VPWR VPWR _10136_ sky130_fd_sc_hd__buf_1
X_20548_ _07838_ VGND VGND VPWR VPWR _07839_ sky130_fd_sc_hd__buf_6
XFILLER_0_85_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26055_ _11353_ net1842 _11350_ _11356_ VGND VGND VPWR VPWR _02988_ sky130_fd_sc_hd__a31o_1
XFILLER_0_21_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20479_ datamem.data_ram\[50\]\[20\] _06609_ _06632_ datamem.data_ram\[51\]\[20\]
+ _06677_ VGND VGND VPWR VPWR _07771_ sky130_fd_sc_hd__o221a_1
X_25006_ _09266_ VGND VGND VPWR VPWR _10724_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_56_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22218_ _08592_ VGND VGND VPWR VPWR _09384_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_56_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23198_ _09248_ net4302 _10115_ VGND VGND VPWR VPWR _10120_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_144_Left_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29814_ net192 _01549_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[1\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_22149_ _09344_ VGND VGND VPWR VPWR _01094_ sky130_fd_sc_hd__clkbuf_1
X_29745_ net1091 _01480_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[21\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26957_ _11849_ net1538 _11853_ _11860_ VGND VGND VPWR VPWR _03386_ sky130_fd_sc_hd__a31o_1
X_14971_ _13518_ _13519_ _13442_ VGND VGND VPWR VPWR _13520_ sky130_fd_sc_hd__a21o_1
X_23943__497 clknet_1_0__leaf__10228_ VGND VGND VPWR VPWR net623 sky130_fd_sc_hd__inv_2
XFILLER_0_22_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16710_ _04599_ VGND VGND VPWR VPWR _01687_ sky130_fd_sc_hd__clkbuf_1
X_25908_ net1657 _11256_ _11258_ _11272_ VGND VGND VPWR VPWR _02925_ sky130_fd_sc_hd__o211a_1
X_17690_ _05119_ VGND VGND VPWR VPWR _01195_ sky130_fd_sc_hd__clkbuf_1
X_29676_ net1022 _01411_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[23\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_26888_ _11813_ net1439 _11809_ _11816_ VGND VGND VPWR VPWR _03361_ sky130_fd_sc_hd__a31o_1
XFILLER_0_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28627_ _12760_ net3472 _12805_ VGND VGND VPWR VPWR _12810_ sky130_fd_sc_hd__mux2_1
X_16641_ _14172_ net4403 _04562_ VGND VGND VPWR VPWR _04563_ sky130_fd_sc_hd__mux2_1
X_25839_ _11221_ _11222_ VGND VGND VPWR VPWR _11223_ sky130_fd_sc_hd__nor2_1
XFILLER_0_199_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26498__51 clknet_1_0__leaf__11601_ VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__inv_2
XFILLER_0_214_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19360_ _06655_ VGND VGND VPWR VPWR _06656_ sky130_fd_sc_hd__buf_4
X_16572_ _14172_ net4434 _04525_ VGND VGND VPWR VPWR _04526_ sky130_fd_sc_hd__mux2_1
X_28558_ _12696_ net3845 _12768_ VGND VGND VPWR VPWR _12773_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_201_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_153_Left_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18311_ _05675_ VGND VGND VPWR VPWR _05676_ sky130_fd_sc_hd__clkbuf_4
X_15523_ _13599_ _14048_ _14049_ VGND VGND VPWR VPWR _14050_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_191_5074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27509_ _12155_ net3610 _12179_ VGND VGND VPWR VPWR _12186_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_191_5085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19291_ _06585_ VGND VGND VPWR VPWR _06587_ sky130_fd_sc_hd__buf_4
XFILLER_0_167_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28489_ _11972_ _12724_ VGND VGND VPWR VPWR _12729_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18242_ _05606_ _05415_ VGND VGND VPWR VPWR _05607_ sky130_fd_sc_hd__or2_1
X_30520_ clknet_leaf_144_clk _02255_ VGND VGND VPWR VPWR datamem.data_ram\[56\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_15454_ _13706_ _13980_ _13983_ _13664_ VGND VGND VPWR VPWR _13984_ sky130_fd_sc_hd__o211a_1
XFILLER_0_182_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18173_ rvcpu.dp.plem.ALUResultM\[27\] _05293_ _05294_ _13194_ VGND VGND VPWR VPWR
+ _05538_ sky130_fd_sc_hd__o22a_1
X_30451_ net789 _02186_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[29\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_15385_ _13528_ _13634_ _13646_ VGND VGND VPWR VPWR _13918_ sky130_fd_sc_hd__o21a_1
XFILLER_0_167_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_182_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17124_ _14179_ net3896 _04815_ VGND VGND VPWR VPWR _04819_ sky130_fd_sc_hd__mux2_1
X_23536__163 clknet_1_0__leaf__10171_ VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__inv_2
XFILLER_0_52_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30382_ clknet_leaf_176_clk _02117_ VGND VGND VPWR VPWR datamem.data_ram\[58\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_150_4092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold508 datamem.data_ram\[27\]\[2\] VGND VGND VPWR VPWR net1658 sky130_fd_sc_hd__dlygate4sd3_1
X_32121_ clknet_leaf_227_clk _03543_ VGND VGND VPWR VPWR datamem.data_ram\[7\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold519 _02936_ VGND VGND VPWR VPWR net1669 sky130_fd_sc_hd__dlygate4sd3_1
X_17055_ _04782_ VGND VGND VPWR VPWR _01509_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_162_Left_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16006_ net2775 _13266_ _14333_ VGND VGND VPWR VPWR _14341_ sky130_fd_sc_hd__mux2_1
X_32052_ clknet_leaf_126_clk _03474_ VGND VGND VPWR VPWR datamem.data_ram\[30\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_206_5438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_206_5449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31003_ clknet_leaf_99_clk _02738_ VGND VGND VPWR VPWR datamem.data_ram\[22\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_209_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_198_5239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17957_ rvcpu.dp.plem.ALUResultM\[12\] _05328_ _05175_ VGND VGND VPWR VPWR _05329_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1208 rvcpu.dp.rf.reg_file_arr\[2\]\[20\] VGND VGND VPWR VPWR net2358 sky130_fd_sc_hd__dlygate4sd3_1
X_24022__554 clknet_1_0__leaf__10242_ VGND VGND VPWR VPWR net680 sky130_fd_sc_hd__inv_2
Xhold1219 datamem.data_ram\[1\]\[18\] VGND VGND VPWR VPWR net2369 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16908_ net2075 _14459_ _04695_ VGND VGND VPWR VPWR _04704_ sky130_fd_sc_hd__mux2_1
X_32954_ clknet_leaf_97_clk _04376_ VGND VGND VPWR VPWR datamem.data_ram\[6\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_17888_ rvcpu.dp.plde.Rs1E\[0\] rvcpu.dp.plmw.RdW\[0\] VGND VGND VPWR VPWR _05261_
+ sky130_fd_sc_hd__or2b_1
XFILLER_0_206_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19627_ _06605_ _06922_ VGND VGND VPWR VPWR _06923_ sky130_fd_sc_hd__nor2_1
X_31905_ _04416_ net120 VGND VGND VPWR VPWR datamem.rd_data_mem\[10\] sky130_fd_sc_hd__dlxtn_1
XFILLER_0_219_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16839_ _04667_ VGND VGND VPWR VPWR _01618_ sky130_fd_sc_hd__clkbuf_1
X_32885_ clknet_leaf_286_clk _04307_ VGND VGND VPWR VPWR datamem.data_ram\[10\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23308__949 clknet_1_0__leaf__10133_ VGND VGND VPWR VPWR net1075 sky130_fd_sc_hd__inv_2
XFILLER_0_75_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19558_ datamem.data_ram\[6\]\[24\] _06718_ _06686_ datamem.data_ram\[4\]\[24\] VGND
+ VGND VPWR VPWR _06854_ sky130_fd_sc_hd__o22a_1
X_31836_ clknet_leaf_213_clk _03290_ VGND VGND VPWR VPWR datamem.data_ram\[3\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_211_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_157_4257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_4268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18509_ _05394_ _05826_ _05870_ _05668_ VGND VGND VPWR VPWR _05871_ sky130_fd_sc_hd__o22a_1
XFILLER_0_146_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19489_ datamem.data_ram\[18\]\[16\] _06611_ _06784_ datamem.data_ram\[23\]\[16\]
+ VGND VGND VPWR VPWR _06785_ sky130_fd_sc_hd__o22a_1
X_23697__292 clknet_1_0__leaf__10195_ VGND VGND VPWR VPWR net418 sky130_fd_sc_hd__inv_2
X_31767_ clknet_leaf_228_clk _03221_ VGND VGND VPWR VPWR datamem.data_ram\[1\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_186_892 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21520_ _08572_ _08774_ VGND VGND VPWR VPWR _08775_ sky130_fd_sc_hd__or2_1
X_30718_ clknet_leaf_178_clk _02453_ VGND VGND VPWR VPWR datamem.data_ram\[49\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31698_ clknet_leaf_42_clk _03156_ VGND VGND VPWR VPWR rvcpu.dp.pcreg.q\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21451_ rvcpu.dp.rf.reg_file_arr\[24\]\[4\] rvcpu.dp.rf.reg_file_arr\[25\]\[4\] rvcpu.dp.rf.reg_file_arr\[26\]\[4\]
+ rvcpu.dp.rf.reg_file_arr\[27\]\[4\] _08517_ _08519_ VGND VGND VPWR VPWR _08709_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_21_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30649_ clknet_leaf_178_clk _02384_ VGND VGND VPWR VPWR datamem.data_ram\[51\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20402_ datamem.data_ram\[34\]\[12\] _06691_ _06778_ datamem.data_ram\[32\]\[12\]
+ _07693_ VGND VGND VPWR VPWR _07694_ sky130_fd_sc_hd__o221a_1
XFILLER_0_189_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_3275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21382_ _08511_ _08642_ VGND VGND VPWR VPWR _08643_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_116_3286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20333_ datamem.data_ram\[43\]\[4\] _06966_ _06977_ datamem.data_ram\[44\]\[4\] _07624_
+ VGND VGND VPWR VPWR _07625_ sky130_fd_sc_hd__a221o_1
XFILLER_0_31_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32319_ clknet_leaf_186_clk _03741_ VGND VGND VPWR VPWR datamem.data_ram\[31\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_187_4976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_187_4987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput17 net17 VGND VGND VPWR VPWR Instr[23] sky130_fd_sc_hd__buf_2
Xoutput28 net28 VGND VGND VPWR VPWR Instr[4] sky130_fd_sc_hd__buf_2
XFILLER_0_222_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20264_ datamem.data_ram\[63\]\[19\] _06760_ _06766_ datamem.data_ram\[60\]\[19\]
+ VGND VGND VPWR VPWR _07557_ sky130_fd_sc_hd__o22a_1
XFILLER_0_113_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_129_3603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold3100 datamem.data_ram\[13\]\[14\] VGND VGND VPWR VPWR net4250 sky130_fd_sc_hd__dlygate4sd3_1
X_22003_ _09224_ net4405 _09232_ VGND VGND VPWR VPWR _09233_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3111 datamem.data_ram\[12\]\[14\] VGND VGND VPWR VPWR net4261 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3122 rvcpu.dp.plem.ALUResultM\[3\] VGND VGND VPWR VPWR net4272 sky130_fd_sc_hd__dlygate4sd3_1
X_27860_ _12378_ VGND VGND VPWR VPWR _03771_ sky130_fd_sc_hd__clkbuf_1
Xhold3133 rvcpu.dp.rf.reg_file_arr\[26\]\[22\] VGND VGND VPWR VPWR net4283 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold3144 datamem.data_ram\[28\]\[16\] VGND VGND VPWR VPWR net4294 sky130_fd_sc_hd__dlygate4sd3_1
X_20195_ datamem.data_ram\[38\]\[11\] _06764_ _07024_ datamem.data_ram\[36\]\[11\]
+ VGND VGND VPWR VPWR _07488_ sky130_fd_sc_hd__o22a_1
Xhold2410 datamem.data_ram\[9\]\[9\] VGND VGND VPWR VPWR net3560 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3155 rvcpu.dp.rf.reg_file_arr\[15\]\[14\] VGND VGND VPWR VPWR net4305 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26811_ _11689_ _11762_ VGND VGND VPWR VPWR _11770_ sky130_fd_sc_hd__and2_1
Xhold3166 rvcpu.dp.plem.ALUResultM\[30\] VGND VGND VPWR VPWR net4316 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2421 datamem.data_ram\[19\]\[15\] VGND VGND VPWR VPWR net3571 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3177 datamem.data_ram\[55\]\[22\] VGND VGND VPWR VPWR net4327 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2432 rvcpu.dp.rf.reg_file_arr\[25\]\[11\] VGND VGND VPWR VPWR net3582 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2443 datamem.data_ram\[10\]\[16\] VGND VGND VPWR VPWR net3593 sky130_fd_sc_hd__dlygate4sd3_1
X_27791_ _12337_ VGND VGND VPWR VPWR _03743_ sky130_fd_sc_hd__clkbuf_1
Xhold3188 rvcpu.dp.rf.reg_file_arr\[24\]\[4\] VGND VGND VPWR VPWR net4338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2454 rvcpu.dp.rf.reg_file_arr\[29\]\[0\] VGND VGND VPWR VPWR net3604 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3199 rvcpu.dp.plfd.InstrD\[6\] VGND VGND VPWR VPWR net4349 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1720 datamem.data_ram\[63\]\[19\] VGND VGND VPWR VPWR net2870 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_3994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2465 rvcpu.dp.rf.reg_file_arr\[2\]\[21\] VGND VGND VPWR VPWR net3615 sky130_fd_sc_hd__dlygate4sd3_1
X_29530_ clknet_leaf_180_clk _01265_ VGND VGND VPWR VPWR datamem.data_ram\[5\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_26742_ _11681_ _11726_ VGND VGND VPWR VPWR _11729_ sky130_fd_sc_hd__and2_1
Xhold2476 rvcpu.dp.rf.reg_file_arr\[20\]\[16\] VGND VGND VPWR VPWR net3626 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1731 rvcpu.dp.rf.reg_file_arr\[0\]\[18\] VGND VGND VPWR VPWR net2881 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1742 datamem.data_ram\[14\]\[17\] VGND VGND VPWR VPWR net2892 sky130_fd_sc_hd__dlygate4sd3_1
X_23954_ _09236_ net4353 _10229_ VGND VGND VPWR VPWR _10231_ sky130_fd_sc_hd__mux2_1
Xhold2487 datamem.data_ram\[60\]\[13\] VGND VGND VPWR VPWR net3637 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1753 rvcpu.dp.rf.reg_file_arr\[1\]\[16\] VGND VGND VPWR VPWR net2903 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2498 datamem.data_ram\[7\]\[13\] VGND VGND VPWR VPWR net3648 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1764 rvcpu.dp.rf.reg_file_arr\[27\]\[18\] VGND VGND VPWR VPWR net2914 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1775 datamem.data_ram\[15\]\[30\] VGND VGND VPWR VPWR net2925 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22905_ _09388_ _10031_ _10035_ _10039_ VGND VGND VPWR VPWR _10040_ sky130_fd_sc_hd__and4_1
Xclkbuf_1_1__f__10242_ clknet_0__10242_ VGND VGND VPWR VPWR clknet_1_1__leaf__10242_
+ sky130_fd_sc_hd__clkbuf_16
X_29461_ net823 _01196_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[2\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_26673_ _11683_ net1757 _11675_ _11688_ VGND VGND VPWR VPWR _03274_ sky130_fd_sc_hd__a31o_1
Xhold1786 datamem.data_ram\[36\]\[9\] VGND VGND VPWR VPWR net2936 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1797 rvcpu.dp.rf.reg_file_arr\[9\]\[16\] VGND VGND VPWR VPWR net2947 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28412_ _12456_ net2842 _12678_ VGND VGND VPWR VPWR _12683_ sky130_fd_sc_hd__mux2_1
X_25624_ _10047_ VGND VGND VPWR VPWR _11078_ sky130_fd_sc_hd__clkbuf_4
X_22836_ _09422_ _09973_ VGND VGND VPWR VPWR _09974_ sky130_fd_sc_hd__nor2_1
X_29392_ clknet_leaf_1_clk _01127_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD2E\[3\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__10173_ clknet_0__10173_ VGND VGND VPWR VPWR clknet_1_1__leaf__10173_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_6_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28343_ _12439_ net3499 _12641_ VGND VGND VPWR VPWR _12646_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25555_ _10762_ net2828 _11030_ VGND VGND VPWR VPWR _11036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22767_ _09903_ _09905_ _09908_ _09412_ _09525_ VGND VGND VPWR VPWR _09909_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24506_ _10445_ VGND VGND VPWR VPWR _02350_ sky130_fd_sc_hd__clkbuf_1
X_21718_ _08835_ _08962_ VGND VGND VPWR VPWR _08963_ sky130_fd_sc_hd__or2_1
X_25486_ _10783_ net35 _10996_ net1301 VGND VGND VPWR VPWR _02779_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_45_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28274_ _12608_ VGND VGND VPWR VPWR _03955_ sky130_fd_sc_hd__clkbuf_1
X_22698_ _09622_ _09841_ _09843_ VGND VGND VPWR VPWR _09844_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_117_Right_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27225_ _12022_ net1587 _12018_ _12024_ VGND VGND VPWR VPWR _03490_ sky130_fd_sc_hd__a31o_1
XFILLER_0_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24437_ _07019_ _10402_ _10044_ VGND VGND VPWR VPWR _10403_ sky130_fd_sc_hd__or3_1
XFILLER_0_137_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21649_ _08817_ _08895_ _08897_ _08700_ VGND VGND VPWR VPWR _08898_ sky130_fd_sc_hd__a211o_1
XFILLER_0_118_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15170_ _13688_ _13702_ _13713_ VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__a21oi_4
XFILLER_0_151_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27156_ _11982_ VGND VGND VPWR VPWR _11983_ sky130_fd_sc_hd__buf_2
XFILLER_0_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24368_ _09318_ net3847 net61 VGND VGND VPWR VPWR _10362_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_90 _06797_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26107_ net1455 _11386_ VGND VGND VPWR VPWR _11389_ sky130_fd_sc_hd__and2_1
XFILLER_0_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27087_ _11918_ VGND VGND VPWR VPWR _11938_ sky130_fd_sc_hd__buf_2
XFILLER_0_205_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24299_ _09288_ net3842 _10316_ VGND VGND VPWR VPWR _10323_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26038_ _11089_ _11340_ VGND VGND VPWR VPWR _11346_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18860_ _05781_ _06079_ _06203_ _05660_ VGND VGND VPWR VPWR _06204_ sky130_fd_sc_hd__a211o_1
XFILLER_0_24_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17811_ rvcpu.dp.plem.ALUResultM\[29\] _05201_ _05178_ VGND VGND VPWR VPWR _05202_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_206_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_201_5313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18791_ _06031_ _06138_ _05819_ VGND VGND VPWR VPWR _06139_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_201_5324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27989_ _12453_ VGND VGND VPWR VPWR _03825_ sky130_fd_sc_hd__clkbuf_1
X_23566__189 clknet_1_0__leaf__10175_ VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__inv_2
X_29728_ net1074 _01463_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[22\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_17742_ _05146_ VGND VGND VPWR VPWR _01170_ sky130_fd_sc_hd__clkbuf_1
X_14954_ _13331_ _13458_ VGND VGND VPWR VPWR _13503_ sky130_fd_sc_hd__nor2_1
XFILLER_0_215_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_199_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_193_5125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29659_ net1005 _01394_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[24\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_17673_ net4205 _13259_ _05104_ VGND VGND VPWR VPWR _05110_ sky130_fd_sc_hd__mux2_1
X_14885_ _13423_ _13427_ _13429_ _13436_ VGND VGND VPWR VPWR _13437_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_193_5136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_195_clk clknet_5_29__leaf_clk VGND VGND VPWR VPWR clknet_leaf_195_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_202_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19412_ datamem.data_ram\[5\]\[16\] _06703_ _06707_ datamem.data_ram\[7\]\[16\] VGND
+ VGND VPWR VPWR _06708_ sky130_fd_sc_hd__o22a_1
X_16624_ _14156_ net2069 _04551_ VGND VGND VPWR VPWR _04554_ sky130_fd_sc_hd__mux2_1
X_32670_ clknet_leaf_284_clk _04092_ VGND VGND VPWR VPWR datamem.data_ram\[19\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
Xmax_cap70 _12896_ VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__buf_4
XFILLER_0_212_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap81 _12233_ VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__buf_4
X_31621_ clknet_leaf_66_clk net1198 VGND VGND VPWR VPWR rvcpu.dp.plmw.lAuiPCW\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_19343_ net122 _06584_ VGND VGND VPWR VPWR _06639_ sky130_fd_sc_hd__nand2_8
Xmax_cap92 _10650_ VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__buf_4
XFILLER_0_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16555_ _14156_ net2484 _04514_ VGND VGND VPWR VPWR _04517_ sky130_fd_sc_hd__mux2_1
XFILLER_0_174_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15506_ _13454_ _13613_ _13597_ VGND VGND VPWR VPWR _14033_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_57_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31552_ clknet_leaf_63_clk datamem.rd_data_mem\[2\] VGND VGND VPWR VPWR rvcpu.dp.plmw.ReadDataW\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_19274_ _06567_ _06569_ _06571_ _06573_ VGND VGND VPWR VPWR _04447_ sky130_fd_sc_hd__a31o_1
XFILLER_0_127_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16486_ _04480_ VGND VGND VPWR VPWR _01800_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_14_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_152_4132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_152_4143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_4154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18225_ _05321_ rvcpu.dp.SrcBFW_Mux.y\[4\] _05362_ VGND VGND VPWR VPWR _05590_ sky130_fd_sc_hd__o21a_4
X_30503_ clknet_leaf_266_clk _02238_ VGND VGND VPWR VPWR datamem.data_ram\[57\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_15437_ _13964_ _13966_ _13967_ _13539_ VGND VGND VPWR VPWR _13968_ sky130_fd_sc_hd__a31o_1
XFILLER_0_143_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31483_ clknet_leaf_65_clk rvcpu.dp.lAuiPCE\[9\] VGND VGND VPWR VPWR rvcpu.dp.plem.lAuiPCM\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_480 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18156_ _05520_ _05479_ _05472_ VGND VGND VPWR VPWR _05521_ sky130_fd_sc_hd__a21o_1
XFILLER_0_41_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30434_ net772 _02169_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[29\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_15368_ _13774_ _13892_ _13895_ _13896_ _13902_ VGND VGND VPWR VPWR _13903_ sky130_fd_sc_hd__a32o_1
Xclkbuf_1_0__f__10262_ clknet_0__10262_ VGND VGND VPWR VPWR clknet_1_0__leaf__10262_
+ sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_170_Left_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17107_ _14162_ net2297 _04804_ VGND VGND VPWR VPWR _04810_ sky130_fd_sc_hd__mux2_1
Xhold305 rvcpu.dp.plfd.PCPlus4D\[10\] VGND VGND VPWR VPWR net1455 sky130_fd_sc_hd__dlygate4sd3_1
Xhold316 datamem.data_ram\[42\]\[4\] VGND VGND VPWR VPWR net1466 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_145_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18087_ rvcpu.dp.plem.ALUResultM\[23\] _05339_ _05340_ _13206_ VGND VGND VPWR VPWR
+ _05455_ sky130_fd_sc_hd__o22a_1
XFILLER_0_29_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30365_ net711 _02100_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[3\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_15299_ _13559_ _13689_ _13639_ VGND VGND VPWR VPWR _13837_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_68_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold327 datamem.data_ram\[56\]\[4\] VGND VGND VPWR VPWR net1477 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__10193_ clknet_0__10193_ VGND VGND VPWR VPWR clknet_1_0__leaf__10193_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_1_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_229_5983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold338 datamem.data_ram\[19\]\[2\] VGND VGND VPWR VPWR net1488 sky130_fd_sc_hd__dlygate4sd3_1
X_32104_ clknet_leaf_114_clk _03526_ VGND VGND VPWR VPWR datamem.data_ram\[23\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_229_5994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold349 datamem.data_ram\[20\]\[2\] VGND VGND VPWR VPWR net1499 sky130_fd_sc_hd__dlygate4sd3_1
X_17038_ _04773_ VGND VGND VPWR VPWR _01517_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_111_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30296_ net642 _02031_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[5\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32035_ clknet_leaf_130_clk _03457_ VGND VGND VPWR VPWR datamem.data_ram\[50\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_182_4862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_4873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18989_ _05305_ _05641_ _06323_ VGND VGND VPWR VPWR _06324_ sky130_fd_sc_hd__a21o_1
X_23052__752 clknet_1_1__leaf__10090_ VGND VGND VPWR VPWR net878 sky130_fd_sc_hd__inv_2
Xhold1005 rvcpu.dp.rf.reg_file_arr\[3\]\[4\] VGND VGND VPWR VPWR net2155 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_175_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1016 rvcpu.dp.rf.reg_file_arr\[7\]\[15\] VGND VGND VPWR VPWR net2166 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1027 datamem.data_ram\[0\]\[31\] VGND VGND VPWR VPWR net2177 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1038 datamem.data_ram\[37\]\[9\] VGND VGND VPWR VPWR net2188 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1049 rvcpu.dp.rf.reg_file_arr\[15\]\[30\] VGND VGND VPWR VPWR net2199 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_219_Right_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_217_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_197_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_159_4308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20951_ _06590_ _08183_ _08240_ _07227_ VGND VGND VPWR VPWR _08241_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_159_4319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32937_ clknet_leaf_156_clk _04359_ VGND VGND VPWR VPWR datamem.data_ram\[6\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_1_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_186_clk clknet_5_22__leaf_clk VGND VGND VPWR VPWR clknet_leaf_186_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_108_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_3880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_3891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20882_ datamem.data_ram\[41\]\[14\] _06658_ _08171_ _07845_ VGND VGND VPWR VPWR
+ _08172_ sky130_fd_sc_hd__o22a_1
X_32868_ clknet_leaf_257_clk _04290_ VGND VGND VPWR VPWR datamem.data_ram\[11\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22621_ _09528_ _09770_ _09426_ VGND VGND VPWR VPWR _09771_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_81_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31819_ clknet_leaf_103_clk _03273_ VGND VGND VPWR VPWR datamem.data_ram\[9\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32799_ clknet_leaf_185_clk _04221_ VGND VGND VPWR VPWR datamem.data_ram\[13\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25340_ _10764_ net2942 _10909_ VGND VGND VPWR VPWR _10916_ sky130_fd_sc_hd__mux2_1
X_22552_ _09388_ VGND VGND VPWR VPWR _09705_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_118_3326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_118_3337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21503_ _08565_ _08756_ _08758_ _08576_ VGND VGND VPWR VPWR _08759_ sky130_fd_sc_hd__o211a_1
X_25271_ _10876_ net1374 _10867_ _10877_ VGND VGND VPWR VPWR _02683_ sky130_fd_sc_hd__a31o_1
XFILLER_0_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22483_ rvcpu.dp.rf.reg_file_arr\[28\]\[9\] rvcpu.dp.rf.reg_file_arr\[30\]\[9\] rvcpu.dp.rf.reg_file_arr\[29\]\[9\]
+ rvcpu.dp.rf.reg_file_arr\[31\]\[9\] _09558_ _09453_ VGND VGND VPWR VPWR _09640_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_1_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27010_ _11889_ net1604 _11885_ _11891_ VGND VGND VPWR VPWR _03408_ sky130_fd_sc_hd__a31o_1
X_24222_ _09240_ net4279 _10279_ VGND VGND VPWR VPWR _10282_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21434_ _08533_ VGND VGND VPWR VPWR _08693_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_40_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21365_ _08557_ VGND VGND VPWR VPWR _08626_ sky130_fd_sc_hd__buf_2
XFILLER_0_86_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_110_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_110_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_47_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20316_ datamem.data_ram\[8\]\[4\] _07138_ _07606_ _07607_ VGND VGND VPWR VPWR _07608_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_124_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28961_ _12987_ VGND VGND VPWR VPWR _12988_ sky130_fd_sc_hd__buf_2
X_24084_ _09282_ net2540 _10249_ VGND VGND VPWR VPWR _10254_ sky130_fd_sc_hd__mux2_1
Xhold850 rvcpu.dp.rf.reg_file_arr\[11\]\[21\] VGND VGND VPWR VPWR net2000 sky130_fd_sc_hd__dlygate4sd3_1
X_21296_ rvcpu.dp.plfd.InstrD\[19\] _08557_ VGND VGND VPWR VPWR _08558_ sky130_fd_sc_hd__nor2_4
Xhold861 datamem.data_ram\[10\]\[15\] VGND VGND VPWR VPWR net2011 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_219_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold872 rvcpu.dp.plfd.PCD\[30\] VGND VGND VPWR VPWR net2022 sky130_fd_sc_hd__dlygate4sd3_1
X_27912_ _12407_ VGND VGND VPWR VPWR _03794_ sky130_fd_sc_hd__clkbuf_1
X_20247_ datamem.data_ram\[34\]\[3\] _06931_ _06924_ datamem.data_ram\[39\]\[3\] VGND
+ VGND VPWR VPWR _07540_ sky130_fd_sc_hd__a22o_1
Xhold883 rvcpu.dp.rf.reg_file_arr\[6\]\[7\] VGND VGND VPWR VPWR net2033 sky130_fd_sc_hd__dlygate4sd3_1
X_28892_ _12734_ net2496 net68 VGND VGND VPWR VPWR _12951_ sky130_fd_sc_hd__mux2_1
Xhold894 rvcpu.dp.rf.reg_file_arr\[7\]\[22\] VGND VGND VPWR VPWR net2044 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27843_ _12368_ VGND VGND VPWR VPWR _03764_ sky130_fd_sc_hd__clkbuf_1
X_23485__132 clknet_1_0__leaf__10159_ VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__inv_2
X_20178_ _06603_ _07463_ _07465_ _07470_ VGND VGND VPWR VPWR _07471_ sky130_fd_sc_hd__a31o_1
Xhold2240 datamem.data_ram\[19\]\[27\] VGND VGND VPWR VPWR net3390 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2251 rvcpu.dp.rf.reg_file_arr\[26\]\[7\] VGND VGND VPWR VPWR net3401 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2262 datamem.data_ram\[27\]\[26\] VGND VGND VPWR VPWR net3412 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_5_5__f_clk clknet_2_0_0_clk VGND VGND VPWR VPWR clknet_5_5__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_27774_ _12083_ net3526 _12326_ VGND VGND VPWR VPWR _12328_ sky130_fd_sc_hd__mux2_1
Xhold2273 rvcpu.dp.rf.reg_file_arr\[25\]\[12\] VGND VGND VPWR VPWR net3423 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24986_ _10713_ VGND VGND VPWR VPWR _02562_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2284 datamem.data_ram\[48\]\[26\] VGND VGND VPWR VPWR net3434 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2295 rvcpu.dp.rf.reg_file_arr\[18\]\[21\] VGND VGND VPWR VPWR net3445 sky130_fd_sc_hd__dlygate4sd3_1
X_29513_ net875 _01248_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[28\]\[20\] sky130_fd_sc_hd__dfxtp_1
Xhold1550 datamem.data_ram\[7\]\[31\] VGND VGND VPWR VPWR net2700 sky130_fd_sc_hd__dlygate4sd3_1
X_26725_ _11718_ VGND VGND VPWR VPWR _03296_ sky130_fd_sc_hd__clkbuf_1
Xhold1561 rvcpu.dp.rf.reg_file_arr\[30\]\[10\] VGND VGND VPWR VPWR net2711 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1572 datamem.data_ram\[38\]\[17\] VGND VGND VPWR VPWR net2722 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_177_clk clknet_5_25__leaf_clk VGND VGND VPWR VPWR clknet_leaf_177_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_19_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1583 rvcpu.dp.rf.reg_file_arr\[27\]\[10\] VGND VGND VPWR VPWR net2733 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1594 rvcpu.dp.rf.reg_file_arr\[22\]\[8\] VGND VGND VPWR VPWR net2744 sky130_fd_sc_hd__dlygate4sd3_1
X_29444_ net806 _01179_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[30\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__10225_ clknet_0__10225_ VGND VGND VPWR VPWR clknet_1_1__leaf__10225_
+ sky130_fd_sc_hd__clkbuf_16
X_26656_ _10268_ _10935_ _11609_ VGND VGND VPWR VPWR _11677_ sky130_fd_sc_hd__and3_2
X_14670_ rvcpu.dp.plmw.ALUResultW\[13\] rvcpu.dp.plmw.ReadDataW\[13\] rvcpu.dp.plmw.PCPlus4W\[13\]
+ rvcpu.dp.plmw.lAuiPCW\[13\] _13169_ _13171_ VGND VGND VPWR VPWR _13237_ sky130_fd_sc_hd__mux4_2
XFILLER_0_19_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25607_ _10727_ net3560 net53 VGND VGND VPWR VPWR _11068_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29375_ clknet_leaf_144_clk _01110_ VGND VGND VPWR VPWR datamem.data_ram\[60\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__10156_ clknet_0__10156_ VGND VGND VPWR VPWR clknet_1_1__leaf__10156_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_39_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22819_ rvcpu.dp.rf.reg_file_arr\[20\]\[27\] rvcpu.dp.rf.reg_file_arr\[21\]\[27\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[27\] rvcpu.dp.rf.reg_file_arr\[23\]\[27\] _09512_
+ _09408_ VGND VGND VPWR VPWR _09958_ sky130_fd_sc_hd__mux4_1
X_26587_ _10297_ _10935_ _11609_ VGND VGND VPWR VPWR _11640_ sky130_fd_sc_hd__and3_2
XFILLER_0_183_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_184_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16340_ net2287 _14438_ _14525_ VGND VGND VPWR VPWR _14534_ sky130_fd_sc_hd__mux2_1
X_28326_ _12365_ net2890 _12632_ VGND VGND VPWR VPWR _12637_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25538_ _10735_ net3383 _11021_ VGND VGND VPWR VPWR _11027_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__10087_ clknet_0__10087_ VGND VGND VPWR VPWR clknet_1_1__leaf__10087_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_137_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28257_ _12598_ VGND VGND VPWR VPWR _03948_ sky130_fd_sc_hd__clkbuf_1
X_16271_ _14497_ VGND VGND VPWR VPWR _01900_ sky130_fd_sc_hd__clkbuf_1
X_25469_ _10954_ net1435 _10984_ _10990_ VGND VGND VPWR VPWR _02768_ sky130_fd_sc_hd__a31o_1
XFILLER_0_192_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18010_ _05321_ rvcpu.dp.SrcBFW_Mux.y\[2\] _05379_ VGND VGND VPWR VPWR _05380_ sky130_fd_sc_hd__o21a_2
X_15222_ _13397_ _13282_ VGND VGND VPWR VPWR _13763_ sky130_fd_sc_hd__nor2_1
X_27208_ _11976_ _12008_ VGND VGND VPWR VPWR _12014_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28188_ _12561_ VGND VGND VPWR VPWR _03916_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15153_ _13333_ _13344_ VGND VGND VPWR VPWR _13697_ sky130_fd_sc_hd__nand2_1
X_27139_ _11956_ net1531 _11964_ _11971_ VGND VGND VPWR VPWR _03457_ sky130_fd_sc_hd__a31o_1
XFILLER_0_62_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_101_clk clknet_5_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_101_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_129_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23337__975 clknet_1_0__leaf__10136_ VGND VGND VPWR VPWR net1101 sky130_fd_sc_hd__inv_2
X_15084_ _13282_ _13317_ VGND VGND VPWR VPWR _13630_ sky130_fd_sc_hd__nand2_1
X_19961_ datamem.data_ram\[2\]\[18\] _06612_ _06648_ datamem.data_ram\[0\]\[18\] _07254_
+ VGND VGND VPWR VPWR _07255_ sky130_fd_sc_hd__o221a_1
X_30150_ net512 _01885_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[0\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18912_ _05535_ _05536_ VGND VGND VPWR VPWR _06252_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19892_ datamem.data_ram\[16\]\[17\] _06648_ _06707_ datamem.data_ram\[23\]\[17\]
+ VGND VGND VPWR VPWR _07187_ sky130_fd_sc_hd__o22a_1
X_30081_ net443 _01816_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[11\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_224_5880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18843_ _05486_ _05785_ _05732_ _05487_ VGND VGND VPWR VPWR _06188_ sky130_fd_sc_hd__o22ai_1
XTAP_TAPCELL_ROW_8_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_220_5766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18774_ _05311_ _06106_ _05335_ VGND VGND VPWR VPWR _06123_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_220_5777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15986_ _14330_ VGND VGND VPWR VPWR _02034_ sky130_fd_sc_hd__clkbuf_1
X_17725_ _05137_ VGND VGND VPWR VPWR _01178_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14937_ _13476_ _13479_ _13480_ _13485_ VGND VGND VPWR VPWR _13486_ sky130_fd_sc_hd__and4b_1
X_30983_ clknet_leaf_115_clk _02718_ VGND VGND VPWR VPWR datamem.data_ram\[39\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_168_clk clknet_5_24__leaf_clk VGND VGND VPWR VPWR clknet_leaf_168_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_175_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32722_ clknet_leaf_212_clk _04144_ VGND VGND VPWR VPWR datamem.data_ram\[16\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17656_ net2714 _13234_ _05093_ VGND VGND VPWR VPWR _05101_ sky130_fd_sc_hd__mux2_1
X_14868_ _13419_ _13293_ VGND VGND VPWR VPWR _13420_ sky130_fd_sc_hd__nand2_4
XFILLER_0_216_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16607_ _14139_ net3303 _04540_ VGND VGND VPWR VPWR _04545_ sky130_fd_sc_hd__mux2_1
X_32653_ clknet_leaf_237_clk _04075_ VGND VGND VPWR VPWR datamem.data_ram\[19\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17587_ _05064_ VGND VGND VPWR VPWR _01243_ sky130_fd_sc_hd__clkbuf_1
X_14799_ _13314_ _13331_ VGND VGND VPWR VPWR _13352_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31604_ clknet_leaf_29_clk net1178 VGND VGND VPWR VPWR rvcpu.dp.plmw.PCPlus4W\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_19326_ rvcpu.dp.plem.ALUResultM\[4\] VGND VGND VPWR VPWR _06622_ sky130_fd_sc_hd__inv_4
XFILLER_0_161_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16538_ _14139_ net2806 _04503_ VGND VGND VPWR VPWR _04508_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32584_ clknet_leaf_183_clk _04006_ VGND VGND VPWR VPWR datamem.data_ram\[21\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_190_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19257_ _06559_ VGND VGND VPWR VPWR rvcpu.dp.lAuiPCE\[30\] sky130_fd_sc_hd__clkbuf_1
X_31535_ clknet_leaf_17_clk net1172 VGND VGND VPWR VPWR rvcpu.dp.plem.PCPlus4M\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16469_ _04471_ VGND VGND VPWR VPWR _01808_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_183_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_4596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18208_ _05563_ _05572_ VGND VGND VPWR VPWR _05573_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_3201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19188_ _06499_ rvcpu.dp.plde.ImmExtE\[21\] _06493_ VGND VGND VPWR VPWR _06500_ sky130_fd_sc_hd__mux2_1
X_31466_ clknet_leaf_2_clk rvcpu.dp.SrcBFW_Mux.y\[24\] VGND VGND VPWR VPWR rvcpu.dp.plem.WriteDataM\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_113_3212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18139_ rvcpu.dp.plem.ALUResultM\[16\] _05268_ VGND VGND VPWR VPWR _05505_ sky130_fd_sc_hd__and2_1
X_30417_ net755 _02152_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[31\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31397_ clknet_leaf_49_clk _03100_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCE\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_184_4902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold102 rvcpu.dp.plde.RdE\[3\] VGND VGND VPWR VPWR net1252 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_184_4913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold113 rvcpu.dp.plde.funct3E\[1\] VGND VGND VPWR VPWR net1263 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__10245_ clknet_0__10245_ VGND VGND VPWR VPWR clknet_1_0__leaf__10245_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_223_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold124 rvcpu.dp.plem.ALUResultM\[27\] VGND VGND VPWR VPWR net1274 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold135 rvcpu.dp.plem.ALUResultM\[21\] VGND VGND VPWR VPWR net1285 sky130_fd_sc_hd__dlygate4sd3_1
X_21150_ datamem.data_ram\[23\]\[23\] _06667_ _06653_ datamem.data_ram\[17\]\[23\]
+ VGND VGND VPWR VPWR _08439_ sky130_fd_sc_hd__o22a_1
X_30348_ net694 _02083_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[4\]\[31\] sky130_fd_sc_hd__dfxtp_1
Xhold146 rvcpu.dp.plfd.InstrD\[25\] VGND VGND VPWR VPWR net1296 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold157 datamem.data_ram\[40\]\[4\] VGND VGND VPWR VPWR net1307 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__10176_ clknet_0__10176_ VGND VGND VPWR VPWR clknet_1_0__leaf__10176_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_74_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold168 datamem.data_ram\[43\]\[0\] VGND VGND VPWR VPWR net1318 sky130_fd_sc_hd__dlygate4sd3_1
X_20101_ datamem.data_ram\[7\]\[10\] _07020_ _07391_ _07394_ VGND VGND VPWR VPWR _07395_
+ sky130_fd_sc_hd__o211a_1
Xhold179 datamem.data_ram\[44\]\[3\] VGND VGND VPWR VPWR net1329 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21081_ _06605_ datamem.data_ram\[35\]\[7\] _07825_ datamem.data_ram\[34\]\[7\] _07844_
+ VGND VGND VPWR VPWR _08370_ sky130_fd_sc_hd__o221a_1
X_30279_ clknet_leaf_144_clk _02014_ VGND VGND VPWR VPWR datamem.data_ram\[58\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32018_ clknet_leaf_129_clk _03440_ VGND VGND VPWR VPWR datamem.data_ram\[51\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_6_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20032_ datamem.data_ram\[24\]\[26\] _06695_ _07243_ datamem.data_ram\[25\]\[26\]
+ _07325_ VGND VGND VPWR VPWR _07326_ sky130_fd_sc_hd__o221a_1
XFILLER_0_42_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_143_3920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24840_ _10446_ net2939 _10631_ VGND VGND VPWR VPWR _10635_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_213_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_159_clk clknet_5_25__leaf_clk VGND VGND VPWR VPWR clknet_leaf_159_clk
+ sky130_fd_sc_hd__clkbuf_8
X_21983_ _06585_ rvcpu.dp.plem.MemWriteM VGND VGND VPWR VPWR _09213_ sky130_fd_sc_hd__nand2_2
X_24771_ _10595_ VGND VGND VPWR VPWR _02465_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20934_ datamem.data_ram\[33\]\[22\] _07133_ _08223_ _06603_ VGND VGND VPWR VPWR
+ _08224_ sky130_fd_sc_hd__a211o_1
X_23722_ clknet_1_1__leaf__10192_ VGND VGND VPWR VPWR _10198_ sky130_fd_sc_hd__buf_1
XFILLER_0_179_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27490_ _12175_ VGND VGND VPWR VPWR _03604_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0__10110_ _10110_ VGND VGND VPWR VPWR clknet_0__10110_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_7_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26441_ _06484_ _11539_ _11529_ _11202_ _11571_ VGND VGND VPWR VPWR _11572_ sky130_fd_sc_hd__a221o_1
XFILLER_0_178_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20865_ datamem.data_ram\[38\]\[14\] _07860_ _07851_ datamem.data_ram\[34\]\[14\]
+ _08154_ VGND VGND VPWR VPWR _08155_ sky130_fd_sc_hd__o221a_1
XFILLER_0_193_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29160_ _09239_ net3544 net64 VGND VGND VPWR VPWR _13097_ sky130_fd_sc_hd__mux2_1
X_22604_ rvcpu.dp.rf.reg_file_arr\[8\]\[15\] rvcpu.dp.rf.reg_file_arr\[10\]\[15\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[15\] rvcpu.dp.rf.reg_file_arr\[11\]\[15\] _09608_
+ _09532_ VGND VGND VPWR VPWR _09755_ sky130_fd_sc_hd__mux4_1
XFILLER_0_3_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26372_ _11517_ net1373 _11510_ _11520_ VGND VGND VPWR VPWR _03141_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_42_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20796_ datamem.data_ram\[38\]\[30\] datamem.data_ram\[39\]\[30\] _07835_ VGND VGND
+ VPWR VPWR _08086_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28111_ _12359_ net3289 net74 VGND VGND VPWR VPWR _12521_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22535_ rvcpu.dp.rf.reg_file_arr\[20\]\[12\] rvcpu.dp.rf.reg_file_arr\[21\]\[12\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[12\] rvcpu.dp.rf.reg_file_arr\[23\]\[12\] _09384_
+ _09430_ VGND VGND VPWR VPWR _09689_ sky130_fd_sc_hd__mux4_1
XFILLER_0_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25323_ _10906_ VGND VGND VPWR VPWR _02706_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_221_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29091_ _13060_ VGND VGND VPWR VPWR _04320_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_137_3779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22963__672 clknet_1_1__leaf__10081_ VGND VGND VPWR VPWR net798 sky130_fd_sc_hd__inv_2
XFILLER_0_174_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28042_ _12484_ VGND VGND VPWR VPWR _03847_ sky130_fd_sc_hd__clkbuf_1
X_25254_ _10142_ _10049_ _10052_ VGND VGND VPWR VPWR _10868_ sky130_fd_sc_hd__and3_2
XFILLER_0_162_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22466_ rvcpu.dp.rf.reg_file_arr\[4\]\[8\] rvcpu.dp.rf.reg_file_arr\[5\]\[8\] rvcpu.dp.rf.reg_file_arr\[6\]\[8\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[8\] _09604_ _09424_ VGND VGND VPWR VPWR _09624_ sky130_fd_sc_hd__mux4_1
XFILLER_0_134_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21417_ rvcpu.dp.rf.reg_file_arr\[28\]\[3\] rvcpu.dp.rf.reg_file_arr\[30\]\[3\] rvcpu.dp.rf.reg_file_arr\[29\]\[3\]
+ rvcpu.dp.rf.reg_file_arr\[31\]\[3\] _08533_ _08636_ VGND VGND VPWR VPWR _08676_
+ sky130_fd_sc_hd__mux4_1
X_24205_ _09310_ net3379 _10270_ VGND VGND VPWR VPWR _10273_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25185_ _10830_ VGND VGND VPWR VPWR _02644_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22397_ _09381_ VGND VGND VPWR VPWR _09558_ sky130_fd_sc_hd__buf_4
X_23059__758 clknet_1_0__leaf__10091_ VGND VGND VPWR VPWR net884 sky130_fd_sc_hd__inv_2
X_21348_ _05747_ _05794_ _08608_ _08609_ VGND VGND VPWR VPWR _08610_ sky130_fd_sc_hd__or4_1
X_29993_ net363 _01728_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[14\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_23436__87 clknet_1_1__leaf__10155_ VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__inv_2
XFILLER_0_102_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28944_ _12734_ net3680 net67 VGND VGND VPWR VPWR _12979_ sky130_fd_sc_hd__mux2_1
Xhold680 rvcpu.dp.pcreg.q\[13\] VGND VGND VPWR VPWR net1830 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21279_ _08540_ VGND VGND VPWR VPWR _08541_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold691 datamem.data_ram\[25\]\[6\] VGND VGND VPWR VPWR net1841 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_200_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28875_ _12751_ net2255 _12941_ VGND VGND VPWR VPWR _12942_ sky130_fd_sc_hd__mux2_1
X_15840_ net2175 _13226_ _14247_ VGND VGND VPWR VPWR _14252_ sky130_fd_sc_hd__mux2_1
X_27826_ _10668_ _12325_ _12356_ VGND VGND VPWR VPWR _12357_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_200_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2070 datamem.data_ram\[49\]\[25\] VGND VGND VPWR VPWR net3220 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2081 datamem.data_ram\[43\]\[24\] VGND VGND VPWR VPWR net3231 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_189_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23721__314 clknet_1_1__leaf__10197_ VGND VGND VPWR VPWR net440 sky130_fd_sc_hd__inv_2
Xhold2092 rvcpu.dp.rf.reg_file_arr\[2\]\[3\] VGND VGND VPWR VPWR net3242 sky130_fd_sc_hd__dlygate4sd3_1
X_27757_ _12318_ VGND VGND VPWR VPWR _03728_ sky130_fd_sc_hd__clkbuf_1
X_15771_ _14160_ net4051 _14210_ VGND VGND VPWR VPWR _14215_ sky130_fd_sc_hd__mux2_1
X_24969_ _10400_ net2190 _10696_ VGND VGND VPWR VPWR _10704_ sky130_fd_sc_hd__mux2_1
Xhold1380 datamem.data_ram\[22\]\[22\] VGND VGND VPWR VPWR net2530 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17510_ _13220_ net3124 _05021_ VGND VGND VPWR VPWR _05024_ sky130_fd_sc_hd__mux2_1
Xhold1391 rvcpu.dp.rf.reg_file_arr\[27\]\[2\] VGND VGND VPWR VPWR net2541 sky130_fd_sc_hd__dlygate4sd3_1
X_26708_ _10820_ net4194 _11704_ VGND VGND VPWR VPWR _11709_ sky130_fd_sc_hd__mux2_1
X_14722_ _13276_ VGND VGND VPWR VPWR _03173_ sky130_fd_sc_hd__clkbuf_1
X_18490_ _05679_ _05664_ _05851_ VGND VGND VPWR VPWR _05852_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_87_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27688_ _12128_ net2920 _12280_ VGND VGND VPWR VPWR _12282_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_520 _13251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_531 _14432_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29427_ clknet_leaf_84_clk _01162_ VGND VGND VPWR VPWR datamem.data_ram\[5\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_542 _06744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_1_1__f__10208_ clknet_0__10208_ VGND VGND VPWR VPWR clknet_1_1__leaf__10208_
+ sky130_fd_sc_hd__clkbuf_16
X_17441_ _04987_ VGND VGND VPWR VPWR _01320_ sky130_fd_sc_hd__clkbuf_1
X_26639_ _11665_ net1794 _11662_ _11666_ VGND VGND VPWR VPWR _03262_ sky130_fd_sc_hd__a31o_1
XANTENNA_553 _07845_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14653_ _13224_ VGND VGND VPWR VPWR _03190_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_564 _13254_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_200_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0__10239_ _10239_ VGND VGND VPWR VPWR clknet_0__10239_ sky130_fd_sc_hd__clkbuf_16
X_29358_ clknet_leaf_173_clk _01093_ VGND VGND VPWR VPWR datamem.data_ram\[61\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__10139_ clknet_0__10139_ VGND VGND VPWR VPWR clknet_1_1__leaf__10139_
+ sky130_fd_sc_hd__clkbuf_16
X_17372_ _14154_ net4274 _04949_ VGND VGND VPWR VPWR _04951_ sky130_fd_sc_hd__mux2_1
X_14584_ _13168_ VGND VGND VPWR VPWR _13169_ sky130_fd_sc_hd__clkbuf_8
X_19111_ _06429_ _06431_ VGND VGND VPWR VPWR _06432_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_188_5002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28309_ _12456_ net3698 net72 VGND VGND VPWR VPWR _12628_ sky130_fd_sc_hd__mux2_1
X_16323_ _14524_ VGND VGND VPWR VPWR _14525_ sky130_fd_sc_hd__buf_4
XFILLER_0_131_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_188_5013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29289_ _09325_ net3793 _13159_ VGND VGND VPWR VPWR _13166_ sky130_fd_sc_hd__mux2_1
X_19042_ _06371_ rvcpu.dp.plde.ImmExtE\[3\] _06355_ VGND VGND VPWR VPWR _06372_ sky130_fd_sc_hd__mux2_1
X_31320_ clknet_leaf_26_clk _03023_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCPlus4E\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16254_ _14234_ _14273_ VGND VGND VPWR VPWR _14488_ sky130_fd_sc_hd__nor2_2
X_15205_ _13350_ _13545_ VGND VGND VPWR VPWR _13747_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_207_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31251_ clknet_leaf_21_clk _02954_ VGND VGND VPWR VPWR rvcpu.dp.plfd.InstrD\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_515 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16185_ _14441_ VGND VGND VPWR VPWR _01938_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_112_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30202_ net556 _01937_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[8\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_226_5920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15136_ _13638_ _13652_ _13662_ _13670_ _13680_ VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__a32o_1
XFILLER_0_11_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_226_5931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31182_ clknet_leaf_37_clk _02885_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCPlus4D\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_147_4020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23270__915 clknet_1_0__leaf__10129_ VGND VGND VPWR VPWR net1041 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_147_4031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30133_ net495 _01868_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[10\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_15067_ _13284_ _13372_ VGND VGND VPWR VPWR _13613_ sky130_fd_sc_hd__nor2_1
X_19944_ datamem.data_ram\[47\]\[18\] _06707_ _07237_ _06602_ VGND VGND VPWR VPWR
+ _07238_ sky130_fd_sc_hd__o211a_1
X_23882__443 clknet_1_1__leaf__10221_ VGND VGND VPWR VPWR net569 sky130_fd_sc_hd__inv_2
XFILLER_0_10_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_222_5817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_1275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_222_5828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30064_ net426 _01799_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[12\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_19875_ datamem.data_ram\[28\]\[1\] _07123_ _07166_ _07169_ VGND VGND VPWR VPWR _07170_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_219_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_207_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18826_ _06171_ VGND VGND VPWR VPWR _06172_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18757_ _05311_ _06106_ VGND VGND VPWR VPWR _06107_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_175_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15969_ _14321_ VGND VGND VPWR VPWR _02042_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_222_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17708_ _05128_ VGND VGND VPWR VPWR _01186_ sky130_fd_sc_hd__clkbuf_1
X_18688_ _05809_ _06040_ _06041_ VGND VGND VPWR VPWR _06042_ sky130_fd_sc_hd__and3_1
X_30966_ clknet_leaf_228_clk _02701_ VGND VGND VPWR VPWR datamem.data_ram\[39\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_177_4750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32705_ clknet_leaf_79_clk _04127_ VGND VGND VPWR VPWR datamem.data_ram\[17\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17639_ net3001 _13209_ _05082_ VGND VGND VPWR VPWR _05092_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30897_ clknet_leaf_151_clk _02632_ VGND VGND VPWR VPWR datamem.data_ram\[41\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_173_4636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_173_4647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_4658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20650_ _07935_ _07940_ _06797_ VGND VGND VPWR VPWR _07941_ sky130_fd_sc_hd__o21a_1
X_32636_ clknet_leaf_255_clk _04058_ VGND VGND VPWR VPWR datamem.data_ram\[1\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19309_ _05185_ VGND VGND VPWR VPWR _06605_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_184_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32567_ clknet_leaf_83_clk _03989_ VGND VGND VPWR VPWR datamem.data_ram\[22\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_20581_ rvcpu.dp.plem.ALUResultM\[7\] _06592_ VGND VGND VPWR VPWR _07872_ sky130_fd_sc_hd__nand2_8
XFILLER_0_2_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22320_ _09484_ VGND VGND VPWR VPWR _09485_ sky130_fd_sc_hd__buf_4
X_31518_ clknet_leaf_52_clk net1239 VGND VGND VPWR VPWR rvcpu.dp.plem.PCPlus4M\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32498_ clknet_leaf_286_clk _03920_ VGND VGND VPWR VPWR datamem.data_ram\[25\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_76_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22251_ _09416_ VGND VGND VPWR VPWR _09417_ sky130_fd_sc_hd__clkbuf_8
X_31449_ clknet_leaf_7_clk rvcpu.dp.SrcBFW_Mux.y\[7\] VGND VGND VPWR VPWR rvcpu.dp.plem.WriteDataM\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_132_3654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_3665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21202_ _08483_ VGND VGND VPWR VPWR _04419_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22182_ _09363_ VGND VGND VPWR VPWR _01108_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__10228_ clknet_0__10228_ VGND VGND VPWR VPWR clknet_1_0__leaf__10228_
+ sky130_fd_sc_hd__clkbuf_16
X_21133_ _06678_ _08412_ _08415_ _08419_ _08421_ VGND VGND VPWR VPWR _08422_ sky130_fd_sc_hd__o32a_1
XFILLER_0_2_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26990_ _11879_ VGND VGND VPWR VPWR _03400_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__10159_ clknet_0__10159_ VGND VGND VPWR VPWR clknet_1_0__leaf__10159_
+ sky130_fd_sc_hd__clkbuf_16
X_23132__808 clknet_1_0__leaf__10106_ VGND VGND VPWR VPWR net934 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_35_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25941_ net1859 _11290_ _11286_ _11292_ VGND VGND VPWR VPWR _02938_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_35_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21064_ _07872_ _08311_ _08325_ _08352_ VGND VGND VPWR VPWR _08353_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_10_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20015_ datamem.data_ram\[55\]\[2\] _06926_ _07305_ _07308_ VGND VGND VPWR VPWR _07309_
+ sky130_fd_sc_hd__a211o_1
X_28660_ _12827_ VGND VGND VPWR VPWR _04122_ sky130_fd_sc_hd__clkbuf_1
X_25872_ rvcpu.dp.plfd.PCPlus4D\[30\] _11249_ _08598_ VGND VGND VPWR VPWR _11250_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_31_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27611_ _12155_ net2563 _12233_ VGND VGND VPWR VPWR _12240_ sky130_fd_sc_hd__mux2_1
X_24823_ _10625_ VGND VGND VPWR VPWR _02487_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_216_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28591_ _12790_ VGND VGND VPWR VPWR _04090_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_214_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_179_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27542_ _12203_ VGND VGND VPWR VPWR _03628_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24754_ _10586_ VGND VGND VPWR VPWR _02457_ sky130_fd_sc_hd__clkbuf_1
X_21966_ rvcpu.dp.rf.reg_file_arr\[28\]\[31\] rvcpu.dp.rf.reg_file_arr\[30\]\[31\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[31\] rvcpu.dp.rf.reg_file_arr\[31\]\[31\] rvcpu.dp.plfd.InstrD\[16\]
+ _08516_ VGND VGND VPWR VPWR _09197_ sky130_fd_sc_hd__mux4_2
XFILLER_0_16_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20917_ datamem.data_ram\[26\]\[22\] _06692_ _06635_ datamem.data_ram\[27\]\[22\]
+ _08206_ VGND VGND VPWR VPWR _08207_ sky130_fd_sc_hd__o221a_1
XFILLER_0_55_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27473_ _12093_ net2219 _12159_ VGND VGND VPWR VPWR _12166_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21897_ _08742_ _09131_ VGND VGND VPWR VPWR _09132_ sky130_fd_sc_hd__or2_1
X_24685_ _10549_ VGND VGND VPWR VPWR _02425_ sky130_fd_sc_hd__clkbuf_1
X_29212_ _11533_ net1667 _13122_ _13125_ VGND VGND VPWR VPWR _04376_ sky130_fd_sc_hd__a31o_1
XFILLER_0_7_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26424_ _11545_ rvcpu.ALUResultE\[14\] VGND VGND VPWR VPWR _11560_ sky130_fd_sc_hd__and2_1
XFILLER_0_167_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23636_ _10184_ VGND VGND VPWR VPWR _01741_ sky130_fd_sc_hd__clkbuf_1
X_20848_ datamem.data_ram\[4\]\[14\] datamem.data_ram\[5\]\[14\] _07849_ VGND VGND
+ VPWR VPWR _08138_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_182_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29143_ _09275_ net2757 net39 VGND VGND VPWR VPWR _13088_ sky130_fd_sc_hd__mux2_1
X_26355_ _09226_ _10935_ _10052_ VGND VGND VPWR VPWR _11511_ sky130_fd_sc_hd__and3_2
XFILLER_0_147_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20779_ _08023_ _08037_ _08053_ _08068_ VGND VGND VPWR VPWR _08069_ sky130_fd_sc_hd__or4_2
XFILLER_0_37_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25306_ _08124_ _07903_ VGND VGND VPWR VPWR _10896_ sky130_fd_sc_hd__or2_2
X_29074_ _13051_ VGND VGND VPWR VPWR _04312_ sky130_fd_sc_hd__clkbuf_1
X_22518_ _09671_ _09672_ _09449_ VGND VGND VPWR VPWR _09673_ sky130_fd_sc_hd__mux2_1
X_26286_ _11475_ VGND VGND VPWR VPWR _03100_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28025_ _12433_ net3364 _12473_ VGND VGND VPWR VPWR _12475_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_21_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22449_ _09430_ VGND VGND VPWR VPWR _09608_ sky130_fd_sc_hd__clkbuf_8
X_25237_ _10858_ VGND VGND VPWR VPWR _02668_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25168_ _10818_ net4022 net58 VGND VGND VPWR VPWR _10819_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_206_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25099_ _10064_ _10779_ _10781_ net1299 VGND VGND VPWR VPWR _02607_ sky130_fd_sc_hd__a22o_1
X_17990_ _05358_ _05359_ VGND VGND VPWR VPWR _05360_ sky130_fd_sc_hd__nor2_1
X_29976_ net346 _01711_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[14\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28927_ _12969_ VGND VGND VPWR VPWR _04247_ sky130_fd_sc_hd__clkbuf_1
X_16941_ net1868 _14424_ _04720_ VGND VGND VPWR VPWR _04722_ sky130_fd_sc_hd__mux2_1
XFILLER_0_202_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_217_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19660_ datamem.data_ram\[38\]\[0\] _06952_ _06955_ datamem.data_ram\[36\]\[0\] VGND
+ VGND VPWR VPWR _06956_ sky130_fd_sc_hd__a22o_1
XFILLER_0_159_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28858_ _12687_ net3491 _12932_ VGND VGND VPWR VPWR _12933_ sky130_fd_sc_hd__mux2_1
X_16872_ _04685_ VGND VGND VPWR VPWR _01603_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_217_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18611_ _05705_ _05850_ _05968_ _05776_ VGND VGND VPWR VPWR _05969_ sky130_fd_sc_hd__a211o_1
X_27809_ _12347_ VGND VGND VPWR VPWR _03751_ sky130_fd_sc_hd__clkbuf_1
X_15823_ net2395 _13201_ _14236_ VGND VGND VPWR VPWR _14243_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19591_ datamem.data_ram\[58\]\[8\] _06610_ _06821_ datamem.data_ram\[56\]\[8\] VGND
+ VGND VPWR VPWR _06887_ sky130_fd_sc_hd__o22a_1
X_28789_ _12601_ _11020_ _12886_ VGND VGND VPWR VPWR _12896_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_189_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18542_ _05704_ _05900_ _05902_ VGND VGND VPWR VPWR _05903_ sky130_fd_sc_hd__o21ai_1
X_30820_ clknet_leaf_172_clk _02555_ VGND VGND VPWR VPWR datamem.data_ram\[45\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15754_ _14143_ net4319 _14199_ VGND VGND VPWR VPWR _14206_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14705_ net2181 _13263_ _13245_ VGND VGND VPWR VPWR _13264_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18473_ _05818_ _05835_ VGND VGND VPWR VPWR _05836_ sky130_fd_sc_hd__or2_1
X_30751_ clknet_leaf_179_clk _02486_ VGND VGND VPWR VPWR datamem.data_ram\[48\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_15685_ _14160_ net4066 _14152_ VGND VGND VPWR VPWR _14161_ sky130_fd_sc_hd__mux2_1
XANTENNA_350 rvcpu.ALUResultE\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_361 rvcpu.dp.SrcBFW_Mux.y\[22\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_372 rvcpu.dp.plem.ALUResultM\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17424_ _04978_ VGND VGND VPWR VPWR _01328_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_383 net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14636_ _13211_ VGND VGND VPWR VPWR _03194_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_215_5654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30682_ clknet_leaf_96_clk _02417_ VGND VGND VPWR VPWR datamem.data_ram\[4\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24131__636 clknet_1_0__leaf__10261_ VGND VGND VPWR VPWR net762 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_215_5665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_394 clknet_1_1__leaf__10087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32421_ clknet_leaf_78_clk _03843_ VGND VGND VPWR VPWR datamem.data_ram\[28\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17355_ _14137_ net2384 _04938_ VGND VGND VPWR VPWR _04942_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16306_ net3418 _14472_ _14511_ VGND VGND VPWR VPWR _14516_ sky130_fd_sc_hd__mux2_1
X_32352_ clknet_leaf_170_clk _03774_ VGND VGND VPWR VPWR datamem.data_ram\[30\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17286_ _04905_ VGND VGND VPWR VPWR _01401_ sky130_fd_sc_hd__clkbuf_1
Xclkload303 clknet_1_1__leaf__10202_ VGND VGND VPWR VPWR clkload303/Y sky130_fd_sc_hd__clkinvlp_4
X_31303_ clknet_leaf_48_clk _03006_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCPlus4E\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_19025_ rvcpu.dp.plde.ImmExtE\[1\] rvcpu.dp.plde.PCE\[1\] VGND VGND VPWR VPWR _06357_
+ sky130_fd_sc_hd__xor2_2
XFILLER_0_181_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload11 clknet_5_13__leaf_clk VGND VGND VPWR VPWR clkload11/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_113_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload314 clknet_1_1__leaf__10179_ VGND VGND VPWR VPWR clkload314/Y sky130_fd_sc_hd__clkinvlp_4
X_16237_ net3264 _14476_ _14464_ VGND VGND VPWR VPWR _14477_ sky130_fd_sc_hd__mux2_1
Xclkload22 clknet_5_27__leaf_clk VGND VGND VPWR VPWR clkload22/Y sky130_fd_sc_hd__inv_6
Xclkload325 clknet_1_1__leaf__11602_ VGND VGND VPWR VPWR clkload325/Y sky130_fd_sc_hd__clkinvlp_4
X_32283_ clknet_leaf_241_clk _03705_ VGND VGND VPWR VPWR datamem.data_ram\[33\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload33 clknet_leaf_13_clk VGND VGND VPWR VPWR clkload33/Y sky130_fd_sc_hd__clkinv_1
Xclkload336 clknet_1_1__leaf__10132_ VGND VGND VPWR VPWR clkload336/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload44 clknet_leaf_34_clk VGND VGND VPWR VPWR clkload44/Y sky130_fd_sc_hd__clkinv_4
Xclkload347 clknet_1_0__leaf__10087_ VGND VGND VPWR VPWR clkload347/X sky130_fd_sc_hd__clkbuf_8
Xclkload358 clknet_1_1__leaf__10082_ VGND VGND VPWR VPWR clkload358/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload55 clknet_leaf_282_clk VGND VGND VPWR VPWR clkload55/Y sky130_fd_sc_hd__clkinv_4
X_31234_ clknet_leaf_31_clk _02937_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCD\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload66 clknet_leaf_63_clk VGND VGND VPWR VPWR clkload66/X sky130_fd_sc_hd__clkbuf_4
X_16168_ _13194_ VGND VGND VPWR VPWR _14430_ sky130_fd_sc_hd__clkbuf_4
Xclkload77 clknet_leaf_38_clk VGND VGND VPWR VPWR clkload77/Y sky130_fd_sc_hd__bufinv_16
Xclkload88 clknet_leaf_52_clk VGND VGND VPWR VPWR clkload88/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_71_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload99 clknet_leaf_85_clk VGND VGND VPWR VPWR clkload99/Y sky130_fd_sc_hd__inv_6
XFILLER_0_62_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15119_ _13412_ _13549_ _13663_ _13357_ VGND VGND VPWR VPWR _13664_ sky130_fd_sc_hd__o31a_1
X_31165_ clknet_leaf_9_clk rvcpu.ALUResultE\[24\] VGND VGND VPWR VPWR rvcpu.dp.plem.ALUResultM\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16099_ _14391_ VGND VGND VPWR VPWR _01974_ sky130_fd_sc_hd__clkbuf_1
X_23415__68 clknet_1_1__leaf__10153_ VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_166_4473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_166_4484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30116_ net478 _01851_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[10\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_19927_ datamem.data_ram\[51\]\[17\] _06863_ _07221_ _06776_ VGND VGND VPWR VPWR
+ _07222_ sky130_fd_sc_hd__o211a_1
Xhold2806 datamem.data_ram\[20\]\[27\] VGND VGND VPWR VPWR net3956 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2817 datamem.data_ram\[31\]\[8\] VGND VGND VPWR VPWR net3967 sky130_fd_sc_hd__dlygate4sd3_1
X_31096_ clknet_leaf_257_clk _02831_ VGND VGND VPWR VPWR datamem.data_ram\[9\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2828 datamem.data_ram\[40\]\[29\] VGND VGND VPWR VPWR net3978 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2839 datamem.data_ram\[63\]\[20\] VGND VGND VPWR VPWR net3989 sky130_fd_sc_hd__dlygate4sd3_1
X_30047_ net409 _01782_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[12\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_19858_ _06916_ _07130_ _07141_ _07152_ VGND VGND VPWR VPWR _07153_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_179_4801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18809_ _05313_ _05334_ _05500_ _05506_ _05664_ _05768_ VGND VGND VPWR VPWR _06156_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_69_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19789_ datamem.data_ram\[55\]\[9\] _06707_ _06783_ datamem.data_ram\[49\]\[9\] VGND
+ VGND VPWR VPWR _07084_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_69_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_3491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21820_ _09057_ _09058_ _08743_ VGND VGND VPWR VPWR _09059_ sky130_fd_sc_hd__mux2_1
XFILLER_0_222_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31998_ clknet_leaf_131_clk _03420_ VGND VGND VPWR VPWR datamem.data_ram\[31\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_65_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_195_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21751_ _08626_ _08987_ _08989_ _08993_ _08808_ VGND VGND VPWR VPWR _08994_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_121_3388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30949_ clknet_leaf_260_clk _02684_ VGND VGND VPWR VPWR datamem.data_ram\[3\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_210_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_90_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_90_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_121_3399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20702_ datamem.data_ram\[14\]\[5\] _07127_ _07000_ datamem.data_ram\[10\]\[5\] VGND
+ VGND VPWR VPWR _07993_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24470_ _09314_ net3272 _10421_ VGND VGND VPWR VPWR _10425_ sky130_fd_sc_hd__mux2_1
X_21682_ _08692_ _08926_ _08928_ VGND VGND VPWR VPWR _08929_ sky130_fd_sc_hd__a21o_1
XFILLER_0_176_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20633_ datamem.data_ram\[3\]\[29\] _06635_ _06783_ datamem.data_ram\[1\]\[29\] _07923_
+ VGND VGND VPWR VPWR _07924_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_134_3705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32619_ clknet_leaf_250_clk _04041_ VGND VGND VPWR VPWR datamem.data_ram\[20\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_3716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_199_Left_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26140_ net1897 _11397_ VGND VGND VPWR VPWR _11406_ sky130_fd_sc_hd__and2_1
Xclkload5 clknet_5_6__leaf_clk VGND VGND VPWR VPWR clkload5/Y sky130_fd_sc_hd__inv_6
XFILLER_0_117_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20564_ _07131_ _07846_ _07854_ _07154_ VGND VGND VPWR VPWR _07855_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_24_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_99_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23889__449 clknet_1_1__leaf__10222_ VGND VGND VPWR VPWR net575 sky130_fd_sc_hd__inv_2
XFILLER_0_229_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23750__340 clknet_1_1__leaf__10200_ VGND VGND VPWR VPWR net466 sky130_fd_sc_hd__inv_2
X_22303_ rvcpu.dp.rf.reg_file_arr\[4\]\[1\] rvcpu.dp.rf.reg_file_arr\[5\]\[1\] rvcpu.dp.rf.reg_file_arr\[6\]\[1\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[1\] _09464_ _09467_ VGND VGND VPWR VPWR _09468_ sky130_fd_sc_hd__mux4_1
XFILLER_0_15_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26071_ _11365_ VGND VGND VPWR VPWR _02994_ sky130_fd_sc_hd__clkbuf_1
X_20495_ datamem.data_ram\[34\]\[21\] _06613_ _06701_ datamem.data_ram\[33\]\[21\]
+ VGND VGND VPWR VPWR _07786_ sky130_fd_sc_hd__o22a_1
XFILLER_0_171_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22234_ _08595_ VGND VGND VPWR VPWR _09400_ sky130_fd_sc_hd__clkbuf_8
X_25022_ _09284_ VGND VGND VPWR VPWR _10735_ sky130_fd_sc_hd__buf_2
XFILLER_0_14_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_384 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_5_30__f_clk clknet_2_3_0_clk VGND VGND VPWR VPWR clknet_5_30__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_29830_ net208 _01565_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[1\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_22165_ _09306_ net3011 _09352_ VGND VGND VPWR VPWR _09354_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_218_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21116_ datamem.data_ram\[27\]\[7\] _06941_ _06946_ datamem.data_ram\[25\]\[7\] _08404_
+ VGND VGND VPWR VPWR _08405_ sky130_fd_sc_hd__a221o_2
XFILLER_0_121_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24165__7 clknet_1_1__leaf__10264_ VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__inv_2
XFILLER_0_100_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29761_ net1107 _01496_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[21\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_26973_ _11863_ net1773 _11865_ _11870_ VGND VGND VPWR VPWR _03392_ sky130_fd_sc_hd__a31o_1
X_22096_ rvcpu.dp.plem.WriteDataM\[2\] _08488_ _09293_ VGND VGND VPWR VPWR _09308_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_79_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_227_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28712_ _12696_ net3137 _12850_ VGND VGND VPWR VPWR _12855_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_54_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25924_ net2115 _11279_ VGND VGND VPWR VPWR _11282_ sky130_fd_sc_hd__or2_1
X_21047_ datamem.data_ram\[4\]\[31\] datamem.data_ram\[5\]\[31\] _07912_ VGND VGND
+ VPWR VPWR _08336_ sky130_fd_sc_hd__mux2_1
X_29692_ net1038 _01427_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[23\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_54_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28643_ _12818_ VGND VGND VPWR VPWR _04114_ sky130_fd_sc_hd__clkbuf_1
X_25855_ _11234_ _11235_ VGND VGND VPWR VPWR _11236_ sky130_fd_sc_hd__nor2_1
XFILLER_0_198_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_198_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24806_ _10616_ VGND VGND VPWR VPWR _02479_ sky130_fd_sc_hd__clkbuf_1
X_28574_ _12781_ VGND VGND VPWR VPWR _04082_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25786_ _11143_ VGND VGND VPWR VPWR _11181_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_201_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27525_ _12194_ VGND VGND VPWR VPWR _03620_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_332 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24737_ _10577_ VGND VGND VPWR VPWR _02449_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21949_ rvcpu.dp.rf.reg_file_arr\[24\]\[30\] rvcpu.dp.rf.reg_file_arr\[25\]\[30\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[30\] rvcpu.dp.rf.reg_file_arr\[27\]\[30\] _08549_
+ _08527_ VGND VGND VPWR VPWR _09181_ sky130_fd_sc_hd__mux4_2
XFILLER_0_96_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_81_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_81_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_16_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15470_ _13496_ _13999_ VGND VGND VPWR VPWR _14000_ sky130_fd_sc_hd__nand2_1
X_27456_ _12156_ VGND VGND VPWR VPWR _03589_ sky130_fd_sc_hd__clkbuf_1
X_24668_ _10418_ _10532_ VGND VGND VPWR VPWR _10540_ sky130_fd_sc_hd__and2_1
XFILLER_0_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26407_ _06411_ _11540_ VGND VGND VPWR VPWR _11548_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27387_ _10735_ net2631 _12107_ VGND VGND VPWR VPWR _12113_ sky130_fd_sc_hd__mux2_1
X_24599_ _10500_ VGND VGND VPWR VPWR _10501_ sky130_fd_sc_hd__buf_8
XFILLER_0_182_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29126_ _09239_ net2853 _13076_ VGND VGND VPWR VPWR _13079_ sky130_fd_sc_hd__mux2_1
X_17140_ _14195_ net2659 _04792_ VGND VGND VPWR VPWR _04827_ sky130_fd_sc_hd__mux2_1
X_26338_ _11501_ net1494 _11496_ _11504_ VGND VGND VPWR VPWR _03123_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_210_5540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17071_ _04790_ VGND VGND VPWR VPWR _01501_ sky130_fd_sc_hd__clkbuf_1
X_29057_ _13042_ VGND VGND VPWR VPWR _04304_ sky130_fd_sc_hd__clkbuf_1
X_23948__502 clknet_1_0__leaf__10228_ VGND VGND VPWR VPWR net628 sky130_fd_sc_hd__inv_2
X_26269_ _11466_ VGND VGND VPWR VPWR _03092_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23000__705 clknet_1_1__leaf__10085_ VGND VGND VPWR VPWR net831 sky130_fd_sc_hd__inv_2
XFILLER_0_123_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28008_ _12359_ net2512 net97 VGND VGND VPWR VPWR _12466_ sky130_fd_sc_hd__mux2_1
X_16022_ net1914 _13184_ _14349_ VGND VGND VPWR VPWR _14351_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_208_5480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_208_5491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17973_ _05342_ _05343_ VGND VGND VPWR VPWR _05344_ sky130_fd_sc_hd__and2_1
X_29959_ net329 _01694_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[15\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19712_ datamem.data_ram\[19\]\[0\] _06966_ _07004_ _07007_ VGND VGND VPWR VPWR _07008_
+ sky130_fd_sc_hd__a211o_1
X_16924_ _04712_ VGND VGND VPWR VPWR _01578_ sky130_fd_sc_hd__clkbuf_1
X_32970_ clknet_leaf_141_clk _04392_ VGND VGND VPWR VPWR datamem.data_ram\[63\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_204_5388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_204_5399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_4370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19643_ datamem.data_ram\[37\]\[0\] _06921_ _06927_ datamem.data_ram\[39\]\[0\] _06938_
+ VGND VGND VPWR VPWR _06939_ sky130_fd_sc_hd__a221o_1
X_31921_ _04433_ net119 VGND VGND VPWR VPWR datamem.rd_data_mem\[26\] sky130_fd_sc_hd__dlxtn_1
X_16855_ net2571 _14474_ _04670_ VGND VGND VPWR VPWR _04676_ sky130_fd_sc_hd__mux2_1
XFILLER_0_204_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15806_ _14195_ net2597 _14198_ VGND VGND VPWR VPWR _14233_ sky130_fd_sc_hd__mux2_1
X_23920__476 clknet_1_0__leaf__10226_ VGND VGND VPWR VPWR net602 sky130_fd_sc_hd__inv_2
X_31852_ clknet_leaf_123_clk _03306_ VGND VGND VPWR VPWR datamem.data_ram\[61\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_19574_ datamem.data_ram\[13\]\[8\] _06724_ _06837_ datamem.data_ram\[8\]\[8\] VGND
+ VGND VPWR VPWR _06870_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_196_5189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16786_ _04639_ VGND VGND VPWR VPWR _01651_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_217_5705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18525_ _05812_ VGND VGND VPWR VPWR _05886_ sky130_fd_sc_hd__buf_4
X_30803_ clknet_leaf_192_clk _02538_ VGND VGND VPWR VPWR datamem.data_ram\[45\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15737_ _14195_ net3604 _14130_ VGND VGND VPWR VPWR _14196_ sky130_fd_sc_hd__mux2_1
X_31783_ clknet_leaf_53_clk _03237_ VGND VGND VPWR VPWR datamem.data_ram\[8\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_72_clk clknet_5_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_72_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_153_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18456_ _05370_ _05380_ _05667_ _05576_ _05590_ VGND VGND VPWR VPWR _05819_ sky130_fd_sc_hd__o41a_2
XFILLER_0_29_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30734_ clknet_leaf_227_clk _02469_ VGND VGND VPWR VPWR datamem.data_ram\[47\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15668_ _13209_ VGND VGND VPWR VPWR _14149_ sky130_fd_sc_hd__buf_4
XFILLER_0_75_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_180 _08988_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_213_1084 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23161__834 clknet_1_0__leaf__10109_ VGND VGND VPWR VPWR net960 sky130_fd_sc_hd__inv_2
XANTENNA_191 _09290_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_2_1_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_1_0_clk sky130_fd_sc_hd__clkbuf_8
X_17407_ _14189_ net4262 _04960_ VGND VGND VPWR VPWR _04969_ sky130_fd_sc_hd__mux2_1
X_14619_ net2399 _13198_ _13181_ VGND VGND VPWR VPWR _13199_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18387_ _05574_ _05570_ _05565_ _05566_ _05683_ _05579_ VGND VGND VPWR VPWR _05751_
+ sky130_fd_sc_hd__mux4_1
X_30665_ clknet_leaf_151_clk _02400_ VGND VGND VPWR VPWR datamem.data_ram\[50\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15599_ _14107_ VGND VGND VPWR VPWR _02206_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32404_ clknet_leaf_254_clk _03826_ VGND VGND VPWR VPWR datamem.data_ram\[29\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_17338_ _04932_ VGND VGND VPWR VPWR _01376_ sky130_fd_sc_hd__clkbuf_1
X_30596_ clknet_leaf_118_clk _02331_ VGND VGND VPWR VPWR datamem.data_ram\[53\]\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_83_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23276__921 clknet_1_1__leaf__10129_ VGND VGND VPWR VPWR net1047 sky130_fd_sc_hd__inv_2
Xclkload100 clknet_leaf_86_clk VGND VGND VPWR VPWR clkload100/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_154_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32335_ clknet_leaf_275_clk _03757_ VGND VGND VPWR VPWR datamem.data_ram\[31\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload111 clknet_leaf_98_clk VGND VGND VPWR VPWR clkload111/Y sky130_fd_sc_hd__clkinv_1
XFILLER_0_126_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17269_ _04895_ VGND VGND VPWR VPWR _01408_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_12_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload122 clknet_leaf_107_clk VGND VGND VPWR VPWR clkload122/Y sky130_fd_sc_hd__clkinvlp_2
XTAP_TAPCELL_ROW_12_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_4524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19008_ _05288_ _05732_ _05730_ _05289_ VGND VGND VPWR VPWR _06342_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_12_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload133 clknet_leaf_287_clk VGND VGND VPWR VPWR clkload133/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_168_4535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload144 clknet_leaf_249_clk VGND VGND VPWR VPWR clkload144/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_222_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20280_ _06716_ _07567_ _07572_ VGND VGND VPWR VPWR _07573_ sky130_fd_sc_hd__or3_1
XFILLER_0_3_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32266_ clknet_leaf_228_clk _03688_ VGND VGND VPWR VPWR datamem.data_ram\[33\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload155 clknet_leaf_278_clk VGND VGND VPWR VPWR clkload155/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_11_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload166 clknet_leaf_267_clk VGND VGND VPWR VPWR clkload166/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload177 clknet_leaf_232_clk VGND VGND VPWR VPWR clkload177/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_23_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31217_ clknet_leaf_37_clk _02920_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCD\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload188 clknet_leaf_222_clk VGND VGND VPWR VPWR clkload188/Y sky130_fd_sc_hd__inv_6
Xclkload199 clknet_leaf_189_clk VGND VGND VPWR VPWR clkload199/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_178_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32197_ clknet_leaf_225_clk _03619_ VGND VGND VPWR VPWR datamem.data_ram\[36\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3304 rvcpu.dp.pcreg.q\[20\] VGND VGND VPWR VPWR net4454 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_90_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31148_ clknet_leaf_63_clk rvcpu.ALUResultE\[7\] VGND VGND VPWR VPWR rvcpu.dp.plem.ALUResultM\[7\]
+ sky130_fd_sc_hd__dfxtp_4
Xhold2603 datamem.data_ram\[21\]\[26\] VGND VGND VPWR VPWR net3753 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2614 rvcpu.dp.rf.reg_file_arr\[15\]\[16\] VGND VGND VPWR VPWR net3764 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold17 rvcpu.dp.plem.PCPlus4M\[4\] VGND VGND VPWR VPWR net1167 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2625 datamem.data_ram\[61\]\[27\] VGND VGND VPWR VPWR net3775 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold28 rvcpu.dp.plem.PCPlus4M\[22\] VGND VGND VPWR VPWR net1178 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2636 datamem.data_ram\[43\]\[20\] VGND VGND VPWR VPWR net3786 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_127_3542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31079_ clknet_leaf_107_clk _02814_ VGND VGND VPWR VPWR datamem.data_ram\[20\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_127_3553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1902 datamem.data_ram\[24\]\[28\] VGND VGND VPWR VPWR net3052 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2647 datamem.data_ram\[4\]\[24\] VGND VGND VPWR VPWR net3797 sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 rvcpu.dp.plem.lAuiPCM\[31\] VGND VGND VPWR VPWR net1189 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2658 datamem.data_ram\[24\]\[17\] VGND VGND VPWR VPWR net3808 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1913 datamem.data_ram\[24\]\[21\] VGND VGND VPWR VPWR net3063 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23780__366 clknet_1_1__leaf__10204_ VGND VGND VPWR VPWR net492 sky130_fd_sc_hd__inv_2
Xhold1924 datamem.data_ram\[25\]\[15\] VGND VGND VPWR VPWR net3074 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2669 datamem.data_ram\[62\]\[12\] VGND VGND VPWR VPWR net3819 sky130_fd_sc_hd__dlygate4sd3_1
X_22921_ _10041_ net1825 _10046_ _10054_ VGND VGND VPWR VPWR _01156_ sky130_fd_sc_hd__a31o_1
Xhold1935 datamem.data_ram\[59\]\[12\] VGND VGND VPWR VPWR net3085 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1946 datamem.data_ram\[55\]\[24\] VGND VGND VPWR VPWR net3096 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1957 datamem.data_ram\[45\]\[21\] VGND VGND VPWR VPWR net3107 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_123_3439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1968 rvcpu.dp.rf.reg_file_arr\[27\]\[28\] VGND VGND VPWR VPWR net3118 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_155_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25640_ _10069_ VGND VGND VPWR VPWR _11089_ sky130_fd_sc_hd__clkbuf_4
Xhold1979 datamem.data_ram\[40\]\[12\] VGND VGND VPWR VPWR net3129 sky130_fd_sc_hd__dlygate4sd3_1
X_22852_ rvcpu.dp.rf.reg_file_arr\[20\]\[29\] rvcpu.dp.rf.reg_file_arr\[21\]\[29\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[29\] rvcpu.dp.rf.reg_file_arr\[23\]\[29\] _09384_
+ _09577_ VGND VGND VPWR VPWR _09989_ sky130_fd_sc_hd__mux4_1
XFILLER_0_223_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21803_ rvcpu.dp.rf.reg_file_arr\[28\]\[22\] rvcpu.dp.rf.reg_file_arr\[30\]\[22\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[22\] rvcpu.dp.rf.reg_file_arr\[31\]\[22\] _08552_
+ _08687_ VGND VGND VPWR VPWR _09043_ sky130_fd_sc_hd__mux4_1
X_25571_ _10413_ _11042_ VGND VGND VPWR VPWR _11046_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22783_ rvcpu.dp.rf.reg_file_arr\[28\]\[25\] rvcpu.dp.rf.reg_file_arr\[30\]\[25\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[25\] rvcpu.dp.rf.reg_file_arr\[31\]\[25\] _09382_
+ _09417_ VGND VGND VPWR VPWR _09924_ sky130_fd_sc_hd__mux4_1
XFILLER_0_211_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_63_clk clknet_5_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_63_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27310_ _11972_ _12066_ VGND VGND VPWR VPWR _12070_ sky130_fd_sc_hd__and2_1
X_24522_ _09351_ _10347_ _10366_ VGND VGND VPWR VPWR _10456_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_52_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28290_ _12617_ VGND VGND VPWR VPWR _03962_ sky130_fd_sc_hd__clkbuf_1
X_21734_ rvcpu.dp.rf.reg_file_arr\[12\]\[18\] rvcpu.dp.rf.reg_file_arr\[13\]\[18\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[18\] rvcpu.dp.rf.reg_file_arr\[15\]\[18\] _08578_
+ _08684_ VGND VGND VPWR VPWR _08978_ sky130_fd_sc_hd__mux4_1
XFILLER_0_149_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27241_ _11970_ _12031_ VGND VGND VPWR VPWR _12034_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24453_ _10067_ _10406_ VGND VGND VPWR VPWR _10415_ sky130_fd_sc_hd__and2_1
XFILLER_0_137_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21665_ rvcpu.dp.rf.reg_file_arr\[12\]\[14\] rvcpu.dp.rf.reg_file_arr\[13\]\[14\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[14\] rvcpu.dp.rf.reg_file_arr\[15\]\[14\] _08696_
+ _08568_ VGND VGND VPWR VPWR _08913_ sky130_fd_sc_hd__mux4_1
XFILLER_0_164_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_97_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23674__271 clknet_1_1__leaf__10193_ VGND VGND VPWR VPWR net397 sky130_fd_sc_hd__inv_2
XFILLER_0_46_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_97_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27172_ _11991_ net1631 _11983_ _11992_ VGND VGND VPWR VPWR _03469_ sky130_fd_sc_hd__a31o_1
X_20616_ datamem.data_ram\[24\]\[13\] _06820_ _06780_ datamem.data_ram\[25\]\[13\]
+ VGND VGND VPWR VPWR _07907_ sky130_fd_sc_hd__o22a_1
X_24384_ _09244_ net3992 _10367_ VGND VGND VPWR VPWR _10371_ sky130_fd_sc_hd__mux2_1
X_21596_ _08514_ _08846_ VGND VGND VPWR VPWR _08847_ sky130_fd_sc_hd__or2_1
XFILLER_0_149_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26123_ _11371_ VGND VGND VPWR VPWR _11397_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_10_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20547_ _06606_ VGND VGND VPWR VPWR _07838_ sky130_fd_sc_hd__buf_8
XFILLER_0_172_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_963 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26054_ _11086_ _11351_ VGND VGND VPWR VPWR _11356_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23138__814 clknet_1_1__leaf__10106_ VGND VGND VPWR VPWR net940 sky130_fd_sc_hd__inv_2
XFILLER_0_127_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20478_ datamem.data_ram\[54\]\[20\] _06743_ _06820_ datamem.data_ram\[48\]\[20\]
+ VGND VGND VPWR VPWR _07770_ sky130_fd_sc_hd__o22a_1
XFILLER_0_104_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25005_ _10723_ VGND VGND VPWR VPWR _02571_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22217_ _09382_ VGND VGND VPWR VPWR _09383_ sky130_fd_sc_hd__clkbuf_4
X_23197_ _10119_ VGND VGND VPWR VPWR _01367_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22148_ _09276_ net3950 net62 VGND VGND VPWR VPWR _09344_ sky130_fd_sc_hd__mux2_1
X_29813_ net191 _01548_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[1\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26956_ _11833_ _11854_ VGND VGND VPWR VPWR _11860_ sky130_fd_sc_hd__and2_1
X_14970_ _13370_ _13472_ _13292_ _13419_ VGND VGND VPWR VPWR _13519_ sky130_fd_sc_hd__a211o_1
X_22079_ rvcpu.dp.plem.MemWriteM rvcpu.dp.plem.ALUResultM\[0\] _06911_ net117 VGND
+ VGND VPWR VPWR _09293_ sky130_fd_sc_hd__and4_2
X_29744_ net1090 _01479_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[21\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_25907_ net1840 _11263_ VGND VGND VPWR VPWR _11272_ sky130_fd_sc_hd__or2_1
X_29675_ net1021 _01410_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[23\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26887_ _11803_ _11810_ VGND VGND VPWR VPWR _11816_ sky130_fd_sc_hd__and2_1
XFILLER_0_92_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28626_ _12809_ VGND VGND VPWR VPWR _04106_ sky130_fd_sc_hd__clkbuf_1
X_16640_ _04539_ VGND VGND VPWR VPWR _04562_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_215_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25838_ rvcpu.dp.pcreg.q\[23\] _11213_ rvcpu.dp.pcreg.q\[24\] VGND VGND VPWR VPWR
+ _11222_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_187_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_214_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23110__788 clknet_1_1__leaf__10104_ VGND VGND VPWR VPWR net914 sky130_fd_sc_hd__inv_2
XFILLER_0_186_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16571_ _04502_ VGND VGND VPWR VPWR _04525_ sky130_fd_sc_hd__clkbuf_4
X_28557_ _12772_ VGND VGND VPWR VPWR _04074_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25769_ _13538_ _11165_ VGND VGND VPWR VPWR _11168_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_54_clk clknet_5_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_54_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_198_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18310_ _05674_ VGND VGND VPWR VPWR _05675_ sky130_fd_sc_hd__buf_2
XFILLER_0_85_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15522_ _13893_ _13959_ _13315_ VGND VGND VPWR VPWR _14049_ sky130_fd_sc_hd__a21o_1
X_27508_ _12185_ VGND VGND VPWR VPWR _03612_ sky130_fd_sc_hd__clkbuf_1
X_19290_ _06585_ rvcpu.dp.plem.ALUResultM\[1\] VGND VGND VPWR VPWR _06586_ sky130_fd_sc_hd__nand2_2
XFILLER_0_85_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_191_5075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28488_ _12727_ net1702 _12723_ _12728_ VGND VGND VPWR VPWR _04049_ sky130_fd_sc_hd__a31o_1
XFILLER_0_31_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23757__346 clknet_1_0__leaf__10201_ VGND VGND VPWR VPWR net472 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_191_5086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_195_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18241_ rvcpu.dp.plde.RD1E\[10\] _05267_ _05271_ _13247_ _05411_ VGND VGND VPWR VPWR
+ _05606_ sky130_fd_sc_hd__a221oi_4
X_15453_ _13514_ _13981_ _13982_ VGND VGND VPWR VPWR _13983_ sky130_fd_sc_hd__a21oi_1
X_27439_ _09272_ VGND VGND VPWR VPWR _12145_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_72_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_210_1268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18172_ _05535_ _05536_ VGND VGND VPWR VPWR _05537_ sky130_fd_sc_hd__nor2_2
X_30450_ net788 _02185_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[29\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_15384_ _13904_ _13908_ _13917_ VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__a21oi_1
XFILLER_0_182_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17123_ _04818_ VGND VGND VPWR VPWR _01477_ sky130_fd_sc_hd__clkbuf_1
X_29109_ _09275_ net2529 _13067_ VGND VGND VPWR VPWR _13070_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30381_ clknet_leaf_267_clk _02116_ VGND VGND VPWR VPWR datamem.data_ram\[58\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32120_ clknet_leaf_83_clk _03542_ VGND VGND VPWR VPWR datamem.data_ram\[0\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_150_4093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold509 datamem.data_ram\[12\]\[5\] VGND VGND VPWR VPWR net1659 sky130_fd_sc_hd__dlygate4sd3_1
X_17054_ net2671 _14468_ _04779_ VGND VGND VPWR VPWR _04782_ sky130_fd_sc_hd__mux2_1
XFILLER_0_204_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_204_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16005_ _14340_ VGND VGND VPWR VPWR _02025_ sky130_fd_sc_hd__clkbuf_1
X_32051_ clknet_leaf_127_clk _03473_ VGND VGND VPWR VPWR datamem.data_ram\[30\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_206_5428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_206_5439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31002_ clknet_leaf_101_clk _02737_ VGND VGND VPWR VPWR datamem.data_ram\[22\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_163_4410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17956_ _13240_ rvcpu.dp.plde.RD2E\[12\] _05194_ VGND VGND VPWR VPWR _05328_ sky130_fd_sc_hd__mux2_1
XFILLER_0_225_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1209 rvcpu.dp.rf.reg_file_arr\[7\]\[18\] VGND VGND VPWR VPWR net2359 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16907_ _04703_ VGND VGND VPWR VPWR _01586_ sky130_fd_sc_hd__clkbuf_1
X_32953_ clknet_leaf_99_clk _04375_ VGND VGND VPWR VPWR datamem.data_ram\[6\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_17887_ rvcpu.dp.plde.Rs1E\[4\] _13176_ VGND VGND VPWR VPWR _05260_ sky130_fd_sc_hd__or2b_1
XFILLER_0_174_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31904_ _04446_ net119 VGND VGND VPWR VPWR datamem.rd_data_mem\[9\] sky130_fd_sc_hd__dlxtn_1
X_19626_ rvcpu.dp.plem.ALUResultM\[4\] _06640_ VGND VGND VPWR VPWR _06922_ sky130_fd_sc_hd__nand2_8
X_16838_ net2381 _14457_ _04659_ VGND VGND VPWR VPWR _04667_ sky130_fd_sc_hd__mux2_1
X_32884_ clknet_leaf_287_clk _04306_ VGND VGND VPWR VPWR datamem.data_ram\[10\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_24137__642 clknet_1_0__leaf__10261_ VGND VGND VPWR VPWR net768 sky130_fd_sc_hd__inv_2
X_23543__168 clknet_1_0__leaf__10173_ VGND VGND VPWR VPWR net294 sky130_fd_sc_hd__inv_2
XFILLER_0_215_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_220_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16769_ _04630_ VGND VGND VPWR VPWR _01659_ sky130_fd_sc_hd__clkbuf_1
X_19557_ datamem.data_ram\[11\]\[24\] _06829_ _06848_ _06852_ VGND VGND VPWR VPWR
+ _06853_ sky130_fd_sc_hd__o211a_1
X_31835_ clknet_leaf_234_clk _03289_ VGND VGND VPWR VPWR datamem.data_ram\[3\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_45_clk clknet_5_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_45_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_87_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_4258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23085__765 clknet_1_1__leaf__10102_ VGND VGND VPWR VPWR net891 sky130_fd_sc_hd__inv_2
XFILLER_0_220_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18508_ _05382_ _05388_ _05662_ VGND VGND VPWR VPWR _05870_ sky130_fd_sc_hd__mux2_1
X_31766_ clknet_leaf_105_clk _03220_ VGND VGND VPWR VPWR datamem.data_ram\[18\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_4269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19488_ _06670_ VGND VGND VPWR VPWR _06784_ sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_83_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30717_ clknet_leaf_179_clk _02452_ VGND VGND VPWR VPWR datamem.data_ram\[49\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_18439_ _05365_ _05662_ VGND VGND VPWR VPWR _05802_ sky130_fd_sc_hd__nand2_1
X_31697_ clknet_leaf_50_clk _03155_ VGND VGND VPWR VPWR rvcpu.dp.pcreg.q\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21450_ _08532_ _08707_ VGND VGND VPWR VPWR _08708_ sky130_fd_sc_hd__nor2_1
XFILLER_0_145_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30648_ clknet_leaf_189_clk _02383_ VGND VGND VPWR VPWR datamem.data_ram\[51\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20401_ datamem.data_ram\[37\]\[12\] _06815_ _06705_ datamem.data_ram\[39\]\[12\]
+ VGND VGND VPWR VPWR _07693_ sky130_fd_sc_hd__o22a_1
XFILLER_0_181_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21381_ _08627_ _08634_ _08639_ _08641_ VGND VGND VPWR VPWR _08642_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_185_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30579_ clknet_leaf_177_clk _02314_ VGND VGND VPWR VPWR datamem.data_ram\[54\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_116_3276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_3287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_92_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20332_ datamem.data_ram\[42\]\[4\] _06989_ _06990_ datamem.data_ram\[40\]\[4\] VGND
+ VGND VPWR VPWR _07624_ sky130_fd_sc_hd__a22o_1
XFILLER_0_141_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_92_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32318_ clknet_leaf_230_clk _03740_ VGND VGND VPWR VPWR datamem.data_ram\[31\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_187_4977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_187_4988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput18 net18 VGND VGND VPWR VPWR Instr[24] sky130_fd_sc_hd__buf_2
X_20263_ datamem.data_ram\[48\]\[19\] _06698_ _06658_ datamem.data_ram\[49\]\[19\]
+ _07555_ VGND VGND VPWR VPWR _07556_ sky130_fd_sc_hd__o221a_1
X_32249_ clknet_leaf_168_clk _03671_ VGND VGND VPWR VPWR datamem.data_ram\[34\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput29 net29 VGND VGND VPWR VPWR Instr[5] sky130_fd_sc_hd__buf_2
X_22002_ _09226_ _09229_ _09231_ VGND VGND VPWR VPWR _09232_ sky130_fd_sc_hd__a21oi_4
Xhold3101 datamem.data_ram\[49\]\[26\] VGND VGND VPWR VPWR net4251 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3112 rvcpu.dp.rf.reg_file_arr\[25\]\[3\] VGND VGND VPWR VPWR net4262 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3123 rvcpu.dp.rf.reg_file_arr\[15\]\[31\] VGND VGND VPWR VPWR net4273 sky130_fd_sc_hd__dlygate4sd3_1
X_20194_ datamem.data_ram\[45\]\[11\] _06865_ _07483_ _07486_ VGND VGND VPWR VPWR
+ _07487_ sky130_fd_sc_hd__o211a_1
Xhold3134 rvcpu.dp.rf.reg_file_arr\[26\]\[2\] VGND VGND VPWR VPWR net4284 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2400 datamem.data_ram\[51\]\[22\] VGND VGND VPWR VPWR net3550 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3145 rvcpu.c.ad.funct7b5 VGND VGND VPWR VPWR net4295 sky130_fd_sc_hd__dlygate4sd3_1
X_26810_ _11767_ net1453 _11761_ _11769_ VGND VGND VPWR VPWR _03330_ sky130_fd_sc_hd__a31o_1
Xhold3156 datamem.data_ram\[55\]\[18\] VGND VGND VPWR VPWR net4306 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2411 datamem.data_ram\[10\]\[24\] VGND VGND VPWR VPWR net3561 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_51_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2422 datamem.data_ram\[0\]\[29\] VGND VGND VPWR VPWR net3572 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3167 datamem.data_ram\[63\]\[8\] VGND VGND VPWR VPWR net4317 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27790_ _12125_ net3029 _12336_ VGND VGND VPWR VPWR _12337_ sky130_fd_sc_hd__mux2_1
Xhold3178 datamem.data_ram\[21\]\[22\] VGND VGND VPWR VPWR net4328 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2433 datamem.data_ram\[8\]\[25\] VGND VGND VPWR VPWR net3583 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2444 datamem.data_ram\[0\]\[11\] VGND VGND VPWR VPWR net3594 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3189 rvcpu.dp.rf.reg_file_arr\[0\]\[10\] VGND VGND VPWR VPWR net4339 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1710 datamem.data_ram\[61\]\[28\] VGND VGND VPWR VPWR net2860 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2455 rvcpu.dp.rf.reg_file_arr\[30\]\[3\] VGND VGND VPWR VPWR net3605 sky130_fd_sc_hd__dlygate4sd3_1
X_26741_ _11700_ net1740 _11724_ _11728_ VGND VGND VPWR VPWR _03302_ sky130_fd_sc_hd__a31o_1
XFILLER_0_215_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_146_3995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1721 rvcpu.dp.rf.reg_file_arr\[17\]\[2\] VGND VGND VPWR VPWR net2871 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2466 datamem.data_ram\[25\]\[31\] VGND VGND VPWR VPWR net3616 sky130_fd_sc_hd__dlygate4sd3_1
X_23953_ _10230_ VGND VGND VPWR VPWR _02012_ sky130_fd_sc_hd__clkbuf_1
Xhold1732 rvcpu.dp.rf.reg_file_arr\[26\]\[10\] VGND VGND VPWR VPWR net2882 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2477 datamem.data_ram\[63\]\[25\] VGND VGND VPWR VPWR net3627 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1743 datamem.data_ram\[38\]\[24\] VGND VGND VPWR VPWR net2893 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2488 datamem.data_ram\[41\]\[11\] VGND VGND VPWR VPWR net3638 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2499 datamem.data_ram\[8\]\[11\] VGND VGND VPWR VPWR net3649 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1754 rvcpu.dp.rf.reg_file_arr\[2\]\[0\] VGND VGND VPWR VPWR net2904 sky130_fd_sc_hd__dlygate4sd3_1
X_29460_ net822 _01195_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[30\]\[31\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_4_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1765 rvcpu.dp.rf.reg_file_arr\[21\]\[29\] VGND VGND VPWR VPWR net2915 sky130_fd_sc_hd__dlygate4sd3_1
X_22904_ _09452_ _10036_ _10038_ _09795_ VGND VGND VPWR VPWR _10039_ sky130_fd_sc_hd__a211o_1
Xclkbuf_1_1__f__10241_ clknet_0__10241_ VGND VGND VPWR VPWR clknet_1_1__leaf__10241_
+ sky130_fd_sc_hd__clkbuf_16
X_26672_ _11687_ _11677_ VGND VGND VPWR VPWR _11688_ sky130_fd_sc_hd__and2_1
Xhold1776 datamem.data_ram\[26\]\[22\] VGND VGND VPWR VPWR net2926 sky130_fd_sc_hd__dlygate4sd3_1
X_23884_ clknet_1_1__leaf__10203_ VGND VGND VPWR VPWR _10222_ sky130_fd_sc_hd__buf_1
Xhold1787 rvcpu.dp.rf.reg_file_arr\[30\]\[24\] VGND VGND VPWR VPWR net2937 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1798 datamem.data_ram\[29\]\[13\] VGND VGND VPWR VPWR net2948 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_155_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28411_ _12682_ VGND VGND VPWR VPWR _04018_ sky130_fd_sc_hd__clkbuf_1
X_25623_ _11076_ VGND VGND VPWR VPWR _11077_ sky130_fd_sc_hd__buf_2
XFILLER_0_224_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29391_ clknet_leaf_1_clk _01126_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD2E\[2\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__10172_ clknet_0__10172_ VGND VGND VPWR VPWR clknet_1_1__leaf__10172_
+ sky130_fd_sc_hd__clkbuf_16
X_22835_ rvcpu.dp.rf.reg_file_arr\[24\]\[28\] rvcpu.dp.rf.reg_file_arr\[25\]\[28\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[28\] rvcpu.dp.rf.reg_file_arr\[27\]\[28\] _09385_
+ _09637_ VGND VGND VPWR VPWR _09973_ sky130_fd_sc_hd__mux4_1
XFILLER_0_6_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28342_ _12645_ VGND VGND VPWR VPWR _03986_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_49_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25554_ _11035_ VGND VGND VPWR VPWR _02808_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22766_ _09906_ _09907_ _09380_ VGND VGND VPWR VPWR _09908_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24505_ _10444_ net4431 _10440_ VGND VGND VPWR VPWR _10445_ sky130_fd_sc_hd__mux2_1
X_28273_ _12365_ net3820 _12603_ VGND VGND VPWR VPWR _12608_ sky130_fd_sc_hd__mux2_1
X_21717_ rvcpu.dp.rf.reg_file_arr\[0\]\[17\] rvcpu.dp.rf.reg_file_arr\[1\]\[17\] rvcpu.dp.rf.reg_file_arr\[2\]\[17\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[17\] _08525_ _08528_ VGND VGND VPWR VPWR _08962_
+ sky130_fd_sc_hd__mux4_1
X_25485_ _10073_ _10995_ _10996_ net1308 VGND VGND VPWR VPWR _02778_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_700 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22697_ _09433_ _09842_ _09789_ VGND VGND VPWR VPWR _09843_ sky130_fd_sc_hd__a21o_1
XFILLER_0_87_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27224_ _11972_ _12019_ VGND VGND VPWR VPWR _12024_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24436_ _10326_ VGND VGND VPWR VPWR _10402_ sky130_fd_sc_hd__buf_2
XFILLER_0_137_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21648_ _08695_ _08896_ VGND VGND VPWR VPWR _08897_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27155_ _07808_ _10326_ _11839_ VGND VGND VPWR VPWR _11982_ sky130_fd_sc_hd__or3_1
X_24367_ _10361_ VGND VGND VPWR VPWR _02295_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_80 _06779_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21579_ _08686_ _08830_ _08748_ VGND VGND VPWR VPWR _08831_ sky130_fd_sc_hd__o21ai_1
XANTENNA_91 _06802_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26106_ _11388_ VGND VGND VPWR VPWR _03006_ sky130_fd_sc_hd__clkbuf_1
X_27086_ net1364 _11933_ _11937_ _10041_ VGND VGND VPWR VPWR _03438_ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24298_ _10322_ VGND VGND VPWR VPWR _02265_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_205_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26037_ _11121_ net1602 _11339_ _11345_ VGND VGND VPWR VPWR _02981_ sky130_fd_sc_hd__a31o_1
XFILLER_0_123_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24006__539 clknet_1_1__leaf__10241_ VGND VGND VPWR VPWR net665 sky130_fd_sc_hd__inv_2
XFILLER_0_101_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17810_ _13186_ rvcpu.dp.plde.RD2E\[29\] _05196_ VGND VGND VPWR VPWR _05201_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18790_ _05275_ _05864_ _05943_ VGND VGND VPWR VPWR _06138_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_201_5314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27988_ _12452_ net2291 net76 VGND VGND VPWR VPWR _12453_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_201_5325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17741_ _13260_ net2961 _05140_ VGND VGND VPWR VPWR _05146_ sky130_fd_sc_hd__mux2_1
X_14953_ _13330_ _13452_ _13501_ VGND VGND VPWR VPWR _13502_ sky130_fd_sc_hd__a21o_1
X_26939_ _11835_ _11842_ VGND VGND VPWR VPWR _11850_ sky130_fd_sc_hd__and2_1
X_29727_ net1073 _01462_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[22\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_222_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23462__111 clknet_1_1__leaf__10157_ VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__inv_2
X_17672_ _05109_ VGND VGND VPWR VPWR _01203_ sky130_fd_sc_hd__clkbuf_1
X_14884_ _13431_ _13432_ _13435_ VGND VGND VPWR VPWR _13436_ sky130_fd_sc_hd__a21o_1
X_29658_ net1004 _01393_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[24\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_193_5126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_193_5137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16623_ _04553_ VGND VGND VPWR VPWR _01728_ sky130_fd_sc_hd__clkbuf_1
X_19411_ _06706_ VGND VGND VPWR VPWR _06707_ sky130_fd_sc_hd__buf_6
XFILLER_0_173_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28609_ _12800_ VGND VGND VPWR VPWR _04098_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29589_ net943 _01324_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[26\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23991__525 clknet_1_1__leaf__10240_ VGND VGND VPWR VPWR net651 sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_27_clk clknet_5_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_27_clk sky130_fd_sc_hd__clkbuf_8
Xmax_cap60 _10466_ VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_4
XFILLER_0_58_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap71 _12814_ VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__buf_4
X_31620_ clknet_leaf_66_clk net1203 VGND VGND VPWR VPWR rvcpu.dp.plmw.lAuiPCW\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_19342_ datamem.data_ram\[10\]\[16\] _06613_ _06621_ datamem.data_ram\[12\]\[16\]
+ _06637_ VGND VGND VPWR VPWR _06638_ sky130_fd_sc_hd__o221a_1
X_16554_ _04516_ VGND VGND VPWR VPWR _01768_ sky130_fd_sc_hd__clkbuf_1
Xmax_cap93 _10641_ VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__buf_4
XFILLER_0_58_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_214_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15505_ _13469_ _14024_ _14032_ VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__o21ai_2
XFILLER_0_35_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31551_ clknet_leaf_63_clk datamem.rd_data_mem\[1\] VGND VGND VPWR VPWR rvcpu.dp.plmw.ReadDataW\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19273_ rvcpu.dp.plfd.InstrD\[6\] rvcpu.c.ad.opb5 _06572_ VGND VGND VPWR VPWR _06573_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_14_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16485_ net3471 _14445_ _04478_ VGND VGND VPWR VPWR _04480_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_532 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_4133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23006__711 clknet_1_0__leaf__10085_ VGND VGND VPWR VPWR net837 sky130_fd_sc_hd__inv_2
XFILLER_0_85_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18224_ _05585_ _05586_ _05368_ _05588_ VGND VGND VPWR VPWR _05589_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_152_4144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30502_ clknet_leaf_175_clk _02237_ VGND VGND VPWR VPWR datamem.data_ram\[57\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15436_ _13451_ _13666_ _13872_ _13483_ _13438_ VGND VGND VPWR VPWR _13967_ sky130_fd_sc_hd__a311o_1
XFILLER_0_182_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31482_ clknet_leaf_48_clk rvcpu.dp.lAuiPCE\[8\] VGND VGND VPWR VPWR rvcpu.dp.plem.lAuiPCM\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_152_4155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18155_ _05469_ _05470_ VGND VGND VPWR VPWR _05520_ sky130_fd_sc_hd__or2_1
X_30433_ net771 _02168_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[29\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_15367_ _13343_ _13897_ _13898_ _13899_ _13901_ VGND VGND VPWR VPWR _13902_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_14_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__10261_ clknet_0__10261_ VGND VGND VPWR VPWR clknet_1_0__leaf__10261_
+ sky130_fd_sc_hd__clkbuf_16
X_17106_ _04809_ VGND VGND VPWR VPWR _01485_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18086_ _05338_ _05453_ VGND VGND VPWR VPWR _05454_ sky130_fd_sc_hd__or2_2
XFILLER_0_13_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30364_ net710 _02099_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[3\]\[15\] sky130_fd_sc_hd__dfxtp_1
Xhold306 datamem.data_ram\[17\]\[7\] VGND VGND VPWR VPWR net1456 sky130_fd_sc_hd__dlygate4sd3_1
X_15298_ _13432_ _13322_ _13796_ _13776_ _13370_ VGND VGND VPWR VPWR _13836_ sky130_fd_sc_hd__o311a_1
Xhold317 datamem.data_ram\[57\]\[4\] VGND VGND VPWR VPWR net1467 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32103_ clknet_leaf_114_clk _03525_ VGND VGND VPWR VPWR datamem.data_ram\[23\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold328 datamem.data_ram\[3\]\[2\] VGND VGND VPWR VPWR net1478 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__10192_ clknet_0__10192_ VGND VGND VPWR VPWR clknet_1_0__leaf__10192_
+ sky130_fd_sc_hd__clkbuf_16
Xhold339 datamem.data_ram\[55\]\[3\] VGND VGND VPWR VPWR net1489 sky130_fd_sc_hd__dlygate4sd3_1
X_17037_ net2896 _14451_ _04768_ VGND VGND VPWR VPWR _04773_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_229_5984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_111_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_229_5995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30295_ net641 _02030_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[5\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_111_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_55 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32034_ clknet_leaf_132_clk _03456_ VGND VGND VPWR VPWR datamem.data_ram\[50\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_182_4852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_4863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_4874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23926__482 clknet_1_0__leaf__10226_ VGND VGND VPWR VPWR net608 sky130_fd_sc_hd__inv_2
X_18988_ _05561_ _05644_ VGND VGND VPWR VPWR _06323_ sky130_fd_sc_hd__nand2_1
Xhold1006 rvcpu.dp.rf.reg_file_arr\[19\]\[31\] VGND VGND VPWR VPWR net2156 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1017 rvcpu.dp.rf.reg_file_arr\[5\]\[21\] VGND VGND VPWR VPWR net2167 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_183_Right_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1028 datamem.data_ram\[32\]\[22\] VGND VGND VPWR VPWR net2178 sky130_fd_sc_hd__dlygate4sd3_1
X_17939_ net105 _05310_ VGND VGND VPWR VPWR _05311_ sky130_fd_sc_hd__xnor2_4
Xhold1039 rvcpu.dp.rf.reg_file_arr\[8\]\[13\] VGND VGND VPWR VPWR net2189 sky130_fd_sc_hd__dlygate4sd3_1
X_23625__243 clknet_1_1__leaf__10180_ VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_159_4309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20950_ _06985_ _08197_ _08210_ _08239_ VGND VGND VPWR VPWR _08240_ sky130_fd_sc_hd__a31oi_4
X_32936_ clknet_leaf_146_clk _04358_ VGND VGND VPWR VPWR datamem.data_ram\[7\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_1_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_3870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19609_ datamem.data_ram\[27\]\[8\] _06828_ _06789_ datamem.data_ram\[25\]\[8\] _06904_
+ VGND VGND VPWR VPWR _06905_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_141_3881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20881_ _08169_ _08170_ _07821_ VGND VGND VPWR VPWR _08171_ sky130_fd_sc_hd__mux2_1
X_32867_ clknet_leaf_251_clk _04289_ VGND VGND VPWR VPWR datamem.data_ram\[11\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_18_clk clknet_5_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_18_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_49_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22620_ rvcpu.dp.rf.reg_file_arr\[4\]\[16\] rvcpu.dp.rf.reg_file_arr\[5\]\[16\] rvcpu.dp.rf.reg_file_arr\[6\]\[16\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[16\] _09604_ _09716_ VGND VGND VPWR VPWR _09770_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_81_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31818_ clknet_leaf_103_clk _03272_ VGND VGND VPWR VPWR datamem.data_ram\[9\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_81_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32798_ clknet_leaf_238_clk _04220_ VGND VGND VPWR VPWR datamem.data_ram\[13\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22551_ _09704_ VGND VGND VPWR VPWR _01136_ sky130_fd_sc_hd__clkbuf_1
X_31749_ _04450_ net126 VGND VGND VPWR VPWR rvcpu.ALUControl\[3\] sky130_fd_sc_hd__dlxtn_1
XTAP_TAPCELL_ROW_118_3316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_3327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23360__996 clknet_1_1__leaf__10138_ VGND VGND VPWR VPWR net1122 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_118_3338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21502_ _08572_ _08757_ VGND VGND VPWR VPWR _08758_ sky130_fd_sc_hd__or2_1
X_25270_ _10076_ _10868_ VGND VGND VPWR VPWR _10877_ sky130_fd_sc_hd__and2_1
XFILLER_0_91_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22482_ _09636_ _09638_ VGND VGND VPWR VPWR _09639_ sky130_fd_sc_hd__nor2_1
XFILLER_0_228_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24221_ _10281_ VGND VGND VPWR VPWR _02229_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21433_ _08523_ VGND VGND VPWR VPWR _08692_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21364_ _08546_ _08564_ _08577_ _08625_ VGND VGND VPWR VPWR _01028_ sky130_fd_sc_hd__o31a_1
XFILLER_0_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20315_ datamem.data_ram\[13\]\[4\] _06969_ _06976_ datamem.data_ram\[12\]\[4\] _06776_
+ VGND VGND VPWR VPWR _07607_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_1058 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28960_ _07791_ _10042_ _10918_ VGND VGND VPWR VPWR _12987_ sky130_fd_sc_hd__or3_1
XFILLER_0_141_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24083_ _10253_ VGND VGND VPWR VPWR _02119_ sky130_fd_sc_hd__clkbuf_1
X_21295_ rvcpu.dp.plfd.InstrD\[18\] VGND VGND VPWR VPWR _08557_ sky130_fd_sc_hd__inv_2
Xhold840 rvcpu.dp.rf.reg_file_arr\[11\]\[16\] VGND VGND VPWR VPWR net1990 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_820 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold851 datamem.data_ram\[28\]\[31\] VGND VGND VPWR VPWR net2001 sky130_fd_sc_hd__dlygate4sd3_1
Xhold862 rvcpu.dp.rf.reg_file_arr\[2\]\[24\] VGND VGND VPWR VPWR net2012 sky130_fd_sc_hd__dlygate4sd3_1
X_20246_ datamem.data_ram\[58\]\[3\] _07136_ _07535_ _07538_ VGND VGND VPWR VPWR _07539_
+ sky130_fd_sc_hd__a211o_1
X_27911_ _12149_ net2488 net47 VGND VGND VPWR VPWR _12407_ sky130_fd_sc_hd__mux2_1
X_23786__372 clknet_1_0__leaf__10204_ VGND VGND VPWR VPWR net498 sky130_fd_sc_hd__inv_2
Xhold873 rvcpu.dp.rf.reg_file_arr\[6\]\[8\] VGND VGND VPWR VPWR net2023 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold884 rvcpu.dp.rf.reg_file_arr\[4\]\[19\] VGND VGND VPWR VPWR net2034 sky130_fd_sc_hd__dlygate4sd3_1
X_28891_ _12178_ _11020_ _12886_ VGND VGND VPWR VPWR _12950_ sky130_fd_sc_hd__a21oi_1
Xhold895 rvcpu.dp.rf.reg_file_arr\[5\]\[12\] VGND VGND VPWR VPWR net2045 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_228_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27842_ _12367_ net3934 _12357_ VGND VGND VPWR VPWR _12368_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20177_ _06680_ _07467_ _07469_ VGND VGND VPWR VPWR _07470_ sky130_fd_sc_hd__and3_1
XFILLER_0_216_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2230 datamem.data_ram\[61\]\[30\] VGND VGND VPWR VPWR net3380 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2241 datamem.data_ram\[51\]\[20\] VGND VGND VPWR VPWR net3391 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2252 datamem.data_ram\[54\]\[15\] VGND VGND VPWR VPWR net3402 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27773_ _12327_ VGND VGND VPWR VPWR _03735_ sky130_fd_sc_hd__clkbuf_1
Xhold2263 rvcpu.dp.rf.reg_file_arr\[16\]\[19\] VGND VGND VPWR VPWR net3413 sky130_fd_sc_hd__dlygate4sd3_1
X_24985_ _10478_ net3116 _10706_ VGND VGND VPWR VPWR _10713_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_150_Right_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2274 rvcpu.dp.rf.reg_file_arr\[16\]\[5\] VGND VGND VPWR VPWR net3424 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1540 datamem.data_ram\[9\]\[23\] VGND VGND VPWR VPWR net2690 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2285 datamem.data_ram\[23\]\[25\] VGND VGND VPWR VPWR net3435 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1551 datamem.data_ram\[3\]\[16\] VGND VGND VPWR VPWR net2701 sky130_fd_sc_hd__dlygate4sd3_1
X_26724_ _10758_ net3302 _11714_ VGND VGND VPWR VPWR _11718_ sky130_fd_sc_hd__mux2_1
Xhold2296 rvcpu.dp.rf.reg_file_arr\[14\]\[25\] VGND VGND VPWR VPWR net3446 sky130_fd_sc_hd__dlygate4sd3_1
X_29512_ net874 _01247_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[28\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1562 rvcpu.dp.rf.reg_file_arr\[21\]\[14\] VGND VGND VPWR VPWR net2712 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1573 rvcpu.dp.rf.reg_file_arr\[16\]\[0\] VGND VGND VPWR VPWR net2723 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_1300 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1584 rvcpu.dp.rf.reg_file_arr\[12\]\[19\] VGND VGND VPWR VPWR net2734 sky130_fd_sc_hd__dlygate4sd3_1
X_29443_ net805 _01178_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[30\]\[14\] sky130_fd_sc_hd__dfxtp_1
Xhold1595 datamem.data_ram\[13\]\[15\] VGND VGND VPWR VPWR net2745 sky130_fd_sc_hd__dlygate4sd3_1
X_26655_ _10047_ VGND VGND VPWR VPWR _11676_ sky130_fd_sc_hd__buf_2
Xclkbuf_1_1__f__10224_ clknet_0__10224_ VGND VGND VPWR VPWR clknet_1_1__leaf__10224_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_200_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_212_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25606_ _11067_ VGND VGND VPWR VPWR _02828_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_196_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29374_ clknet_leaf_140_clk _01109_ VGND VGND VPWR VPWR datamem.data_ram\[60\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_22818_ rvcpu.dp.rf.reg_file_arr\[16\]\[27\] rvcpu.dp.rf.reg_file_arr\[17\]\[27\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[27\] rvcpu.dp.rf.reg_file_arr\[19\]\[27\] _09406_
+ _09408_ VGND VGND VPWR VPWR _09957_ sky130_fd_sc_hd__mux4_1
X_26586_ _11638_ VGND VGND VPWR VPWR _11639_ sky130_fd_sc_hd__buf_2
XFILLER_0_39_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__10155_ clknet_0__10155_ VGND VGND VPWR VPWR clknet_1_1__leaf__10155_
+ sky130_fd_sc_hd__clkbuf_16
X_28325_ _12636_ VGND VGND VPWR VPWR _03978_ sky130_fd_sc_hd__clkbuf_1
X_25537_ _11026_ VGND VGND VPWR VPWR _02800_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22749_ _09510_ _09885_ _09887_ _09891_ _09525_ VGND VGND VPWR VPWR _09892_ sky130_fd_sc_hd__a311o_1
Xclkbuf_1_1__f__10086_ clknet_0__10086_ VGND VGND VPWR VPWR clknet_1_1__leaf__10086_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_165_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28256_ _12458_ net3551 net44 VGND VGND VPWR VPWR _12598_ sky130_fd_sc_hd__mux2_1
X_16270_ net3066 _14436_ _14489_ VGND VGND VPWR VPWR _14497_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25468_ _10067_ _10985_ VGND VGND VPWR VPWR _10990_ sky130_fd_sc_hd__and2_1
XFILLER_0_180_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27207_ _12005_ net1474 _12007_ _12013_ VGND VGND VPWR VPWR _03483_ sky130_fd_sc_hd__a31o_1
X_15221_ _13466_ _13761_ VGND VGND VPWR VPWR _13762_ sky130_fd_sc_hd__and2_1
XFILLER_0_168_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24419_ _10390_ datamem.data_ram\[53\]\[10\] _10386_ VGND VGND VPWR VPWR _10391_
+ sky130_fd_sc_hd__mux2_1
X_28187_ _12441_ net4121 _12555_ VGND VGND VPWR VPWR _12561_ sky130_fd_sc_hd__mux2_1
X_25399_ _10055_ VGND VGND VPWR VPWR _10954_ sky130_fd_sc_hd__buf_2
XFILLER_0_191_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15152_ _13447_ _13434_ VGND VGND VPWR VPWR _13696_ sky130_fd_sc_hd__nor2_1
X_27138_ _11970_ _11966_ VGND VGND VPWR VPWR _11971_ sky130_fd_sc_hd__and2_1
XFILLER_0_50_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_270 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27069_ _11919_ net1658 _11923_ _11927_ VGND VGND VPWR VPWR _03431_ sky130_fd_sc_hd__a31o_1
X_15083_ _13628_ _13359_ _13608_ VGND VGND VPWR VPWR _13629_ sky130_fd_sc_hd__o21a_1
X_19960_ datamem.data_ram\[5\]\[18\] _06663_ _06784_ datamem.data_ram\[7\]\[18\] VGND
+ VGND VPWR VPWR _07254_ sky130_fd_sc_hd__o22a_1
XFILLER_0_120_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18911_ _05619_ _05620_ _05629_ VGND VGND VPWR VPWR _06251_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30080_ net442 _01815_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[11\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19891_ datamem.data_ram\[22\]\[17\] _06630_ _06701_ datamem.data_ram\[17\]\[17\]
+ _07185_ VGND VGND VPWR VPWR _07186_ sky130_fd_sc_hd__o221a_1
XFILLER_0_129_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23036__737 clknet_1_1__leaf__10089_ VGND VGND VPWR VPWR net863 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_224_5870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18842_ _05990_ _06058_ _06185_ _06109_ _06186_ VGND VGND VPWR VPWR _06187_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_224_5881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23116__794 clknet_1_0__leaf__10104_ VGND VGND VPWR VPWR net920 sky130_fd_sc_hd__inv_2
X_18773_ _05318_ _05612_ _06104_ _06121_ _05655_ VGND VGND VPWR VPWR _06122_ sky130_fd_sc_hd__a311oi_1
X_15985_ net1941 _13235_ _14322_ VGND VGND VPWR VPWR _14330_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_220_5767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_220_5778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14936_ _13481_ _13483_ _13484_ VGND VGND VPWR VPWR _13485_ sky130_fd_sc_hd__or3b_1
X_17724_ _13235_ net1946 _05129_ VGND VGND VPWR VPWR _05137_ sky130_fd_sc_hd__mux2_1
X_30982_ clknet_leaf_94_clk _02717_ VGND VGND VPWR VPWR datamem.data_ram\[39\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24182__23 clknet_1_0__leaf__10265_ VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__inv_2
XFILLER_0_199_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32721_ clknet_leaf_244_clk _04143_ VGND VGND VPWR VPWR datamem.data_ram\[16\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_14867_ _13371_ VGND VGND VPWR VPWR _13419_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_199_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17655_ _05100_ VGND VGND VPWR VPWR _01211_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_19_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Left_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16606_ _04544_ VGND VGND VPWR VPWR _01736_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32652_ clknet_leaf_244_clk _04074_ VGND VGND VPWR VPWR datamem.data_ram\[19\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_17586_ _13232_ net3128 _05057_ VGND VGND VPWR VPWR _05064_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14798_ _13349_ _13350_ VGND VGND VPWR VPWR _13351_ sky130_fd_sc_hd__or2_1
XFILLER_0_212_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31603_ clknet_leaf_45_clk net1168 VGND VGND VPWR VPWR rvcpu.dp.plmw.PCPlus4W\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_19325_ _06620_ VGND VGND VPWR VPWR _06621_ sky130_fd_sc_hd__buf_4
XFILLER_0_128_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16537_ _04507_ VGND VGND VPWR VPWR _01776_ sky130_fd_sc_hd__clkbuf_1
X_32583_ clknet_leaf_184_clk _04005_ VGND VGND VPWR VPWR datamem.data_ram\[21\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19256_ _06558_ rvcpu.dp.plde.ImmExtE\[30\] rvcpu.dp.plde.luiE VGND VGND VPWR VPWR
+ _06559_ sky130_fd_sc_hd__mux2_1
X_31534_ clknet_leaf_24_clk net1217 VGND VGND VPWR VPWR rvcpu.dp.plem.PCPlus4M\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_16468_ net3917 _14428_ _04467_ VGND VGND VPWR VPWR _04471_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15419_ _13459_ _13526_ _13509_ _13950_ VGND VGND VPWR VPWR _13951_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_171_4597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18207_ _05497_ _05569_ _05571_ VGND VGND VPWR VPWR _05572_ sky130_fd_sc_hd__o21ai_1
X_19187_ _06497_ _06498_ VGND VGND VPWR VPWR _06499_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_170_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31465_ clknet_leaf_5_clk rvcpu.dp.SrcBFW_Mux.y\[23\] VGND VGND VPWR VPWR rvcpu.dp.plem.WriteDataM\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_113_3202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16399_ _14565_ VGND VGND VPWR VPWR _01840_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_113_3213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18138_ _05502_ _05503_ VGND VGND VPWR VPWR _05504_ sky130_fd_sc_hd__nor2_2
XFILLER_0_53_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30416_ net754 _02151_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[31\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_31396_ clknet_leaf_50_clk _03099_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCE\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_184_4903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold103 rvcpu.dp.plem.ALUResultM\[17\] VGND VGND VPWR VPWR net1253 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__10244_ clknet_0__10244_ VGND VGND VPWR VPWR clknet_1_0__leaf__10244_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_130_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Left_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_184_4914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold114 rvcpu.dp.plem.ALUResultM\[15\] VGND VGND VPWR VPWR net1264 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold125 rvcpu.dp.plem.ALUResultM\[26\] VGND VGND VPWR VPWR net1275 sky130_fd_sc_hd__dlygate4sd3_1
X_18069_ rvcpu.dp.plde.RD1E\[13\] _05266_ _05270_ _13237_ _05319_ VGND VGND VPWR VPWR
+ _05437_ sky130_fd_sc_hd__a221oi_4
X_30347_ net693 _02082_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[4\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold136 rvcpu.dp.plem.ALUResultM\[11\] VGND VGND VPWR VPWR net1286 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_7_clk clknet_5_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_223_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold147 datamem.data_ram\[45\]\[5\] VGND VGND VPWR VPWR net1297 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold158 datamem.data_ram\[41\]\[6\] VGND VGND VPWR VPWR net1308 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__10175_ clknet_0__10175_ VGND VGND VPWR VPWR clknet_1_0__leaf__10175_
+ sky130_fd_sc_hd__clkbuf_16
X_20100_ datamem.data_ram\[0\]\[10\] _06837_ _07392_ _07393_ VGND VGND VPWR VPWR _07394_
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_74_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold169 datamem.data_ram\[47\]\[6\] VGND VGND VPWR VPWR net1319 sky130_fd_sc_hd__dlygate4sd3_1
X_21080_ _08355_ _08361_ _08368_ _06733_ VGND VGND VPWR VPWR _08369_ sky130_fd_sc_hd__a211o_1
X_30278_ clknet_leaf_141_clk _02013_ VGND VGND VPWR VPWR datamem.data_ram\[58\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_223_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23469__117 clknet_1_0__leaf__10158_ VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__inv_2
X_32017_ clknet_leaf_129_clk _03439_ VGND VGND VPWR VPWR datamem.data_ram\[51\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_20031_ datamem.data_ram\[26\]\[26\] _06609_ _06632_ datamem.data_ram\[27\]\[26\]
+ VGND VGND VPWR VPWR _07325_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_6_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23549__174 clknet_1_1__leaf__10173_ VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_143_3932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24770_ _10476_ net4197 _10589_ VGND VGND VPWR VPWR _10595_ sky130_fd_sc_hd__mux2_1
XFILLER_0_213_539 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21982_ _09212_ VGND VGND VPWR VPWR _01059_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_206_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32919_ clknet_leaf_157_clk _04341_ VGND VGND VPWR VPWR datamem.data_ram\[0\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_20933_ datamem.data_ram\[32\]\[22\] _06973_ _08220_ _07868_ _08222_ VGND VGND VPWR
+ VPWR _08223_ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_221_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26440_ _11545_ rvcpu.ALUResultE\[19\] VGND VGND VPWR VPWR _11571_ sky130_fd_sc_hd__and2_1
XFILLER_0_179_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20864_ datamem.data_ram\[36\]\[14\] _07862_ _06934_ datamem.data_ram\[32\]\[14\]
+ VGND VGND VPWR VPWR _08154_ sky130_fd_sc_hd__o22a_1
XFILLER_0_178_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_102_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22603_ _09622_ _09751_ _09753_ VGND VGND VPWR VPWR _09754_ sky130_fd_sc_hd__a21o_1
X_26371_ _11064_ _11511_ VGND VGND VPWR VPWR _11520_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23583_ clknet_1_0__leaf__10172_ VGND VGND VPWR VPWR _10177_ sky130_fd_sc_hd__buf_1
XFILLER_0_7_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20795_ datamem.data_ram\[36\]\[30\] datamem.data_ram\[37\]\[30\] _07835_ VGND VGND
+ VPWR VPWR _08085_ sky130_fd_sc_hd__mux2_1
XFILLER_0_187_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28110_ _12520_ VGND VGND VPWR VPWR _03879_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_187_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25322_ _10824_ net2271 _10899_ VGND VGND VPWR VPWR _10906_ sky130_fd_sc_hd__mux2_1
X_22534_ rvcpu.dp.rf.reg_file_arr\[16\]\[12\] rvcpu.dp.rf.reg_file_arr\[17\]\[12\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[12\] rvcpu.dp.rf.reg_file_arr\[19\]\[12\] _09384_
+ _09577_ VGND VGND VPWR VPWR _09688_ sky130_fd_sc_hd__mux4_1
X_29090_ _09305_ net2730 net40 VGND VGND VPWR VPWR _13060_ sky130_fd_sc_hd__mux2_1
XFILLER_0_221_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28041_ _12447_ net3937 net96 VGND VGND VPWR VPWR _12484_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25253_ _10866_ VGND VGND VPWR VPWR _10867_ sky130_fd_sc_hd__buf_2
X_22465_ rvcpu.dp.rf.reg_file_arr\[0\]\[8\] rvcpu.dp.rf.reg_file_arr\[1\]\[8\] rvcpu.dp.rf.reg_file_arr\[2\]\[8\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[8\] _09417_ _09585_ VGND VGND VPWR VPWR _09623_ sky130_fd_sc_hd__mux4_1
X_24204_ _10272_ VGND VGND VPWR VPWR _02221_ sky130_fd_sc_hd__clkbuf_1
X_21416_ _08673_ _08674_ VGND VGND VPWR VPWR _08675_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25184_ _10724_ net3431 net57 VGND VGND VPWR VPWR _10830_ sky130_fd_sc_hd__mux2_1
X_22396_ rvcpu.dp.rf.reg_file_arr\[16\]\[5\] rvcpu.dp.rf.reg_file_arr\[17\]\[5\] rvcpu.dp.rf.reg_file_arr\[18\]\[5\]
+ rvcpu.dp.rf.reg_file_arr\[19\]\[5\] _09445_ _09447_ VGND VGND VPWR VPWR _09557_
+ sky130_fd_sc_hd__mux4_1
X_21347_ rvcpu.ALUResultE\[22\] rvcpu.ALUResultE\[25\] rvcpu.ALUResultE\[26\] rvcpu.ALUResultE\[28\]
+ VGND VGND VPWR VPWR _08609_ sky130_fd_sc_hd__or4_1
X_29992_ net362 _01727_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[14\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_198_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_202_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28943_ _09350_ _11020_ _12977_ VGND VGND VPWR VPWR _12978_ sky130_fd_sc_hd__a21oi_2
Xhold670 datamem.data_ram\[8\]\[6\] VGND VGND VPWR VPWR net1820 sky130_fd_sc_hd__dlygate4sd3_1
X_21278_ rvcpu.dp.plfd.InstrD\[17\] VGND VGND VPWR VPWR _08540_ sky130_fd_sc_hd__buf_4
Xhold681 datamem.data_ram\[16\]\[5\] VGND VGND VPWR VPWR net1831 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold692 datamem.data_ram\[34\]\[3\] VGND VGND VPWR VPWR net1842 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20229_ datamem.data_ram\[14\]\[3\] _07127_ _07518_ _07521_ VGND VGND VPWR VPWR _07522_
+ sky130_fd_sc_hd__a211o_1
X_28874_ _12178_ _10960_ _12886_ VGND VGND VPWR VPWR _12941_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_198_1277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27825_ _10500_ VGND VGND VPWR VPWR _12356_ sky130_fd_sc_hd__buf_6
Xhold2060 datamem.data_ram\[46\]\[15\] VGND VGND VPWR VPWR net3210 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2071 datamem.data_ram\[9\]\[29\] VGND VGND VPWR VPWR net3221 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2082 datamem.data_ram\[31\]\[17\] VGND VGND VPWR VPWR net3232 sky130_fd_sc_hd__dlygate4sd3_1
X_15770_ _14214_ VGND VGND VPWR VPWR _02142_ sky130_fd_sc_hd__clkbuf_1
X_24968_ _10703_ VGND VGND VPWR VPWR _02554_ sky130_fd_sc_hd__clkbuf_1
Xhold2093 rvcpu.dp.rf.reg_file_arr\[13\]\[6\] VGND VGND VPWR VPWR net3243 sky130_fd_sc_hd__dlygate4sd3_1
X_27756_ _12145_ net2808 _12316_ VGND VGND VPWR VPWR _12318_ sky130_fd_sc_hd__mux2_1
Xhold1370 rvcpu.dp.rf.reg_file_arr\[23\]\[4\] VGND VGND VPWR VPWR net2520 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1381 rvcpu.dp.rf.reg_file_arr\[8\]\[23\] VGND VGND VPWR VPWR net2531 sky130_fd_sc_hd__dlygate4sd3_1
X_14721_ net3655 _13275_ _13180_ VGND VGND VPWR VPWR _13276_ sky130_fd_sc_hd__mux2_1
X_26707_ _11708_ VGND VGND VPWR VPWR _03288_ sky130_fd_sc_hd__clkbuf_1
X_27687_ _12281_ VGND VGND VPWR VPWR _03695_ sky130_fd_sc_hd__clkbuf_1
Xhold1392 datamem.data_ram\[53\]\[18\] VGND VGND VPWR VPWR net2542 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_419 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24899_ _10666_ VGND VGND VPWR VPWR _02522_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_510 _13216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_200_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_521 _13251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_532 rvcpu.dp.SrcBFW_Mux.y\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17440_ _14154_ net4002 _04985_ VGND VGND VPWR VPWR _04987_ sky130_fd_sc_hd__mux2_1
X_26638_ _11081_ _11663_ VGND VGND VPWR VPWR _11666_ sky130_fd_sc_hd__and2_1
XFILLER_0_196_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29426_ clknet_leaf_98_clk _01161_ VGND VGND VPWR VPWR datamem.data_ram\[5\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14652_ net2246 _13223_ _13214_ VGND VGND VPWR VPWR _13224_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1__f__10207_ clknet_0__10207_ VGND VGND VPWR VPWR clknet_1_1__leaf__10207_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_197_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_543 _06753_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_196_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_554 _07845_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_565 _13254_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0__10238_ _10238_ VGND VGND VPWR VPWR clknet_0__10238_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_71_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17371_ _04950_ VGND VGND VPWR VPWR _01353_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_185_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14583_ rvcpu.dp.plmw.ResultSrcW\[0\] VGND VGND VPWR VPWR _13168_ sky130_fd_sc_hd__clkbuf_8
Xclkbuf_1_1__f__10138_ clknet_0__10138_ VGND VGND VPWR VPWR clknet_1_1__leaf__10138_
+ sky130_fd_sc_hd__clkbuf_16
X_26569_ _10724_ net2414 _11629_ VGND VGND VPWR VPWR _11630_ sky130_fd_sc_hd__mux2_1
X_29357_ clknet_leaf_267_clk _01092_ VGND VGND VPWR VPWR datamem.data_ram\[61\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_211_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19110_ _06421_ _06430_ VGND VGND VPWR VPWR _06431_ sky130_fd_sc_hd__nand2_1
X_16322_ _13177_ _14347_ VGND VGND VPWR VPWR _14524_ sky130_fd_sc_hd__nor2_2
X_28308_ _12627_ VGND VGND VPWR VPWR _03970_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_188_5003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29288_ _13165_ VGND VGND VPWR VPWR _04412_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_188_5014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19041_ _06369_ _06370_ VGND VGND VPWR VPWR _06371_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_153_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28239_ _12441_ net3063 _12583_ VGND VGND VPWR VPWR _12589_ sky130_fd_sc_hd__mux2_1
X_16253_ _14487_ VGND VGND VPWR VPWR _01916_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15204_ _13298_ _13589_ _13616_ VGND VGND VPWR VPWR _13746_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_113_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_680 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31250_ clknet_leaf_21_clk _02953_ VGND VGND VPWR VPWR rvcpu.dp.plfd.InstrD\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16184_ net2346 _14440_ _14422_ VGND VGND VPWR VPWR _14441_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30201_ net555 _01936_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[8\]\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_226_5910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15135_ _13676_ _13679_ _13638_ VGND VGND VPWR VPWR _13680_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_226_5921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31181_ clknet_leaf_38_clk _02884_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCPlus4D\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_147_4021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_147_4032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30132_ net494 _01867_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[10\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15066_ _13572_ _13596_ _13602_ _13612_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__o22a_1
X_19943_ datamem.data_ram\[40\]\[18\] _06778_ _06619_ datamem.data_ram\[44\]\[18\]
+ _07236_ VGND VGND VPWR VPWR _07237_ sky130_fd_sc_hd__o221a_1
XFILLER_0_227_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_222_5818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_222_5829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30063_ net425 _01798_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[12\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19874_ datamem.data_ram\[31\]\[1\] _06927_ _07167_ _07168_ VGND VGND VPWR VPWR _07169_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18825_ _05313_ _05500_ _05506_ _05490_ _05768_ _05769_ VGND VGND VPWR VPWR _06171_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_65_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23997__531 clknet_1_0__leaf__10240_ VGND VGND VPWR VPWR net657 sky130_fd_sc_hd__inv_2
X_18756_ _05436_ _06082_ _05438_ _05333_ VGND VGND VPWR VPWR _06106_ sky130_fd_sc_hd__a31o_1
X_15968_ net2543 _13210_ _14311_ VGND VGND VPWR VPWR _14321_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_106_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17707_ _13210_ net2134 _05118_ VGND VGND VPWR VPWR _05128_ sky130_fd_sc_hd__mux2_1
X_14919_ _13457_ _13461_ _13468_ _13405_ VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_177_4740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18687_ _05419_ _06039_ VGND VGND VPWR VPWR _06041_ sky130_fd_sc_hd__or2_1
XFILLER_0_136_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30965_ clknet_leaf_227_clk _02700_ VGND VGND VPWR VPWR datamem.data_ram\[39\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15899_ _14284_ VGND VGND VPWR VPWR _02075_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_177_4751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32704_ clknet_leaf_181_clk _04126_ VGND VGND VPWR VPWR datamem.data_ram\[17\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17638_ _05091_ VGND VGND VPWR VPWR _01219_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_216_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30896_ clknet_leaf_155_clk _02631_ VGND VGND VPWR VPWR datamem.data_ram\[41\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_173_4637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_4648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32635_ clknet_leaf_255_clk _04057_ VGND VGND VPWR VPWR datamem.data_ram\[1\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_173_4659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17569_ _13207_ net2041 _05046_ VGND VGND VPWR VPWR _05055_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19308_ _06603_ VGND VGND VPWR VPWR _06604_ sky130_fd_sc_hd__buf_4
XFILLER_0_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20580_ _07858_ _07870_ _06603_ VGND VGND VPWR VPWR _07871_ sky130_fd_sc_hd__a21oi_1
X_32566_ clknet_leaf_82_clk _03988_ VGND VGND VPWR VPWR datamem.data_ram\[22\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_31517_ clknet_leaf_51_clk net1230 VGND VGND VPWR VPWR rvcpu.dp.plem.PCPlus4M\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_19239_ _06535_ _06543_ VGND VGND VPWR VPWR _06544_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32497_ clknet_leaf_248_clk _03919_ VGND VGND VPWR VPWR datamem.data_ram\[25\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22250_ _09401_ VGND VGND VPWR VPWR _09416_ sky130_fd_sc_hd__buf_4
XFILLER_0_108_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31448_ clknet_leaf_76_clk rvcpu.dp.SrcBFW_Mux.y\[6\] VGND VGND VPWR VPWR rvcpu.dp.plem.WriteDataM\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_132_3655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_1142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21201_ _08471_ _08482_ VGND VGND VPWR VPWR _08483_ sky130_fd_sc_hd__or2b_1
XFILLER_0_170_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22181_ _09224_ net4160 _09362_ VGND VGND VPWR VPWR _09363_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31379_ clknet_leaf_24_clk _03082_ VGND VGND VPWR VPWR rvcpu.dp.plde.ImmExtE\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_223_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__10227_ clknet_0__10227_ VGND VGND VPWR VPWR clknet_1_0__leaf__10227_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_2_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21132_ _07844_ _08420_ _06599_ VGND VGND VPWR VPWR _08421_ sky130_fd_sc_hd__a21o_1
Xclkbuf_1_0__f__10158_ clknet_0__10158_ VGND VGND VPWR VPWR clknet_1_0__leaf__10158_
+ sky130_fd_sc_hd__clkbuf_16
X_25940_ net1802 _11279_ VGND VGND VPWR VPWR _11292_ sky130_fd_sc_hd__or2_1
X_21063_ _07154_ _08331_ _08338_ _08345_ _08351_ VGND VGND VPWR VPWR _08352_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_35_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22993__699 clknet_1_0__leaf__10084_ VGND VGND VPWR VPWR net825 sky130_fd_sc_hd__inv_2
X_20014_ datamem.data_ram\[53\]\[2\] _06920_ _07306_ _07307_ VGND VGND VPWR VPWR _07308_
+ sky130_fd_sc_hd__a211o_1
Xclkbuf_1_0__f__10089_ clknet_0__10089_ VGND VGND VPWR VPWR clknet_1_0__leaf__10089_
+ sky130_fd_sc_hd__clkbuf_16
X_25871_ _11247_ _11248_ VGND VGND VPWR VPWR _11249_ sky130_fd_sc_hd__nor2_1
X_27610_ _12239_ VGND VGND VPWR VPWR _03660_ sky130_fd_sc_hd__clkbuf_1
X_24822_ _10392_ net2822 _10621_ VGND VGND VPWR VPWR _10625_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28590_ _12741_ net2897 _12786_ VGND VGND VPWR VPWR _12790_ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27541_ _12136_ net2795 _12197_ VGND VGND VPWR VPWR _12203_ sky130_fd_sc_hd__mux2_1
X_24753_ _10396_ net2320 _10580_ VGND VGND VPWR VPWR _10586_ sky130_fd_sc_hd__mux2_1
X_21965_ _08742_ _09195_ VGND VGND VPWR VPWR _09196_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20916_ _07863_ _08205_ VGND VGND VPWR VPWR _08206_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27472_ _12165_ VGND VGND VPWR VPWR _03596_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24684_ _10396_ net3926 _10543_ VGND VGND VPWR VPWR _10549_ sky130_fd_sc_hd__mux2_1
X_21896_ rvcpu.dp.rf.reg_file_arr\[24\]\[27\] rvcpu.dp.rf.reg_file_arr\[25\]\[27\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[27\] rvcpu.dp.rf.reg_file_arr\[27\]\[27\] rvcpu.dp.plfd.InstrD\[15\]
+ _08526_ VGND VGND VPWR VPWR _09131_ sky130_fd_sc_hd__mux4_1
XFILLER_0_84_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_221_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26423_ net1830 _11542_ _11559_ _11534_ VGND VGND VPWR VPWR _03153_ sky130_fd_sc_hd__o211a_1
X_29211_ _10057_ _13123_ VGND VGND VPWR VPWR _13125_ sky130_fd_sc_hd__and2_1
XFILLER_0_166_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23635_ _09273_ net2906 _10182_ VGND VGND VPWR VPWR _10184_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_194_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20847_ datamem.data_ram\[23\]\[14\] _07021_ _06621_ datamem.data_ram\[20\]\[14\]
+ _08136_ VGND VGND VPWR VPWR _08137_ sky130_fd_sc_hd__o221a_1
XFILLER_0_154_608 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29142_ _13087_ VGND VGND VPWR VPWR _04344_ sky130_fd_sc_hd__clkbuf_1
X_26354_ _11509_ VGND VGND VPWR VPWR _11510_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_193_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20778_ _08058_ _08059_ _08067_ VGND VGND VPWR VPWR _08068_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25305_ _10895_ VGND VGND VPWR VPWR _02699_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29073_ _12754_ net3102 _13049_ VGND VGND VPWR VPWR _13051_ sky130_fd_sc_hd__mux2_1
X_22517_ rvcpu.dp.rf.reg_file_arr\[20\]\[11\] rvcpu.dp.rf.reg_file_arr\[21\]\[11\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[11\] rvcpu.dp.rf.reg_file_arr\[23\]\[11\] _09434_
+ _09558_ VGND VGND VPWR VPWR _09672_ sky130_fd_sc_hd__mux4_1
XFILLER_0_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26285_ net1783 _11467_ VGND VGND VPWR VPWR _11475_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_663 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28024_ _12474_ VGND VGND VPWR VPWR _03839_ sky130_fd_sc_hd__clkbuf_1
X_25236_ _10724_ net3318 net55 VGND VGND VPWR VPWR _10858_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22448_ _09415_ _09603_ _09606_ VGND VGND VPWR VPWR _09607_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_21_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_590 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25167_ _09313_ VGND VGND VPWR VPWR _10818_ sky130_fd_sc_hd__buf_2
X_23866__428 clknet_1_1__leaf__10220_ VGND VGND VPWR VPWR net554 sky130_fd_sc_hd__inv_2
XFILLER_0_0_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22379_ rvcpu.dp.rf.reg_file_arr\[28\]\[4\] rvcpu.dp.rf.reg_file_arr\[30\]\[4\] rvcpu.dp.rf.reg_file_arr\[29\]\[4\]
+ rvcpu.dp.rf.reg_file_arr\[31\]\[4\] _09446_ _09402_ VGND VGND VPWR VPWR _09541_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_27_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24118_ clknet_1_0__leaf__10244_ VGND VGND VPWR VPWR _10260_ sky130_fd_sc_hd__buf_1
XFILLER_0_103_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25098_ _10061_ _10779_ _10781_ net1317 VGND VGND VPWR VPWR _02606_ sky130_fd_sc_hd__a22o_1
X_29975_ net345 _01710_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[14\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28926_ _12751_ net2284 _12968_ VGND VGND VPWR VPWR _12969_ sky130_fd_sc_hd__mux2_1
X_16940_ _04721_ VGND VGND VPWR VPWR _01571_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_198_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23409__1024 clknet_1_1__leaf__10140_ VGND VGND VPWR VPWR net1150 sky130_fd_sc_hd__inv_2
XFILLER_0_217_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16871_ net3037 _14420_ _04684_ VGND VGND VPWR VPWR _04685_ sky130_fd_sc_hd__mux2_1
X_28857_ _12178_ _10997_ _12886_ VGND VGND VPWR VPWR _12932_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_216_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18610_ _05799_ _05855_ VGND VGND VPWR VPWR _05968_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_240_clk clknet_5_17__leaf_clk VGND VGND VPWR VPWR clknet_leaf_240_clk
+ sky130_fd_sc_hd__clkbuf_8
X_27808_ _12142_ net3967 net78 VGND VGND VPWR VPWR _12347_ sky130_fd_sc_hd__mux2_1
X_15822_ _14242_ VGND VGND VPWR VPWR _02110_ sky130_fd_sc_hd__clkbuf_1
X_19590_ _06714_ _06880_ _06885_ VGND VGND VPWR VPWR _06886_ sky130_fd_sc_hd__or3_1
XFILLER_0_204_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28788_ _12895_ VGND VGND VPWR VPWR _04182_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18541_ _05674_ _05901_ VGND VGND VPWR VPWR _05902_ sky130_fd_sc_hd__or2_1
X_15753_ _14205_ VGND VGND VPWR VPWR _02150_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_172_1247 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27739_ _12128_ net3385 _12307_ VGND VGND VPWR VPWR _12309_ sky130_fd_sc_hd__mux2_1
X_14704_ _13262_ VGND VGND VPWR VPWR _13263_ sky130_fd_sc_hd__buf_4
XFILLER_0_158_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18472_ _05669_ _05665_ _05821_ _05834_ _05749_ VGND VGND VPWR VPWR _05835_ sky130_fd_sc_hd__a32o_1
X_30750_ clknet_leaf_191_clk _02485_ VGND VGND VPWR VPWR datamem.data_ram\[48\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15684_ _13225_ VGND VGND VPWR VPWR _14160_ sky130_fd_sc_hd__buf_4
XFILLER_0_206_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_340 _14466_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_351 rvcpu.ALUResultE\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_200_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29409_ clknet_leaf_290_clk _01144_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD2E\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_362 rvcpu.dp.SrcBFW_Mux.y\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14635_ net2331 _13210_ _13181_ VGND VGND VPWR VPWR _13211_ sky130_fd_sc_hd__mux2_1
X_17423_ _14137_ net4032 _04974_ VGND VGND VPWR VPWR _04978_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_215_5644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30681_ clknet_leaf_96_clk _02416_ VGND VGND VPWR VPWR datamem.data_ram\[4\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_373 rvcpu.dp.plem.ALUResultM\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_215_5655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_384 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_395 _01052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_215_5666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32420_ clknet_leaf_80_clk _03842_ VGND VGND VPWR VPWR datamem.data_ram\[28\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17354_ _04941_ VGND VGND VPWR VPWR _01361_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16305_ _14515_ VGND VGND VPWR VPWR _01884_ sky130_fd_sc_hd__clkbuf_1
X_32351_ clknet_leaf_87_clk _03773_ VGND VGND VPWR VPWR datamem.data_ram\[30\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_17285_ rvcpu.dp.rf.reg_file_arr\[24\]\[29\] _13186_ _04902_ VGND VGND VPWR VPWR
+ _04905_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31302_ clknet_leaf_51_clk _03005_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCPlus4E\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_19024_ _06356_ VGND VGND VPWR VPWR rvcpu.dp.lAuiPCE\[0\] sky130_fd_sc_hd__clkbuf_1
X_16236_ _13262_ VGND VGND VPWR VPWR _14476_ sky130_fd_sc_hd__buf_4
XFILLER_0_113_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload304 clknet_1_1__leaf__10201_ VGND VGND VPWR VPWR clkload304/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload12 clknet_5_14__leaf_clk VGND VGND VPWR VPWR clkload12/Y sky130_fd_sc_hd__inv_6
XFILLER_0_183_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload315 clknet_1_0__leaf__10178_ VGND VGND VPWR VPWR clkload315/Y sky130_fd_sc_hd__clkinvlp_4
X_32282_ clknet_leaf_260_clk _03704_ VGND VGND VPWR VPWR datamem.data_ram\[33\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload23 clknet_5_28__leaf_clk VGND VGND VPWR VPWR clkload23/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_125_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload326 clknet_1_1__leaf__11601_ VGND VGND VPWR VPWR clkload326/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_152_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload34 clknet_leaf_14_clk VGND VGND VPWR VPWR clkload34/Y sky130_fd_sc_hd__inv_8
Xclkload337 clknet_1_0__leaf__10131_ VGND VGND VPWR VPWR clkload337/Y sky130_fd_sc_hd__clkinvlp_4
X_31233_ clknet_leaf_32_clk net1669 VGND VGND VPWR VPWR rvcpu.dp.plfd.PCD\[22\] sky130_fd_sc_hd__dfxtp_1
Xclkload45 clknet_leaf_35_clk VGND VGND VPWR VPWR clkload45/Y sky130_fd_sc_hd__clkinv_1
Xclkload348 clknet_1_0__leaf__10107_ VGND VGND VPWR VPWR clkload348/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_2_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16167_ _14429_ VGND VGND VPWR VPWR _01944_ sky130_fd_sc_hd__clkbuf_1
Xclkload56 clknet_leaf_283_clk VGND VGND VPWR VPWR clkload56/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload359 clknet_1_1__leaf__10081_ VGND VGND VPWR VPWR clkload359/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload67 clknet_leaf_65_clk VGND VGND VPWR VPWR clkload67/X sky130_fd_sc_hd__clkbuf_4
Xclkload78 clknet_leaf_40_clk VGND VGND VPWR VPWR clkload78/Y sky130_fd_sc_hd__clkinv_1
XFILLER_0_140_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_71_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15118_ _13417_ _13590_ VGND VGND VPWR VPWR _13663_ sky130_fd_sc_hd__nor2_1
Xclkload89 clknet_leaf_61_clk VGND VGND VPWR VPWR clkload89/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_11_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31164_ clknet_leaf_28_clk rvcpu.ALUResultE\[23\] VGND VGND VPWR VPWR rvcpu.dp.plem.ALUResultM\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_16098_ net2592 _13198_ _14385_ VGND VGND VPWR VPWR _14391_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_166_4474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24064__591 clknet_1_0__leaf__10247_ VGND VGND VPWR VPWR net717 sky130_fd_sc_hd__inv_2
XFILLER_0_227_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_4485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30115_ net477 _01850_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[10\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_15049_ _13580_ _13584_ _13595_ VGND VGND VPWR VPWR _13596_ sky130_fd_sc_hd__a21oi_1
X_19926_ datamem.data_ram\[55\]\[17\] _06784_ _06806_ datamem.data_ram\[52\]\[17\]
+ _07220_ VGND VGND VPWR VPWR _07221_ sky130_fd_sc_hd__o221a_1
XFILLER_0_76_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31095_ clknet_leaf_254_clk _02830_ VGND VGND VPWR VPWR datamem.data_ram\[9\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2807 datamem.data_ram\[8\]\[9\] VGND VGND VPWR VPWR net3957 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_177_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2818 datamem.data_ram\[29\]\[27\] VGND VGND VPWR VPWR net3968 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2829 datamem.data_ram\[5\]\[23\] VGND VGND VPWR VPWR net3979 sky130_fd_sc_hd__dlygate4sd3_1
X_30046_ net408 _01781_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[12\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_19857_ _07071_ _07146_ _07151_ _06985_ VGND VGND VPWR VPWR _07152_ sky130_fd_sc_hd__a31o_1
XFILLER_0_177_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_179_4802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_231_clk clknet_5_20__leaf_clk VGND VGND VPWR VPWR clknet_leaf_231_clk
+ sky130_fd_sc_hd__clkbuf_8
X_18808_ _05698_ _06004_ _05798_ _05703_ VGND VGND VPWR VPWR _06155_ sky130_fd_sc_hd__a31o_1
XFILLER_0_78_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19788_ datamem.data_ram\[43\]\[9\] _07077_ _07078_ _07082_ VGND VGND VPWR VPWR _07083_
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_69_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_69_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18739_ _06081_ _06069_ _06089_ _06085_ VGND VGND VPWR VPWR _06090_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_125_3492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31997_ clknet_leaf_128_clk _03419_ VGND VGND VPWR VPWR datamem.data_ram\[31\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_65_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21750_ _08798_ _08990_ _08992_ _08806_ VGND VGND VPWR VPWR _08993_ sky130_fd_sc_hd__o211a_1
X_30948_ clknet_leaf_86_clk _02683_ VGND VGND VPWR VPWR datamem.data_ram\[3\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_121_3389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20701_ datamem.data_ram\[1\]\[5\] _07133_ _07988_ _07991_ VGND VGND VPWR VPWR _07992_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_19_603 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21681_ _08813_ _08927_ _08689_ VGND VGND VPWR VPWR _08928_ sky130_fd_sc_hd__a21o_1
XFILLER_0_175_243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30879_ clknet_leaf_265_clk _02614_ VGND VGND VPWR VPWR datamem.data_ram\[42\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20632_ datamem.data_ram\[6\]\[29\] _06628_ _07230_ datamem.data_ram\[4\]\[29\] VGND
+ VGND VPWR VPWR _07923_ sky130_fd_sc_hd__o22a_1
X_32618_ clknet_leaf_285_clk _04040_ VGND VGND VPWR VPWR datamem.data_ram\[20\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_3706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_184_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_3717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20563_ datamem.data_ram\[9\]\[21\] _07808_ _07847_ _07853_ VGND VGND VPWR VPWR _07854_
+ sky130_fd_sc_hd__o211a_1
Xclkload6 clknet_5_7__leaf_clk VGND VGND VPWR VPWR clkload6/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_18_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32549_ clknet_leaf_288_clk _03971_ VGND VGND VPWR VPWR datamem.data_ram\[23\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_99_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22302_ _09466_ VGND VGND VPWR VPWR _09467_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_229_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26070_ _06568_ rvcpu.dp.plfd.InstrD\[13\] _06567_ _03029_ VGND VGND VPWR VPWR _11365_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_171_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20494_ _07784_ _07785_ VGND VGND VPWR VPWR _04441_ sky130_fd_sc_hd__nand2_1
XFILLER_0_144_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25021_ _10734_ VGND VGND VPWR VPWR _02576_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22233_ _09398_ VGND VGND VPWR VPWR _09399_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_95_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23253__900 clknet_1_1__leaf__10127_ VGND VGND VPWR VPWR net1026 sky130_fd_sc_hd__inv_2
XFILLER_0_14_396 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22164_ _09353_ VGND VGND VPWR VPWR _01100_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21115_ datamem.data_ram\[26\]\[7\] _06929_ _06935_ datamem.data_ram\[24\]\[7\] _08403_
+ VGND VGND VPWR VPWR _08404_ sky130_fd_sc_hd__a221o_1
X_29760_ net1106 _01495_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[21\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_26972_ _11829_ _11866_ VGND VGND VPWR VPWR _11870_ sky130_fd_sc_hd__and2_1
X_22095_ _09307_ VGND VGND VPWR VPWR _01077_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28711_ _12854_ VGND VGND VPWR VPWR _04146_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_227_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25923_ net1869 _11275_ _11273_ _11281_ VGND VGND VPWR VPWR _02931_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_54_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21046_ _08333_ _08334_ _07819_ VGND VGND VPWR VPWR _08335_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29691_ net1037 _01426_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[23\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_54_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_222_clk clknet_5_21__leaf_clk VGND VGND VPWR VPWR clknet_leaf_222_clk
+ sky130_fd_sc_hd__clkbuf_8
X_25854_ rvcpu.dp.pcreg.q\[26\] _11226_ rvcpu.dp.pcreg.q\[27\] VGND VGND VPWR VPWR
+ _11235_ sky130_fd_sc_hd__a21oi_1
X_28642_ _12741_ net4191 net71 VGND VGND VPWR VPWR _12818_ sky130_fd_sc_hd__mux2_1
XFILLER_0_214_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24805_ _10446_ net3537 _10612_ VGND VGND VPWR VPWR _10616_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25785_ net1736 _11144_ _11177_ _11180_ VGND VGND VPWR VPWR _02894_ sky130_fd_sc_hd__o211a_1
XFILLER_0_202_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28573_ _12758_ net3152 _12777_ VGND VGND VPWR VPWR _12781_ sky130_fd_sc_hd__mux2_1
X_24736_ _10450_ net3927 _10571_ VGND VGND VPWR VPWR _10577_ sky130_fd_sc_hd__mux2_1
X_27524_ _12091_ net3340 net99 VGND VGND VPWR VPWR _12194_ sky130_fd_sc_hd__mux2_1
X_21948_ _09178_ _09179_ _08540_ VGND VGND VPWR VPWR _09180_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27455_ _12155_ net3925 _12143_ VGND VGND VPWR VPWR _12156_ sky130_fd_sc_hd__mux2_1
X_24667_ _10538_ net1567 _10531_ _10539_ VGND VGND VPWR VPWR _02417_ sky130_fd_sc_hd__a31o_1
X_21879_ _08686_ _09114_ _08806_ VGND VGND VPWR VPWR _09115_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_127_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26406_ _13439_ _11542_ _11547_ _11534_ VGND VGND VPWR VPWR _03148_ sky130_fd_sc_hd__o211a_1
XFILLER_0_194_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27386_ _12112_ VGND VGND VPWR VPWR _03563_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24598_ _06591_ VGND VGND VPWR VPWR _10500_ sky130_fd_sc_hd__buf_4
XFILLER_0_108_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26337_ _11089_ _11497_ VGND VGND VPWR VPWR _11504_ sky130_fd_sc_hd__and2_1
XFILLER_0_181_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29125_ _13078_ VGND VGND VPWR VPWR _04336_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_210_5530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_210_5541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17070_ net2632 _14484_ _04756_ VGND VGND VPWR VPWR _04790_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29056_ _09272_ net3829 net65 VGND VGND VPWR VPWR _13042_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26268_ net1854 _11432_ VGND VGND VPWR VPWR _11466_ sky130_fd_sc_hd__and2_1
XFILLER_0_134_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16021_ _14350_ VGND VGND VPWR VPWR _02011_ sky130_fd_sc_hd__clkbuf_1
X_25219_ _10751_ net4168 _10848_ VGND VGND VPWR VPWR _10849_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28007_ _12465_ VGND VGND VPWR VPWR _03831_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26199_ _11437_ VGND VGND VPWR VPWR _03051_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_208_5481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_390 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_208_5492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17972_ rvcpu.dp.plde.ImmExtE\[7\] rvcpu.dp.SrcBFW_Mux.y\[7\] _05278_ VGND VGND VPWR
+ VPWR _05343_ sky130_fd_sc_hd__mux2_1
X_29958_ net328 _01693_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[15\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19711_ datamem.data_ram\[18\]\[0\] _06989_ _07005_ _07006_ VGND VGND VPWR VPWR _07007_
+ sky130_fd_sc_hd__a211o_1
X_16923_ net2707 _14474_ _04706_ VGND VGND VPWR VPWR _04712_ sky130_fd_sc_hd__mux2_1
X_28909_ _12687_ net3040 _12959_ VGND VGND VPWR VPWR _12960_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29889_ net267 _01624_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[17\]\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_204_5389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_4360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_213_clk clknet_5_20__leaf_clk VGND VGND VPWR VPWR clknet_leaf_213_clk
+ sky130_fd_sc_hd__clkbuf_8
X_19642_ datamem.data_ram\[34\]\[0\] _06932_ _06937_ datamem.data_ram\[32\]\[0\] VGND
+ VGND VPWR VPWR _06938_ sky130_fd_sc_hd__a22o_1
X_31920_ _04432_ net119 VGND VGND VPWR VPWR datamem.rd_data_mem\[25\] sky130_fd_sc_hd__dlxtn_1
XTAP_TAPCELL_ROW_161_4371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16854_ _04675_ VGND VGND VPWR VPWR _01611_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_172_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15805_ _14232_ VGND VGND VPWR VPWR _02125_ sky130_fd_sc_hd__clkbuf_1
X_31851_ clknet_leaf_124_clk _03305_ VGND VGND VPWR VPWR datamem.data_ram\[61\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19573_ datamem.data_ram\[4\]\[8\] _06620_ _06868_ _06776_ VGND VGND VPWR VPWR _06869_
+ sky130_fd_sc_hd__o211a_1
X_16785_ net2073 _14472_ _04634_ VGND VGND VPWR VPWR _04639_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_217_5706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18524_ _05585_ _05809_ _05884_ VGND VGND VPWR VPWR _05885_ sky130_fd_sc_hd__and3_1
X_30802_ clknet_leaf_221_clk _02537_ VGND VGND VPWR VPWR datamem.data_ram\[45\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15736_ _13277_ VGND VGND VPWR VPWR _14195_ sky130_fd_sc_hd__buf_4
XFILLER_0_87_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31782_ clknet_leaf_278_clk _03236_ VGND VGND VPWR VPWR datamem.data_ram\[6\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18455_ _05696_ _05702_ _05798_ _05807_ _05817_ VGND VGND VPWR VPWR _05818_ sky130_fd_sc_hd__a311o_1
X_30733_ clknet_leaf_223_clk _02468_ VGND VGND VPWR VPWR datamem.data_ram\[47\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_170 _08693_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15667_ _14148_ VGND VGND VPWR VPWR _02179_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_608 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_181 _09024_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17406_ _04968_ VGND VGND VPWR VPWR _01336_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_192 _09297_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_213_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14618_ _13197_ VGND VGND VPWR VPWR _13198_ sky130_fd_sc_hd__buf_4
XFILLER_0_200_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18386_ _05590_ _05749_ VGND VGND VPWR VPWR _05750_ sky130_fd_sc_hd__nand2_2
X_30664_ clknet_leaf_143_clk _02399_ VGND VGND VPWR VPWR datamem.data_ram\[50\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15598_ net3644 _13223_ _14103_ VGND VGND VPWR VPWR _14107_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32403_ clknet_leaf_247_clk _03825_ VGND VGND VPWR VPWR datamem.data_ram\[29\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_23734__325 clknet_1_0__leaf__10199_ VGND VGND VPWR VPWR net451 sky130_fd_sc_hd__inv_2
XFILLER_0_55_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17337_ net4338 _13265_ _04924_ VGND VGND VPWR VPWR _04932_ sky130_fd_sc_hd__mux2_1
X_30595_ clknet_leaf_117_clk _02330_ VGND VGND VPWR VPWR datamem.data_ram\[53\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_279 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32334_ clknet_leaf_250_clk _03756_ VGND VGND VPWR VPWR datamem.data_ram\[31\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload101 clknet_leaf_87_clk VGND VGND VPWR VPWR clkload101/Y sky130_fd_sc_hd__clkinvlp_2
X_17268_ _14187_ net2520 _04887_ VGND VGND VPWR VPWR _04895_ sky130_fd_sc_hd__mux2_1
Xclkload112 clknet_leaf_99_clk VGND VGND VPWR VPWR clkload112/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_12_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload123 clknet_leaf_250_clk VGND VGND VPWR VPWR clkload123/Y sky130_fd_sc_hd__clkinvlp_2
XTAP_TAPCELL_ROW_168_4525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19007_ _05776_ _05960_ VGND VGND VPWR VPWR _06341_ sky130_fd_sc_hd__nor2_1
Xclkload134 clknet_leaf_288_clk VGND VGND VPWR VPWR clkload134/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_109_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_168_4536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16219_ net2556 _14463_ _14464_ VGND VGND VPWR VPWR _14465_ sky130_fd_sc_hd__mux2_1
Xclkload145 clknet_leaf_263_clk VGND VGND VPWR VPWR clkload145/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_102_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_183_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17199_ _04858_ VGND VGND VPWR VPWR _01441_ sky130_fd_sc_hd__clkbuf_1
X_32265_ clknet_leaf_226_clk _03687_ VGND VGND VPWR VPWR datamem.data_ram\[33\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload156 clknet_leaf_279_clk VGND VGND VPWR VPWR clkload156/Y sky130_fd_sc_hd__clkinv_4
Xclkload167 clknet_leaf_268_clk VGND VGND VPWR VPWR clkload167/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload178 clknet_leaf_233_clk VGND VGND VPWR VPWR clkload178/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_0_87_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31216_ clknet_leaf_37_clk _02919_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCD\[5\] sky130_fd_sc_hd__dfxtp_1
Xclkload189 clknet_leaf_223_clk VGND VGND VPWR VPWR clkload189/Y sky130_fd_sc_hd__inv_8
XFILLER_0_87_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32196_ clknet_leaf_225_clk _03618_ VGND VGND VPWR VPWR datamem.data_ram\[36\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_90_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_1192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_90_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31147_ clknet_leaf_64_clk rvcpu.ALUResultE\[6\] VGND VGND VPWR VPWR rvcpu.dp.plem.ALUResultM\[6\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_227_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2604 datamem.data_ram\[55\]\[11\] VGND VGND VPWR VPWR net3754 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2615 datamem.data_ram\[63\]\[21\] VGND VGND VPWR VPWR net3765 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19909_ datamem.data_ram\[45\]\[17\] _06665_ _06701_ datamem.data_ram\[41\]\[17\]
+ VGND VGND VPWR VPWR _07204_ sky130_fd_sc_hd__o22a_1
Xhold2626 rvcpu.dp.rf.reg_file_arr\[22\]\[18\] VGND VGND VPWR VPWR net3776 sky130_fd_sc_hd__dlygate4sd3_1
X_31078_ clknet_leaf_101_clk _02813_ VGND VGND VPWR VPWR datamem.data_ram\[20\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold18 rvcpu.dp.plem.PCPlus4M\[21\] VGND VGND VPWR VPWR net1168 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_127_3532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold29 rvcpu.dp.plde.ResultSrcE\[1\] VGND VGND VPWR VPWR net1179 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_127_3543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2637 datamem.data_ram\[58\]\[23\] VGND VGND VPWR VPWR net3787 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2648 datamem.data_ram\[27\]\[21\] VGND VGND VPWR VPWR net3798 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_127_3554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1903 rvcpu.dp.rf.reg_file_arr\[1\]\[21\] VGND VGND VPWR VPWR net3053 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1914 datamem.data_ram\[28\]\[21\] VGND VGND VPWR VPWR net3064 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_204_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_204_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold2659 datamem.data_ram\[50\]\[8\] VGND VGND VPWR VPWR net3809 sky130_fd_sc_hd__dlygate4sd3_1
X_22920_ _10048_ _10053_ VGND VGND VPWR VPWR _10054_ sky130_fd_sc_hd__and2_1
Xhold1925 datamem.data_ram\[21\]\[19\] VGND VGND VPWR VPWR net3075 sky130_fd_sc_hd__dlygate4sd3_1
X_30029_ net391 _01764_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[13\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1936 datamem.data_ram\[40\]\[27\] VGND VGND VPWR VPWR net3086 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1947 rvcpu.dp.rf.reg_file_arr\[21\]\[2\] VGND VGND VPWR VPWR net3097 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_3_Left_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1958 rvcpu.dp.rf.reg_file_arr\[12\]\[24\] VGND VGND VPWR VPWR net3108 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1969 datamem.data_ram\[38\]\[27\] VGND VGND VPWR VPWR net3119 sky130_fd_sc_hd__dlygate4sd3_1
X_22851_ _09380_ _09987_ VGND VGND VPWR VPWR _09988_ sky130_fd_sc_hd__or2_1
X_23283__926 clknet_1_1__leaf__10131_ VGND VGND VPWR VPWR net1052 sky130_fd_sc_hd__inv_2
XFILLER_0_97_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21802_ _08522_ _09041_ VGND VGND VPWR VPWR _09042_ sky130_fd_sc_hd__or2_1
XFILLER_0_223_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25570_ _11018_ net1499 _11041_ _11045_ VGND VGND VPWR VPWR _02814_ sky130_fd_sc_hd__a31o_1
XFILLER_0_195_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22782_ _09422_ _09922_ VGND VGND VPWR VPWR _09923_ sky130_fd_sc_hd__nor2_1
XFILLER_0_190_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24521_ _10455_ VGND VGND VPWR VPWR _02355_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21733_ _08510_ _08976_ VGND VGND VPWR VPWR _08977_ sky130_fd_sc_hd__nor2_1
X_24114__621 clknet_1_1__leaf__10259_ VGND VGND VPWR VPWR net747 sky130_fd_sc_hd__inv_2
XFILLER_0_137_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27240_ _12022_ net1443 _12030_ _12033_ VGND VGND VPWR VPWR _03496_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_26_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24452_ _10412_ net4411 _10404_ _10414_ VGND VGND VPWR VPWR _02327_ sky130_fd_sc_hd__a31o_1
XFILLER_0_143_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21664_ rvcpu.dp.rf.reg_file_arr\[8\]\[14\] rvcpu.dp.rf.reg_file_arr\[10\]\[14\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[14\] rvcpu.dp.rf.reg_file_arr\[11\]\[14\] _08693_
+ _08818_ VGND VGND VPWR VPWR _08912_ sky130_fd_sc_hd__mux4_2
X_23408__1023 clknet_1_1__leaf__10140_ VGND VGND VPWR VPWR net1149 sky130_fd_sc_hd__inv_2
XFILLER_0_149_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27171_ _11978_ _11984_ VGND VGND VPWR VPWR _11992_ sky130_fd_sc_hd__and2_1
X_20615_ datamem.data_ram\[31\]\[13\] _06705_ _06618_ datamem.data_ram\[28\]\[13\]
+ _07905_ VGND VGND VPWR VPWR _07906_ sky130_fd_sc_hd__o221a_1
X_24383_ _10370_ VGND VGND VPWR VPWR _02302_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21595_ rvcpu.dp.rf.reg_file_arr\[16\]\[11\] rvcpu.dp.rf.reg_file_arr\[17\]\[11\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[11\] rvcpu.dp.rf.reg_file_arr\[19\]\[11\] _08524_
+ _08527_ VGND VGND VPWR VPWR _08846_ sky130_fd_sc_hd__mux4_1
XFILLER_0_89_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26122_ _11396_ VGND VGND VPWR VPWR _03014_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_49_Left_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20546_ _07836_ VGND VGND VPWR VPWR _07837_ sky130_fd_sc_hd__buf_6
XFILLER_0_127_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26053_ _11353_ net1805 _11350_ _11355_ VGND VGND VPWR VPWR _02987_ sky130_fd_sc_hd__a31o_1
XFILLER_0_43_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20477_ datamem.data_ram\[53\]\[20\] _06662_ _06705_ datamem.data_ram\[55\]\[20\]
+ VGND VGND VPWR VPWR _07769_ sky130_fd_sc_hd__o22a_1
XFILLER_0_63_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25004_ _10454_ net1952 _10715_ VGND VGND VPWR VPWR _10723_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_197_Right_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22216_ _09381_ VGND VGND VPWR VPWR _09382_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_63_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23196_ _09244_ datamem.data_ram\[5\]\[19\] _10115_ VGND VGND VPWR VPWR _10119_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_56_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29812_ net1150 _01547_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[1\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_22147_ _09343_ VGND VGND VPWR VPWR _01093_ sky130_fd_sc_hd__clkbuf_1
X_24160__663 clknet_1_1__leaf__10263_ VGND VGND VPWR VPWR net789 sky130_fd_sc_hd__inv_2
X_29743_ net1089 _01478_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[21\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_26955_ _11849_ net1514 _11853_ _11859_ VGND VGND VPWR VPWR _03385_ sky130_fd_sc_hd__a31o_1
X_22078_ _09292_ VGND VGND VPWR VPWR _01075_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_195_1044 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25906_ net1690 _11256_ _11258_ _11271_ VGND VGND VPWR VPWR _02924_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_58_Left_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21029_ datamem.data_ram\[16\]\[31\] _07912_ VGND VGND VPWR VPWR _08318_ sky130_fd_sc_hd__or2_1
X_29674_ net1020 _01409_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[23\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_26886_ _11813_ net1447 _11809_ _11815_ VGND VGND VPWR VPWR _03360_ sky130_fd_sc_hd__a31o_1
X_28625_ _12758_ net3176 _12805_ VGND VGND VPWR VPWR _12809_ sky130_fd_sc_hd__mux2_1
X_25837_ rvcpu.dp.pcreg.q\[24\] rvcpu.dp.pcreg.q\[23\] _11213_ VGND VGND VPWR VPWR
+ _11221_ sky130_fd_sc_hd__and3_1
XFILLER_0_214_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_202_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16570_ _04524_ VGND VGND VPWR VPWR _01760_ sky130_fd_sc_hd__clkbuf_1
X_28556_ _12694_ net3390 _12768_ VGND VGND VPWR VPWR _12772_ sky130_fd_sc_hd__mux2_1
X_25768_ net1776 _11144_ _11147_ _11167_ VGND VGND VPWR VPWR _02890_ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15521_ _13949_ _14020_ _13304_ VGND VGND VPWR VPWR _14048_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27507_ _12153_ net2245 _12179_ VGND VGND VPWR VPWR _12185_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24719_ _10567_ VGND VGND VPWR VPWR _02441_ sky130_fd_sc_hd__clkbuf_1
X_25699_ _11064_ _11113_ VGND VGND VPWR VPWR _11122_ sky130_fd_sc_hd__and2_1
XFILLER_0_201_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_191_5076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28487_ _11970_ _12724_ VGND VGND VPWR VPWR _12728_ sky130_fd_sc_hd__and2_1
XFILLER_0_210_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_191_5087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15452_ _13506_ _13399_ _13593_ _13504_ VGND VGND VPWR VPWR _13982_ sky130_fd_sc_hd__o31a_1
X_18240_ _05604_ _05424_ _05431_ _05430_ net102 VGND VGND VPWR VPWR _05605_ sky130_fd_sc_hd__o32a_1
XFILLER_0_127_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27438_ _12144_ VGND VGND VPWR VPWR _03583_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15383_ _13911_ _13916_ _13895_ VGND VGND VPWR VPWR _13917_ sky130_fd_sc_hd__and3b_1
X_18171_ _05533_ _05534_ VGND VGND VPWR VPWR _05536_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_67_Left_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27369_ _12091_ net3695 _12097_ VGND VGND VPWR VPWR _12103_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_663 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17122_ _14177_ net4211 _04815_ VGND VGND VPWR VPWR _04818_ sky130_fd_sc_hd__mux2_1
X_29108_ _13069_ VGND VGND VPWR VPWR _04328_ sky130_fd_sc_hd__clkbuf_1
X_30380_ net726 _02115_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[3\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_150_4094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17053_ _04781_ VGND VGND VPWR VPWR _01510_ sky130_fd_sc_hd__clkbuf_1
X_29039_ _10057_ _13031_ VGND VGND VPWR VPWR _13033_ sky130_fd_sc_hd__and2_1
XFILLER_0_208_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16004_ net1942 _13263_ _14333_ VGND VGND VPWR VPWR _14340_ sky130_fd_sc_hd__mux2_1
X_32050_ clknet_leaf_126_clk _03472_ VGND VGND VPWR VPWR datamem.data_ram\[30\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_164_Right_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_206_5429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_4400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31001_ clknet_leaf_101_clk _02736_ VGND VGND VPWR VPWR datamem.data_ram\[22\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_163_4411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24189__29 clknet_1_1__leaf__10266_ VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__inv_2
XFILLER_0_21_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17955_ rvcpu.dp.plde.RD1E\[12\] _05265_ _05269_ _13240_ _05326_ VGND VGND VPWR VPWR
+ _05327_ sky130_fd_sc_hd__a221o_2
XFILLER_0_225_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16906_ net1989 _14457_ _04695_ VGND VGND VPWR VPWR _04703_ sky130_fd_sc_hd__mux2_1
X_32952_ clknet_leaf_193_clk _04374_ VGND VGND VPWR VPWR datamem.data_ram\[6\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_17886_ rvcpu.dp.plmw.RdW\[2\] rvcpu.dp.plde.Rs1E\[2\] VGND VGND VPWR VPWR _05259_
+ sky130_fd_sc_hd__or2b_1
X_19625_ _06920_ VGND VGND VPWR VPWR _06921_ sky130_fd_sc_hd__buf_4
X_31903_ _04445_ net118 VGND VGND VPWR VPWR datamem.rd_data_mem\[8\] sky130_fd_sc_hd__dlxtn_1
X_16837_ _04666_ VGND VGND VPWR VPWR _01619_ sky130_fd_sc_hd__clkbuf_1
X_32883_ clknet_leaf_250_clk _04305_ VGND VGND VPWR VPWR datamem.data_ram\[10\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_475 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19556_ datamem.data_ram\[12\]\[24\] _06805_ _06850_ _06851_ VGND VGND VPWR VPWR
+ _06852_ sky130_fd_sc_hd__o211a_1
X_31834_ clknet_leaf_215_clk _03288_ VGND VGND VPWR VPWR datamem.data_ram\[3\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_16768_ net2419 _14455_ _04623_ VGND VGND VPWR VPWR _04630_ sky130_fd_sc_hd__mux2_1
XFILLER_0_220_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18507_ _05383_ _05726_ _05808_ _05399_ _05868_ VGND VGND VPWR VPWR _05869_ sky130_fd_sc_hd__a221o_1
XFILLER_0_38_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_4259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15719_ _14183_ net2805 _14173_ VGND VGND VPWR VPWR _14184_ sky130_fd_sc_hd__mux2_1
X_31765_ clknet_leaf_106_clk _03219_ VGND VGND VPWR VPWR datamem.data_ram\[18\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_19487_ _06782_ VGND VGND VPWR VPWR _06783_ sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_83_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16699_ _04593_ VGND VGND VPWR VPWR _01692_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_83_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30716_ clknet_leaf_136_clk _02451_ VGND VGND VPWR VPWR datamem.data_ram\[49\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_18438_ _05581_ _05709_ VGND VGND VPWR VPWR _05801_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31696_ clknet_leaf_50_clk _03154_ VGND VGND VPWR VPWR rvcpu.dp.pcreg.q\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18369_ _05275_ _05733_ VGND VGND VPWR VPWR _05734_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30647_ clknet_leaf_185_clk _02382_ VGND VGND VPWR VPWR datamem.data_ram\[51\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20400_ _05391_ _06586_ _07691_ VGND VGND VPWR VPWR _07692_ sky130_fd_sc_hd__or3_1
XFILLER_0_43_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21380_ _08515_ _08640_ _08513_ VGND VGND VPWR VPWR _08641_ sky130_fd_sc_hd__o21ai_1
X_30578_ clknet_leaf_189_clk _02313_ VGND VGND VPWR VPWR datamem.data_ram\[54\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_116_3277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_3288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20331_ datamem.data_ram\[46\]\[4\] _07159_ _06949_ datamem.data_ram\[41\]\[4\] _07622_
+ VGND VGND VPWR VPWR _07623_ sky130_fd_sc_hd__a221o_1
X_32317_ clknet_leaf_229_clk _03739_ VGND VGND VPWR VPWR datamem.data_ram\[31\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_189_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_187_4978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput19 net19 VGND VGND VPWR VPWR Instr[25] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_187_4989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20262_ datamem.data_ram\[53\]\[19\] _06703_ _06707_ datamem.data_ram\[55\]\[19\]
+ VGND VGND VPWR VPWR _07555_ sky130_fd_sc_hd__o22a_1
X_32248_ clknet_leaf_208_clk _03670_ VGND VGND VPWR VPWR datamem.data_ram\[34\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_131_Right_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22001_ _09230_ VGND VGND VPWR VPWR _09231_ sky130_fd_sc_hd__buf_8
Xhold3102 rvcpu.dp.rf.reg_file_arr\[19\]\[6\] VGND VGND VPWR VPWR net4252 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3113 datamem.data_ram\[54\]\[23\] VGND VGND VPWR VPWR net4263 sky130_fd_sc_hd__dlygate4sd3_1
X_20193_ datamem.data_ram\[47\]\[11\] _06761_ _07485_ _06742_ VGND VGND VPWR VPWR
+ _07486_ sky130_fd_sc_hd__o211a_1
X_32179_ clknet_leaf_168_clk _03601_ VGND VGND VPWR VPWR datamem.data_ram\[37\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3124 rvcpu.dp.rf.reg_file_arr\[25\]\[20\] VGND VGND VPWR VPWR net4274 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3135 datamem.data_ram\[54\]\[30\] VGND VGND VPWR VPWR net4285 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2401 datamem.data_ram\[24\]\[13\] VGND VGND VPWR VPWR net3551 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3146 rvcpu.dp.rf.reg_file_arr\[13\]\[31\] VGND VGND VPWR VPWR net4296 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3157 datamem.data_ram\[2\]\[18\] VGND VGND VPWR VPWR net4307 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2412 datamem.data_ram\[20\]\[9\] VGND VGND VPWR VPWR net3562 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2423 datamem.data_ram\[33\]\[21\] VGND VGND VPWR VPWR net3573 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3168 datamem.data_ram\[5\]\[16\] VGND VGND VPWR VPWR net4318 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3179 rvcpu.dp.rf.reg_file_arr\[24\]\[24\] VGND VGND VPWR VPWR net4329 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2434 datamem.data_ram\[21\]\[31\] VGND VGND VPWR VPWR net3584 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2445 datamem.data_ram\[0\]\[16\] VGND VGND VPWR VPWR net3595 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1700 datamem.data_ram\[1\]\[16\] VGND VGND VPWR VPWR net2850 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1711 datamem.data_ram\[37\]\[12\] VGND VGND VPWR VPWR net2861 sky130_fd_sc_hd__dlygate4sd3_1
X_26740_ _11679_ _11726_ VGND VGND VPWR VPWR _11728_ sky130_fd_sc_hd__and2_1
X_23952_ _09224_ net4421 _10229_ VGND VGND VPWR VPWR _10230_ sky130_fd_sc_hd__mux2_1
Xhold2456 datamem.data_ram\[60\]\[12\] VGND VGND VPWR VPWR net3606 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_3996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2467 datamem.data_ram\[17\]\[10\] VGND VGND VPWR VPWR net3617 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1722 datamem.data_ram\[31\]\[31\] VGND VGND VPWR VPWR net2872 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2478 datamem.data_ram\[48\]\[22\] VGND VGND VPWR VPWR net3628 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1733 rvcpu.dp.rf.reg_file_arr\[3\]\[1\] VGND VGND VPWR VPWR net2883 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2489 datamem.data_ram\[47\]\[17\] VGND VGND VPWR VPWR net3639 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1744 rvcpu.dp.rf.reg_file_arr\[4\]\[27\] VGND VGND VPWR VPWR net2894 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1755 datamem.data_ram\[19\]\[12\] VGND VGND VPWR VPWR net2905 sky130_fd_sc_hd__dlygate4sd3_1
X_22903_ _09481_ _10037_ VGND VGND VPWR VPWR _10038_ sky130_fd_sc_hd__and2_1
X_26671_ _10069_ VGND VGND VPWR VPWR _11687_ sky130_fd_sc_hd__buf_2
Xhold1766 datamem.data_ram\[60\]\[24\] VGND VGND VPWR VPWR net2916 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f__10240_ clknet_0__10240_ VGND VGND VPWR VPWR clknet_1_1__leaf__10240_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_169_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_224_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1777 datamem.data_ram\[33\]\[29\] VGND VGND VPWR VPWR net2927 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_223_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1788 datamem.data_ram\[38\]\[28\] VGND VGND VPWR VPWR net2938 sky130_fd_sc_hd__dlygate4sd3_1
X_28410_ _12454_ net2772 _12678_ VGND VGND VPWR VPWR _12682_ sky130_fd_sc_hd__mux2_1
Xhold1799 rvcpu.dp.rf.reg_file_arr\[19\]\[0\] VGND VGND VPWR VPWR net2949 sky130_fd_sc_hd__dlygate4sd3_1
X_25622_ _10946_ _11075_ VGND VGND VPWR VPWR _11076_ sky130_fd_sc_hd__or2_1
X_22834_ _09970_ _09971_ _09449_ VGND VGND VPWR VPWR _09972_ sky130_fd_sc_hd__mux2_1
XFILLER_0_212_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29390_ clknet_leaf_0_clk _01125_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD2E\[1\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__10171_ clknet_0__10171_ VGND VGND VPWR VPWR clknet_1_1__leaf__10171_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_195_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23602__222 clknet_1_1__leaf__10178_ VGND VGND VPWR VPWR net348 sky130_fd_sc_hd__inv_2
XFILLER_0_155_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28341_ _12437_ net3212 _12641_ VGND VGND VPWR VPWR _12645_ sky130_fd_sc_hd__mux2_1
X_25553_ _10760_ net2716 _11030_ VGND VGND VPWR VPWR _11035_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22765_ rvcpu.dp.rf.reg_file_arr\[20\]\[24\] rvcpu.dp.rf.reg_file_arr\[21\]\[24\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[24\] rvcpu.dp.rf.reg_file_arr\[23\]\[24\] _09512_
+ _09408_ VGND VGND VPWR VPWR _09907_ sky130_fd_sc_hd__mux4_1
XFILLER_0_78_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24504_ _09239_ VGND VGND VPWR VPWR _10444_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_17_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28272_ _12607_ VGND VGND VPWR VPWR _03954_ sky130_fd_sc_hd__clkbuf_1
X_21716_ rvcpu.dp.rf.reg_file_arr\[4\]\[17\] rvcpu.dp.rf.reg_file_arr\[5\]\[17\] rvcpu.dp.rf.reg_file_arr\[6\]\[17\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[17\] _08578_ _08684_ VGND VGND VPWR VPWR _08961_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_94_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25484_ _10070_ net35 _10996_ net1314 VGND VGND VPWR VPWR _02777_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22696_ rvcpu.dp.rf.reg_file_arr\[4\]\[20\] rvcpu.dp.rf.reg_file_arr\[5\]\[20\] rvcpu.dp.rf.reg_file_arr\[6\]\[20\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[20\] _09604_ _09716_ VGND VGND VPWR VPWR _09842_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_19_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27223_ _12022_ net1530 _12018_ _12023_ VGND VGND VPWR VPWR _03489_ sky130_fd_sc_hd__a31o_1
X_24435_ _10401_ VGND VGND VPWR VPWR _02323_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_712 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21647_ rvcpu.dp.rf.reg_file_arr\[12\]\[13\] rvcpu.dp.rf.reg_file_arr\[13\]\[13\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[13\] rvcpu.dp.rf.reg_file_arr\[15\]\[13\] _08696_
+ _08568_ VGND VGND VPWR VPWR _08896_ sky130_fd_sc_hd__mux4_1
XFILLER_0_136_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_227_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27154_ _11974_ net1576 _11964_ _11981_ VGND VGND VPWR VPWR _03462_ sky130_fd_sc_hd__a31o_1
XFILLER_0_227_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24366_ _09314_ net2660 net61 VGND VGND VPWR VPWR _10361_ sky130_fd_sc_hd__mux2_1
XANTENNA_70 _06769_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21578_ rvcpu.dp.rf.reg_file_arr\[24\]\[10\] rvcpu.dp.rf.reg_file_arr\[25\]\[10\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[10\] rvcpu.dp.rf.reg_file_arr\[27\]\[10\] _08536_
+ _08519_ VGND VGND VPWR VPWR _08830_ sky130_fd_sc_hd__mux4_1
XANTENNA_81 _06780_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26105_ net1890 _11386_ VGND VGND VPWR VPWR _11388_ sky130_fd_sc_hd__and2_1
XFILLER_0_34_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_92 _06806_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27085_ _11526_ _11936_ VGND VGND VPWR VPWR _11937_ sky130_fd_sc_hd__or2_1
X_20529_ _07819_ VGND VGND VPWR VPWR _07820_ sky130_fd_sc_hd__buf_8
X_24297_ _09285_ net3457 _10316_ VGND VGND VPWR VPWR _10322_ sky130_fd_sc_hd__mux2_1
X_26036_ _11047_ _11340_ VGND VGND VPWR VPWR _11345_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_203_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_0_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_0_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_203_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27987_ _09275_ VGND VGND VPWR VPWR _12452_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_201_5315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_201_5326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29726_ net1072 _01461_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[22\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_17740_ _05145_ VGND VGND VPWR VPWR _01171_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_206_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_197_5230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26938_ _11752_ VGND VGND VPWR VPWR _11849_ sky130_fd_sc_hd__clkbuf_4
X_14952_ _13357_ VGND VGND VPWR VPWR _13501_ sky130_fd_sc_hd__clkbuf_4
X_23231__880 clknet_1_1__leaf__10125_ VGND VGND VPWR VPWR net1006 sky130_fd_sc_hd__inv_2
XFILLER_0_27_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2990 datamem.data_ram\[22\]\[8\] VGND VGND VPWR VPWR net4140 sky130_fd_sc_hd__dlygate4sd3_1
X_17671_ net4331 _13256_ _05104_ VGND VGND VPWR VPWR _05109_ sky130_fd_sc_hd__mux2_1
X_29657_ net1003 _01392_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[24\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_26869_ _11687_ _11798_ VGND VGND VPWR VPWR _11805_ sky130_fd_sc_hd__and2_1
X_14883_ _13289_ _13434_ VGND VGND VPWR VPWR _13435_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_193_5116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_193_5127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_193_5138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19410_ _06705_ VGND VGND VPWR VPWR _06706_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_203_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16622_ _14154_ net3110 _04551_ VGND VGND VPWR VPWR _04553_ sky130_fd_sc_hd__mux2_1
X_28608_ _12694_ net3748 _12796_ VGND VGND VPWR VPWR _12800_ sky130_fd_sc_hd__mux2_1
XFILLER_0_202_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29588_ net942 _01323_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[26\]\[23\] sky130_fd_sc_hd__dfxtp_1
Xmax_cap50 _12289_ VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__buf_4
XFILLER_0_202_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_212_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap61 _10357_ VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__buf_4
XFILLER_0_186_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19341_ datamem.data_ram\[14\]\[16\] _06630_ _06636_ datamem.data_ram\[11\]\[16\]
+ VGND VGND VPWR VPWR _06637_ sky130_fd_sc_hd__o22a_1
Xmax_cap72 _12623_ VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__buf_4
X_28539_ _12761_ VGND VGND VPWR VPWR _04067_ sky130_fd_sc_hd__clkbuf_1
X_16553_ _14154_ net2645 _04514_ VGND VGND VPWR VPWR _04516_ sky130_fd_sc_hd__mux2_1
Xmax_cap83 _12159_ VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__buf_4
X_15504_ _13499_ _14028_ _14031_ _13638_ VGND VGND VPWR VPWR _14032_ sky130_fd_sc_hd__o22a_1
XFILLER_0_155_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_75_Left_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31550_ clknet_leaf_72_clk datamem.rd_data_mem\[0\] VGND VGND VPWR VPWR rvcpu.dp.plmw.ReadDataW\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_19272_ rvcpu.dp.plfd.InstrD\[4\] _06566_ VGND VGND VPWR VPWR _06572_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_14_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16484_ _04479_ VGND VGND VPWR VPWR _01801_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_14_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18223_ _05587_ _05359_ VGND VGND VPWR VPWR _05588_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_155_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_4134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30501_ clknet_leaf_268_clk _02236_ VGND VGND VPWR VPWR datamem.data_ram\[57\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_15435_ _13517_ _13965_ _13953_ _13448_ _13442_ VGND VGND VPWR VPWR _13966_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_152_4145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31481_ clknet_leaf_65_clk rvcpu.dp.lAuiPCE\[7\] VGND VGND VPWR VPWR rvcpu.dp.plem.lAuiPCM\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15366_ _13549_ _13900_ _13409_ VGND VGND VPWR VPWR _13901_ sky130_fd_sc_hd__o21ai_1
X_18154_ _05518_ VGND VGND VPWR VPWR _05519_ sky130_fd_sc_hd__inv_2
X_30432_ net770 _02167_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[29\]\[11\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f__10260_ clknet_0__10260_ VGND VGND VPWR VPWR clknet_1_0__leaf__10260_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_81_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17105_ _14160_ net4277 _04804_ VGND VGND VPWR VPWR _04809_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15297_ _13496_ _13831_ _13832_ _13834_ VGND VGND VPWR VPWR _13835_ sky130_fd_sc_hd__a31o_1
X_18085_ _05406_ _05433_ _05440_ _05452_ VGND VGND VPWR VPWR _05453_ sky130_fd_sc_hd__a31o_1
X_30363_ net709 _02098_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[3\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold307 datamem.data_ram\[18\]\[3\] VGND VGND VPWR VPWR net1457 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__10191_ clknet_0__10191_ VGND VGND VPWR VPWR clknet_1_0__leaf__10191_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_41_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold318 datamem.data_ram\[21\]\[0\] VGND VGND VPWR VPWR net1468 sky130_fd_sc_hd__dlygate4sd3_1
X_32102_ clknet_leaf_114_clk _03524_ VGND VGND VPWR VPWR datamem.data_ram\[23\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold329 datamem.data_ram\[21\]\[7\] VGND VGND VPWR VPWR net1479 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17036_ _04772_ VGND VGND VPWR VPWR _01518_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_229_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_229_5985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23382__1016 clknet_1_0__leaf__10140_ VGND VGND VPWR VPWR net1142 sky130_fd_sc_hd__inv_2
X_30294_ net640 _02029_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[5\]\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_229_5996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32033_ clknet_leaf_131_clk _03455_ VGND VGND VPWR VPWR datamem.data_ram\[50\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_84_Left_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_182_4853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_4864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_182_4875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18987_ _05302_ _06320_ _05561_ VGND VGND VPWR VPWR _06322_ sky130_fd_sc_hd__o21ai_1
X_23407__1022 clknet_1_1__leaf__10140_ VGND VGND VPWR VPWR net1148 sky130_fd_sc_hd__inv_2
Xhold1007 rvcpu.dp.rf.reg_file_arr\[2\]\[13\] VGND VGND VPWR VPWR net2157 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_175_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17938_ rvcpu.dp.plde.ImmExtE\[14\] rvcpu.dp.SrcBFW_Mux.y\[14\] _05277_ VGND VGND
+ VPWR VPWR _05310_ sky130_fd_sc_hd__mux2_2
Xhold1018 rvcpu.dp.rf.reg_file_arr\[2\]\[1\] VGND VGND VPWR VPWR net2168 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1029 rvcpu.dp.rf.reg_file_arr\[17\]\[7\] VGND VGND VPWR VPWR net2179 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32935_ clknet_leaf_139_clk _04357_ VGND VGND VPWR VPWR datamem.data_ram\[7\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_17869_ rvcpu.dp.plde.Rs1E\[1\] rvcpu.dp.plde.Rs1E\[0\] rvcpu.dp.plde.Rs1E\[2\] rvcpu.dp.plde.Rs1E\[4\]
+ VGND VGND VPWR VPWR _05242_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_1_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19608_ datamem.data_ram\[30\]\[8\] _06717_ _06685_ datamem.data_ram\[28\]\[8\] VGND
+ VGND VPWR VPWR _06904_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_141_3871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_3882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20880_ datamem.data_ram\[46\]\[14\] datamem.data_ram\[47\]\[14\] _07827_ VGND VGND
+ VPWR VPWR _08170_ sky130_fd_sc_hd__mux2_1
X_32866_ clknet_leaf_273_clk _04288_ VGND VGND VPWR VPWR datamem.data_ram\[11\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_93_Left_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31817_ clknet_leaf_104_clk _03271_ VGND VGND VPWR VPWR datamem.data_ram\[9\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_19539_ _06827_ _06714_ _06834_ VGND VGND VPWR VPWR _06835_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_81_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_193_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32797_ clknet_leaf_236_clk _04219_ VGND VGND VPWR VPWR datamem.data_ram\[13\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22550_ _09389_ _09695_ _09699_ _09703_ VGND VGND VPWR VPWR _09704_ sky130_fd_sc_hd__and4_1
XFILLER_0_192_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31748_ _04449_ net125 VGND VGND VPWR VPWR rvcpu.ALUControl\[2\] sky130_fd_sc_hd__dlxtn_1
XFILLER_0_146_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_3317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_200_Right_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21501_ rvcpu.dp.rf.reg_file_arr\[0\]\[6\] rvcpu.dp.rf.reg_file_arr\[1\]\[6\] rvcpu.dp.rf.reg_file_arr\[2\]\[6\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[6\] _08566_ _08569_ VGND VGND VPWR VPWR _08757_ sky130_fd_sc_hd__mux4_1
XFILLER_0_173_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22481_ rvcpu.dp.rf.reg_file_arr\[24\]\[9\] rvcpu.dp.rf.reg_file_arr\[25\]\[9\] rvcpu.dp.rf.reg_file_arr\[26\]\[9\]
+ rvcpu.dp.rf.reg_file_arr\[27\]\[9\] _09463_ _09637_ VGND VGND VPWR VPWR _09638_
+ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_44_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31679_ clknet_leaf_9_clk net1274 VGND VGND VPWR VPWR rvcpu.dp.plmw.ALUResultW\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24220_ _09236_ net4369 _10279_ VGND VGND VPWR VPWR _10281_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21432_ _08682_ _08685_ _08690_ VGND VGND VPWR VPWR _08691_ sky130_fd_sc_hd__a21o_1
XFILLER_0_72_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24151_ clknet_1_0__leaf__10244_ VGND VGND VPWR VPWR _10263_ sky130_fd_sc_hd__buf_1
XFILLER_0_31_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21363_ _08624_ VGND VGND VPWR VPWR _08625_ sky130_fd_sc_hd__buf_2
XFILLER_0_114_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20314_ datamem.data_ram\[11\]\[4\] _06943_ _06993_ datamem.data_ram\[15\]\[4\] VGND
+ VGND VPWR VPWR _07606_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24082_ _09279_ net3309 _10249_ VGND VGND VPWR VPWR _10253_ sky130_fd_sc_hd__mux2_1
X_21294_ rvcpu.dp.rf.reg_file_arr\[12\]\[0\] rvcpu.dp.rf.reg_file_arr\[13\]\[0\] rvcpu.dp.rf.reg_file_arr\[14\]\[0\]
+ rvcpu.dp.rf.reg_file_arr\[15\]\[0\] _08551_ _08555_ VGND VGND VPWR VPWR _08556_
+ sky130_fd_sc_hd__mux4_1
Xhold830 rvcpu.dp.rf.reg_file_arr\[11\]\[3\] VGND VGND VPWR VPWR net1980 sky130_fd_sc_hd__dlygate4sd3_1
X_23174__845 clknet_1_0__leaf__10111_ VGND VGND VPWR VPWR net971 sky130_fd_sc_hd__inv_2
Xhold841 rvcpu.dp.rf.reg_file_arr\[9\]\[3\] VGND VGND VPWR VPWR net1991 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold852 datamem.data_ram\[30\]\[14\] VGND VGND VPWR VPWR net2002 sky130_fd_sc_hd__dlygate4sd3_1
X_27910_ _12406_ VGND VGND VPWR VPWR _03793_ sky130_fd_sc_hd__clkbuf_1
X_23033_ clknet_1_0__leaf__10087_ VGND VGND VPWR VPWR _10089_ sky130_fd_sc_hd__buf_1
XFILLER_0_229_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20245_ datamem.data_ram\[61\]\[3\] _06921_ _06680_ _07536_ _07537_ VGND VGND VPWR
+ VPWR _07538_ sky130_fd_sc_hd__a2111o_1
Xhold863 datamem.data_ram\[48\]\[13\] VGND VGND VPWR VPWR net2013 sky130_fd_sc_hd__dlygate4sd3_1
X_28890_ _12949_ VGND VGND VPWR VPWR _04230_ sky130_fd_sc_hd__clkbuf_1
Xhold874 rvcpu.dp.rf.reg_file_arr\[3\]\[30\] VGND VGND VPWR VPWR net2024 sky130_fd_sc_hd__dlygate4sd3_1
Xhold885 datamem.data_ram\[18\]\[22\] VGND VGND VPWR VPWR net2035 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_219_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold896 datamem.data_ram\[12\]\[15\] VGND VGND VPWR VPWR net2046 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_200_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_38_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27841_ _09321_ VGND VGND VPWR VPWR _12367_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_200_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20176_ datamem.data_ram\[22\]\[11\] _06719_ _06754_ datamem.data_ram\[18\]\[11\]
+ _07468_ VGND VGND VPWR VPWR _07469_ sky130_fd_sc_hd__o221a_1
X_23289__932 clknet_1_0__leaf__10131_ VGND VGND VPWR VPWR net1058 sky130_fd_sc_hd__inv_2
Xhold2220 datamem.data_ram\[13\]\[28\] VGND VGND VPWR VPWR net3370 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2231 rvcpu.dp.rf.reg_file_arr\[31\]\[14\] VGND VGND VPWR VPWR net3381 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2242 datamem.data_ram\[10\]\[13\] VGND VGND VPWR VPWR net3392 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27772_ _12080_ net3970 _12326_ VGND VGND VPWR VPWR _12327_ sky130_fd_sc_hd__mux2_1
Xhold2253 datamem.data_ram\[7\]\[12\] VGND VGND VPWR VPWR net3403 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2264 datamem.data_ram\[42\]\[23\] VGND VGND VPWR VPWR net3414 sky130_fd_sc_hd__dlygate4sd3_1
X_24984_ _10712_ VGND VGND VPWR VPWR _02561_ sky130_fd_sc_hd__clkbuf_1
Xhold1530 datamem.data_ram\[0\]\[30\] VGND VGND VPWR VPWR net2680 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2275 datamem.data_ram\[10\]\[8\] VGND VGND VPWR VPWR net3425 sky130_fd_sc_hd__dlygate4sd3_1
X_29511_ net873 _01246_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[28\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_26723_ _11717_ VGND VGND VPWR VPWR _03295_ sky130_fd_sc_hd__clkbuf_1
Xhold1541 datamem.data_ram\[51\]\[30\] VGND VGND VPWR VPWR net2691 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2286 datamem.data_ram\[8\]\[10\] VGND VGND VPWR VPWR net3436 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1552 datamem.data_ram\[6\]\[18\] VGND VGND VPWR VPWR net2702 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2297 datamem.data_ram\[2\]\[9\] VGND VGND VPWR VPWR net3447 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1563 datamem.data_ram\[16\]\[26\] VGND VGND VPWR VPWR net2713 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1574 datamem.data_ram\[24\]\[23\] VGND VGND VPWR VPWR net2724 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1585 rvcpu.dp.rf.reg_file_arr\[4\]\[25\] VGND VGND VPWR VPWR net2735 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29442_ net804 _01177_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[30\]\[13\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__10223_ clknet_0__10223_ VGND VGND VPWR VPWR clknet_1_1__leaf__10223_
+ sky130_fd_sc_hd__clkbuf_16
X_26654_ _11674_ VGND VGND VPWR VPWR _11675_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_170_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1596 datamem.data_ram\[48\]\[31\] VGND VGND VPWR VPWR net2746 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_1128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169_647 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25605_ _10724_ net3623 net53 VGND VGND VPWR VPWR _11067_ sky130_fd_sc_hd__mux2_1
X_22817_ _09451_ _09955_ _09404_ VGND VGND VPWR VPWR _09956_ sky130_fd_sc_hd__o21a_1
X_29373_ clknet_leaf_144_clk _01108_ VGND VGND VPWR VPWR datamem.data_ram\[60\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__10154_ clknet_0__10154_ VGND VGND VPWR VPWR clknet_1_1__leaf__10154_
+ sky130_fd_sc_hd__clkbuf_16
X_26585_ _07191_ _10932_ _11494_ VGND VGND VPWR VPWR _11638_ sky130_fd_sc_hd__or3_1
XFILLER_0_212_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28324_ _12363_ net2922 _12632_ VGND VGND VPWR VPWR _12636_ sky130_fd_sc_hd__mux2_1
X_25536_ _10733_ net4091 net54 VGND VGND VPWR VPWR _11026_ sky130_fd_sc_hd__mux2_1
X_22748_ _09516_ _09888_ _09890_ _09523_ VGND VGND VPWR VPWR _09891_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__10085_ clknet_0__10085_ VGND VGND VPWR VPWR clknet_1_1__leaf__10085_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_149_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26483__37 clknet_1_0__leaf__10267_ VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__inv_2
X_25467_ _10954_ net1545 _10984_ _10989_ VGND VGND VPWR VPWR _02767_ sky130_fd_sc_hd__a31o_1
X_28255_ _12597_ VGND VGND VPWR VPWR _03947_ sky130_fd_sc_hd__clkbuf_1
X_22679_ _09622_ _09823_ _09825_ VGND VGND VPWR VPWR _09826_ sky130_fd_sc_hd__a21o_1
XFILLER_0_165_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15220_ _13385_ _13759_ _13760_ VGND VGND VPWR VPWR _13761_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27206_ _11946_ _12008_ VGND VGND VPWR VPWR _12013_ sky130_fd_sc_hd__and2_1
X_24418_ _09275_ VGND VGND VPWR VPWR _10390_ sky130_fd_sc_hd__buf_2
X_23492__138 clknet_1_0__leaf__10160_ VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__inv_2
X_25398_ _10938_ net1605 _10949_ _10953_ VGND VGND VPWR VPWR _02734_ sky130_fd_sc_hd__a31o_1
X_28186_ _12560_ VGND VGND VPWR VPWR _03915_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15151_ _13692_ _13403_ _13693_ _13694_ VGND VGND VPWR VPWR _13695_ sky130_fd_sc_hd__a31o_1
X_27137_ _10060_ VGND VGND VPWR VPWR _11970_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_180_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24349_ _09279_ net3754 _10348_ VGND VGND VPWR VPWR _10352_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15082_ _13320_ _13346_ VGND VGND VPWR VPWR _13628_ sky130_fd_sc_hd__nor2_2
X_27068_ _11827_ _11924_ VGND VGND VPWR VPWR _11927_ sky130_fd_sc_hd__and2_1
XFILLER_0_132_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26019_ net23 _11152_ VGND VGND VPWR VPWR _11335_ sky130_fd_sc_hd__or2_1
X_18910_ _05525_ _05537_ VGND VGND VPWR VPWR _06250_ sky130_fd_sc_hd__nand2_1
X_19890_ datamem.data_ram\[18\]\[17\] _06612_ _06664_ datamem.data_ram\[21\]\[17\]
+ VGND VGND VPWR VPWR _07185_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_224_5860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18841_ _05698_ _06004_ _05878_ _05703_ VGND VGND VPWR VPWR _06186_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_224_5871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_224_5882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23609__228 clknet_1_1__leaf__10179_ VGND VGND VPWR VPWR net354 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_8_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18772_ _05612_ _06104_ _05318_ VGND VGND VPWR VPWR _06121_ sky130_fd_sc_hd__a21oi_1
X_15984_ _14329_ VGND VGND VPWR VPWR _02035_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_220_5768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_220_5779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29709_ net1055 _01444_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[22\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_17723_ _05136_ VGND VGND VPWR VPWR _01179_ sky130_fd_sc_hd__clkbuf_1
X_14935_ _13284_ _13287_ VGND VGND VPWR VPWR _13484_ sky130_fd_sc_hd__nand2_4
XFILLER_0_145_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30981_ clknet_leaf_116_clk _02716_ VGND VGND VPWR VPWR datamem.data_ram\[39\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_188_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32720_ clknet_leaf_284_clk _04142_ VGND VGND VPWR VPWR datamem.data_ram\[17\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_17654_ net3755 _13231_ _05093_ VGND VGND VPWR VPWR _05100_ sky130_fd_sc_hd__mux2_1
X_14866_ _13417_ _13351_ VGND VGND VPWR VPWR _13418_ sky130_fd_sc_hd__or2b_1
XFILLER_0_159_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16605_ _14137_ net2619 _04540_ VGND VGND VPWR VPWR _04544_ sky130_fd_sc_hd__mux2_1
XFILLER_0_202_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32651_ clknet_leaf_239_clk _04073_ VGND VGND VPWR VPWR datamem.data_ram\[19\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_17585_ _05063_ VGND VGND VPWR VPWR _01244_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_225_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14797_ _13284_ _13305_ VGND VGND VPWR VPWR _13350_ sky130_fd_sc_hd__nand2_4
XFILLER_0_216_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31602_ clknet_leaf_45_clk net1205 VGND VGND VPWR VPWR rvcpu.dp.plmw.PCPlus4W\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19324_ _06619_ VGND VGND VPWR VPWR _06620_ sky130_fd_sc_hd__buf_8
X_16536_ _14137_ net3487 _04503_ VGND VGND VPWR VPWR _04507_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32582_ clknet_leaf_247_clk _04004_ VGND VGND VPWR VPWR datamem.data_ram\[21\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_175_4690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19255_ _06555_ _06557_ VGND VGND VPWR VPWR _06558_ sky130_fd_sc_hd__xnor2_1
X_31533_ clknet_leaf_25_clk net1219 VGND VGND VPWR VPWR rvcpu.dp.plem.PCPlus4M\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_16467_ _04470_ VGND VGND VPWR VPWR _01809_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_186_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18206_ _05570_ _05493_ VGND VGND VPWR VPWR _05571_ sky130_fd_sc_hd__or2_1
XFILLER_0_115_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15418_ _13425_ _13390_ _13317_ VGND VGND VPWR VPWR _13950_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_171_4598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19186_ _06487_ _06491_ VGND VGND VPWR VPWR _06498_ sky130_fd_sc_hd__nand2_1
X_31464_ clknet_leaf_75_clk rvcpu.dp.SrcBFW_Mux.y\[22\] VGND VGND VPWR VPWR rvcpu.dp.plem.WriteDataM\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_113_3203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16398_ net2065 _14428_ _14561_ VGND VGND VPWR VPWR _14565_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_3214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18137_ _05500_ _05501_ VGND VGND VPWR VPWR _05503_ sky130_fd_sc_hd__nor2_1
X_30415_ net753 _02150_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[31\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15349_ _13431_ _13526_ _13428_ _13737_ _13312_ VGND VGND VPWR VPWR _13885_ sky130_fd_sc_hd__a41o_1
X_31395_ clknet_leaf_50_clk _03098_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCE\[12\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f__10243_ clknet_0__10243_ VGND VGND VPWR VPWR clknet_1_0__leaf__10243_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_170_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_184_4904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold104 rvcpu.dp.plem.ALUResultM\[13\] VGND VGND VPWR VPWR net1254 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_184_4915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold115 rvcpu.dp.plem.ALUResultM\[29\] VGND VGND VPWR VPWR net1265 sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 rvcpu.dp.plem.ALUResultM\[20\] VGND VGND VPWR VPWR net1276 sky130_fd_sc_hd__dlygate4sd3_1
X_18068_ _05435_ VGND VGND VPWR VPWR _05436_ sky130_fd_sc_hd__buf_2
XFILLER_0_151_580 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30346_ net692 _02081_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[4\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold137 datamem.data_ram\[0\]\[3\] VGND VGND VPWR VPWR net1287 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__10174_ clknet_0__10174_ VGND VGND VPWR VPWR clknet_1_0__leaf__10174_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_223_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold148 rvcpu.dp.plem.ALUResultM\[16\] VGND VGND VPWR VPWR net1298 sky130_fd_sc_hd__dlygate4sd3_1
X_23238__886 clknet_1_1__leaf__10126_ VGND VGND VPWR VPWR net1012 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_74_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold159 datamem.data_ram\[46\]\[6\] VGND VGND VPWR VPWR net1309 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_145_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17019_ _04763_ VGND VGND VPWR VPWR _01526_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_74_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30277_ clknet_leaf_144_clk _02012_ VGND VGND VPWR VPWR datamem.data_ram\[58\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32016_ clknet_leaf_42_clk _03438_ VGND VGND VPWR VPWR rvcpu.dp.pcreg.q\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20030_ datamem.data_ram\[30\]\[26\] _06763_ _06766_ datamem.data_ram\[28\]\[26\]
+ VGND VGND VPWR VPWR _07324_ sky130_fd_sc_hd__o22a_1
XFILLER_0_106_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_193_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_3922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21981_ _08624_ _09211_ VGND VGND VPWR VPWR _09212_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_33_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32918_ clknet_leaf_91_clk _04340_ VGND VGND VPWR VPWR datamem.data_ram\[0\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_20932_ datamem.data_ram\[34\]\[22\] _07849_ _08221_ _07636_ VGND VGND VPWR VPWR
+ _08222_ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23974__510 clknet_1_0__leaf__10238_ VGND VGND VPWR VPWR net636 sky130_fd_sc_hd__inv_2
XFILLER_0_7_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32849_ clknet_leaf_234_clk _04271_ VGND VGND VPWR VPWR datamem.data_ram\[11\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_20863_ _08133_ _08137_ _08145_ _08152_ VGND VGND VPWR VPWR _08153_ sky130_fd_sc_hd__o211a_1
XFILLER_0_135_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22602_ _09528_ _09752_ _09426_ VGND VGND VPWR VPWR _09753_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_102_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26370_ _11517_ net1722 _11510_ _11519_ VGND VGND VPWR VPWR _03140_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_102_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20794_ datamem.data_ram\[32\]\[30\] _06990_ _08083_ _07636_ _07903_ VGND VGND VPWR
+ VPWR _08084_ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25321_ _10905_ VGND VGND VPWR VPWR _02705_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22533_ _09679_ _09683_ _09687_ _09491_ VGND VGND VPWR VPWR _01135_ sky130_fd_sc_hd__o31a_1
XFILLER_0_88_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_174_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25252_ _07077_ _10042_ _10044_ VGND VGND VPWR VPWR _10866_ sky130_fd_sc_hd__or3_1
XFILLER_0_151_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28040_ _09350_ _12345_ _12482_ VGND VGND VPWR VPWR _12483_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_161_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22464_ _09399_ VGND VGND VPWR VPWR _09622_ sky130_fd_sc_hd__clkbuf_4
X_22998__704 clknet_1_1__leaf__10084_ VGND VGND VPWR VPWR net830 sky130_fd_sc_hd__inv_2
XFILLER_0_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24203_ _09306_ net2257 _10270_ VGND VGND VPWR VPWR _10272_ sky130_fd_sc_hd__mux2_1
X_21415_ rvcpu.dp.rf.reg_file_arr\[24\]\[3\] rvcpu.dp.rf.reg_file_arr\[25\]\[3\] rvcpu.dp.rf.reg_file_arr\[26\]\[3\]
+ rvcpu.dp.rf.reg_file_arr\[27\]\[3\] _08549_ _08527_ VGND VGND VPWR VPWR _08674_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_45_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25183_ _10570_ _10640_ _10828_ VGND VGND VPWR VPWR _10829_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_32_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22395_ _09556_ VGND VGND VPWR VPWR _01128_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21346_ rvcpu.ALUResultE\[19\] rvcpu.ALUResultE\[21\] _08605_ _08607_ VGND VGND VPWR
+ VPWR _08608_ sky130_fd_sc_hd__or4_1
X_29991_ net361 _01726_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[14\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_28942_ _06591_ VGND VGND VPWR VPWR _12977_ sky130_fd_sc_hd__buf_8
Xhold660 datamem.data_ram\[34\]\[0\] VGND VGND VPWR VPWR net1810 sky130_fd_sc_hd__dlygate4sd3_1
X_21277_ _08532_ _08538_ VGND VGND VPWR VPWR _08539_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold671 rvcpu.dp.plfd.PCD\[13\] VGND VGND VPWR VPWR net1821 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_5_13__f_clk clknet_2_1_0_clk VGND VGND VPWR VPWR clknet_5_13__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_102_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold682 datamem.data_ram\[9\]\[6\] VGND VGND VPWR VPWR net1832 sky130_fd_sc_hd__dlygate4sd3_1
X_20228_ datamem.data_ram\[11\]\[3\] _06943_ _07520_ _07031_ VGND VGND VPWR VPWR _07521_
+ sky130_fd_sc_hd__a211o_1
Xhold693 rvcpu.dp.plfd.PCD\[23\] VGND VGND VPWR VPWR net1843 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28873_ _12940_ VGND VGND VPWR VPWR _04222_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_198_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27824_ _09297_ VGND VGND VPWR VPWR _12355_ sky130_fd_sc_hd__clkbuf_2
X_20159_ datamem.data_ram\[30\]\[27\] _06718_ _06696_ datamem.data_ram\[24\]\[27\]
+ _07451_ VGND VGND VPWR VPWR _07452_ sky130_fd_sc_hd__o221a_1
Xhold2050 datamem.data_ram\[25\]\[11\] VGND VGND VPWR VPWR net3200 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2061 datamem.data_ram\[46\]\[16\] VGND VGND VPWR VPWR net3211 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2072 datamem.data_ram\[6\]\[9\] VGND VGND VPWR VPWR net3222 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27755_ _12317_ VGND VGND VPWR VPWR _03727_ sky130_fd_sc_hd__clkbuf_1
X_22970__678 clknet_1_1__leaf__10082_ VGND VGND VPWR VPWR net804 sky130_fd_sc_hd__inv_2
Xhold2083 rvcpu.dp.rf.reg_file_arr\[29\]\[26\] VGND VGND VPWR VPWR net3233 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2094 datamem.data_ram\[44\]\[20\] VGND VGND VPWR VPWR net3244 sky130_fd_sc_hd__dlygate4sd3_1
X_24967_ _10398_ net2120 _10696_ VGND VGND VPWR VPWR _10703_ sky130_fd_sc_hd__mux2_1
Xhold1360 rvcpu.dp.rf.reg_file_arr\[4\]\[4\] VGND VGND VPWR VPWR net2510 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14720_ _13274_ VGND VGND VPWR VPWR _13275_ sky130_fd_sc_hd__buf_4
Xhold1371 datamem.data_ram\[3\]\[10\] VGND VGND VPWR VPWR net2521 sky130_fd_sc_hd__dlygate4sd3_1
X_26706_ _10818_ net3148 _11704_ VGND VGND VPWR VPWR _11708_ sky130_fd_sc_hd__mux2_1
Xhold1382 rvcpu.dp.rf.reg_file_arr\[28\]\[21\] VGND VGND VPWR VPWR net2532 sky130_fd_sc_hd__dlygate4sd3_1
X_23918_ clknet_1_1__leaf__10224_ VGND VGND VPWR VPWR _10226_ sky130_fd_sc_hd__buf_1
XANTENNA_500 _11157_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27686_ _12125_ net3080 _12280_ VGND VGND VPWR VPWR _12281_ sky130_fd_sc_hd__mux2_1
Xhold1393 rvcpu.dp.rf.reg_file_arr\[5\]\[22\] VGND VGND VPWR VPWR net2543 sky130_fd_sc_hd__dlygate4sd3_1
X_24898_ _10452_ net1911 _10659_ VGND VGND VPWR VPWR _10666_ sky130_fd_sc_hd__mux2_1
XFILLER_0_212_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_511 _13216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29425_ clknet_leaf_100_clk _01160_ VGND VGND VPWR VPWR datamem.data_ram\[5\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_522 _13257_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_1_1__f__10206_ clknet_0__10206_ VGND VGND VPWR VPWR clknet_1_1__leaf__10206_
+ sky130_fd_sc_hd__clkbuf_16
X_26637_ _11104_ VGND VGND VPWR VPWR _11665_ sky130_fd_sc_hd__buf_2
XANTENNA_533 rvcpu.dp.plmw.ReadDataW\[24\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14651_ _13222_ VGND VGND VPWR VPWR _13223_ sky130_fd_sc_hd__clkbuf_8
XANTENNA_544 _06753_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_555 _07845_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23381__1015 clknet_1_0__leaf__10140_ VGND VGND VPWR VPWR net1141 sky130_fd_sc_hd__inv_2
XFILLER_0_19_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_566 _14175_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_200_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29356_ clknet_leaf_145_clk _01091_ VGND VGND VPWR VPWR datamem.data_ram\[61\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__10137_ clknet_0__10137_ VGND VGND VPWR VPWR clknet_1_1__leaf__10137_
+ sky130_fd_sc_hd__clkbuf_16
X_17370_ _14151_ net2169 _04949_ VGND VGND VPWR VPWR _04950_ sky130_fd_sc_hd__mux2_1
X_23343__981 clknet_1_0__leaf__10136_ VGND VGND VPWR VPWR net1107 sky130_fd_sc_hd__inv_2
XFILLER_0_67_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26568_ _10668_ _10092_ _10998_ VGND VGND VPWR VPWR _11629_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_55_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28307_ _12454_ net3689 net72 VGND VGND VPWR VPWR _12627_ sky130_fd_sc_hd__mux2_1
X_23500__145 clknet_1_1__leaf__10161_ VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__inv_2
XFILLER_0_67_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16321_ _14523_ VGND VGND VPWR VPWR _01876_ sky130_fd_sc_hd__clkbuf_1
X_25519_ _10416_ _11010_ VGND VGND VPWR VPWR _11016_ sky130_fd_sc_hd__and2_1
X_29287_ _09321_ net2147 _13159_ VGND VGND VPWR VPWR _13165_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_188_5004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_188_5015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19040_ _06362_ _06364_ _06360_ VGND VGND VPWR VPWR _06370_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_164_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28238_ _12588_ VGND VGND VPWR VPWR _03939_ sky130_fd_sc_hd__clkbuf_1
X_16252_ net2076 _14486_ _14421_ VGND VGND VPWR VPWR _14487_ sky130_fd_sc_hd__mux2_1
X_23406__1021 clknet_1_1__leaf__10140_ VGND VGND VPWR VPWR net1147 sky130_fd_sc_hd__inv_2
XFILLER_0_35_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15203_ _13575_ _13744_ _13581_ VGND VGND VPWR VPWR _13745_ sky130_fd_sc_hd__a21oi_1
X_28169_ _12551_ VGND VGND VPWR VPWR _03907_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16183_ _13209_ VGND VGND VPWR VPWR _14440_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_152_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30200_ net554 _01935_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[8\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_15134_ _13533_ _13677_ _13678_ _13573_ _13438_ VGND VGND VPWR VPWR _13679_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_226_5911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31180_ clknet_leaf_209_clk _02883_ VGND VGND VPWR VPWR datamem.data_ram\[5\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_226_5922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_147_4022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15065_ _13540_ _13606_ _13609_ _13611_ VGND VGND VPWR VPWR _13612_ sky130_fd_sc_hd__or4_1
X_19942_ datamem.data_ram\[46\]\[18\] _06627_ _06803_ datamem.data_ram\[42\]\[18\]
+ VGND VGND VPWR VPWR _07236_ sky130_fd_sc_hd__o22a_1
X_30131_ net493 _01866_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[10\]\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_147_4033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_222_5819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30062_ net424 _01797_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[12\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19873_ datamem.data_ram\[29\]\[1\] _06969_ _06943_ datamem.data_ram\[27\]\[1\] _07031_
+ VGND VGND VPWR VPWR _07168_ sky130_fd_sc_hd__a221o_1
XFILLER_0_219_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_208_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18824_ _05497_ _06168_ _05809_ VGND VGND VPWR VPWR _06170_ sky130_fd_sc_hd__o21a_1
XFILLER_0_175_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_218_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18755_ _05311_ _05611_ _06091_ VGND VGND VPWR VPWR _06105_ sky130_fd_sc_hd__nand3_1
XFILLER_0_207_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15967_ _14320_ VGND VGND VPWR VPWR _02043_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_106_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17706_ _05127_ VGND VGND VPWR VPWR _01187_ sky130_fd_sc_hd__clkbuf_1
X_14918_ _13439_ _13464_ _13465_ _13467_ VGND VGND VPWR VPWR _13468_ sky130_fd_sc_hd__a2bb2o_1
X_18686_ _05419_ _06039_ VGND VGND VPWR VPWR _06040_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30964_ clknet_leaf_152_clk _02699_ VGND VGND VPWR VPWR datamem.data_ram\[3\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15898_ net2493 _13207_ _14275_ VGND VGND VPWR VPWR _14284_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_177_4741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_177_4752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32703_ clknet_leaf_185_clk _04125_ VGND VGND VPWR VPWR datamem.data_ram\[17\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_216_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17637_ net2424 _13206_ _05082_ VGND VGND VPWR VPWR _05091_ sky130_fd_sc_hd__mux2_1
X_14849_ _13399_ _13401_ VGND VGND VPWR VPWR _13402_ sky130_fd_sc_hd__nor2_4
X_30895_ clknet_leaf_150_clk _02630_ VGND VGND VPWR VPWR datamem.data_ram\[41\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_173_4638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32634_ clknet_leaf_273_clk _04056_ VGND VGND VPWR VPWR datamem.data_ram\[1\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_173_4649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17568_ _05054_ VGND VGND VPWR VPWR _01252_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_175_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19307_ _06602_ VGND VGND VPWR VPWR _06603_ sky130_fd_sc_hd__buf_8
XFILLER_0_46_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16519_ _04497_ VGND VGND VPWR VPWR _01784_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32565_ clknet_leaf_78_clk _03987_ VGND VGND VPWR VPWR datamem.data_ram\[22\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_17499_ _13204_ net3733 _05010_ VGND VGND VPWR VPWR _05018_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31516_ clknet_leaf_51_clk net1237 VGND VGND VPWR VPWR rvcpu.dp.plem.PCPlus4M\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_19238_ _06533_ _06530_ _06536_ _06527_ VGND VGND VPWR VPWR _06543_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_143_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_3770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32496_ clknet_leaf_3_clk _03918_ VGND VGND VPWR VPWR datamem.data_ram\[25\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19169_ _06473_ _06476_ VGND VGND VPWR VPWR _06483_ sky130_fd_sc_hd__nand2_1
XFILLER_0_186_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31447_ clknet_leaf_6_clk rvcpu.dp.SrcBFW_Mux.y\[5\] VGND VGND VPWR VPWR rvcpu.dp.plem.WriteDataM\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_76_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21200_ _08468_ _07920_ _07965_ _06580_ VGND VGND VPWR VPWR _08482_ sky130_fd_sc_hd__o22a_1
XFILLER_0_143_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_132_3667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22180_ _09351_ _09229_ _09361_ VGND VGND VPWR VPWR _09362_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_83_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_223_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_197_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31378_ clknet_leaf_22_clk _03081_ VGND VGND VPWR VPWR rvcpu.dp.plde.ImmExtE\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__10226_ clknet_0__10226_ VGND VGND VPWR VPWR clknet_1_0__leaf__10226_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_14_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21131_ datamem.data_ram\[32\]\[23\] datamem.data_ram\[33\]\[23\] datamem.data_ram\[34\]\[23\]
+ datamem.data_ram\[35\]\[23\] _07874_ _07820_ VGND VGND VPWR VPWR _08420_ sky130_fd_sc_hd__mux4_1
XFILLER_0_160_1344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30329_ net675 _02064_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[4\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_223_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__10157_ clknet_0__10157_ VGND VGND VPWR VPWR clknet_1_0__leaf__10157_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_1_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21062_ _06599_ _08347_ _08350_ _07903_ VGND VGND VPWR VPWR _08351_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_35_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__10088_ clknet_0__10088_ VGND VGND VPWR VPWR clknet_1_0__leaf__10088_
+ sky130_fd_sc_hd__clkbuf_16
X_20013_ datamem.data_ram\[51\]\[2\] _06941_ _06947_ datamem.data_ram\[49\]\[2\] _06600_
+ VGND VGND VPWR VPWR _07307_ sky130_fd_sc_hd__a221o_1
XFILLER_0_226_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25870_ rvcpu.dp.pcreg.q\[29\] _11239_ rvcpu.dp.pcreg.q\[30\] VGND VGND VPWR VPWR
+ _11248_ sky130_fd_sc_hd__a21oi_1
X_23441__92 clknet_1_0__leaf__10155_ VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__inv_2
X_24041__570 clknet_1_1__leaf__10245_ VGND VGND VPWR VPWR net696 sky130_fd_sc_hd__inv_2
XFILLER_0_214_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24821_ _10624_ VGND VGND VPWR VPWR _02486_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_193_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27540_ _12202_ VGND VGND VPWR VPWR _03627_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21964_ rvcpu.dp.rf.reg_file_arr\[24\]\[31\] rvcpu.dp.rf.reg_file_arr\[25\]\[31\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[31\] rvcpu.dp.rf.reg_file_arr\[27\]\[31\] _08548_
+ _08552_ VGND VGND VPWR VPWR _09195_ sky130_fd_sc_hd__mux4_2
X_24752_ _10585_ VGND VGND VPWR VPWR _02456_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_179_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20915_ datamem.data_ram\[28\]\[22\] datamem.data_ram\[29\]\[22\] _07827_ VGND VGND
+ VPWR VPWR _08205_ sky130_fd_sc_hd__mux2_1
X_27471_ _12091_ net2446 net83 VGND VGND VPWR VPWR _12165_ sky130_fd_sc_hd__mux2_1
X_24683_ _10548_ VGND VGND VPWR VPWR _02424_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_194_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21895_ rvcpu.dp.rf.reg_file_arr\[28\]\[27\] rvcpu.dp.rf.reg_file_arr\[30\]\[27\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[27\] rvcpu.dp.rf.reg_file_arr\[31\]\[27\] _08552_
+ _08687_ VGND VGND VPWR VPWR _09130_ sky130_fd_sc_hd__mux4_1
XFILLER_0_16_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29210_ _13018_ net1566 _13122_ _13124_ VGND VGND VPWR VPWR _04375_ sky130_fd_sc_hd__a31o_1
XFILLER_0_193_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26422_ _06438_ _11539_ _11529_ _11184_ _11558_ VGND VGND VPWR VPWR _11559_ sky130_fd_sc_hd__a221o_1
X_23634_ _10183_ VGND VGND VPWR VPWR _01740_ sky130_fd_sc_hd__clkbuf_1
X_20846_ datamem.data_ram\[22\]\[14\] _06629_ _06664_ datamem.data_ram\[21\]\[14\]
+ _08135_ VGND VGND VPWR VPWR _08136_ sky130_fd_sc_hd__o221a_1
XFILLER_0_193_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29141_ _09272_ net3600 net39 VGND VGND VPWR VPWR _13087_ sky130_fd_sc_hd__mux2_1
X_26353_ _07028_ _10932_ _11494_ VGND VGND VPWR VPWR _11509_ sky130_fd_sc_hd__or3_1
XFILLER_0_92_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20777_ _08063_ _08064_ _08065_ _08066_ VGND VGND VPWR VPWR _08067_ sky130_fd_sc_hd__o31a_1
XFILLER_0_9_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25304_ _10766_ net2666 _10887_ VGND VGND VPWR VPWR _10895_ sky130_fd_sc_hd__mux2_1
X_22516_ rvcpu.dp.rf.reg_file_arr\[16\]\[11\] rvcpu.dp.rf.reg_file_arr\[17\]\[11\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[11\] rvcpu.dp.rf.reg_file_arr\[19\]\[11\] _09445_
+ _09447_ VGND VGND VPWR VPWR _09671_ sky130_fd_sc_hd__mux4_1
XFILLER_0_36_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26284_ _11474_ VGND VGND VPWR VPWR _03099_ sky130_fd_sc_hd__clkbuf_1
X_29072_ _13050_ VGND VGND VPWR VPWR _04311_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28023_ _12430_ net4294 _12473_ VGND VGND VPWR VPWR _12474_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25235_ _10838_ _10640_ _10828_ VGND VGND VPWR VPWR _10857_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_91_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22447_ _09528_ _09605_ _09426_ VGND VGND VPWR VPWR _09606_ sky130_fd_sc_hd__a21o_1
XFILLER_0_162_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25166_ _10817_ VGND VGND VPWR VPWR _02638_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22378_ _09391_ _09539_ VGND VGND VPWR VPWR _09540_ sky130_fd_sc_hd__or2_1
X_21329_ rvcpu.dp.plfd.InstrD\[23\] _08582_ rvcpu.dp.plde.RdE\[4\] _08589_ _08590_
+ VGND VGND VPWR VPWR _08591_ sky130_fd_sc_hd__a221o_1
X_25097_ _10058_ _10779_ _10781_ net1616 VGND VGND VPWR VPWR _02605_ sky130_fd_sc_hd__a22o_1
X_29974_ net344 _01709_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[14\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28925_ _09350_ _10960_ _12886_ VGND VGND VPWR VPWR _12968_ sky130_fd_sc_hd__a21oi_4
Xhold490 datamem.data_ram\[1\]\[7\] VGND VGND VPWR VPWR net1640 sky130_fd_sc_hd__dlygate4sd3_1
X_16870_ _04683_ VGND VGND VPWR VPWR _04684_ sky130_fd_sc_hd__clkbuf_4
X_28856_ _12931_ VGND VGND VPWR VPWR _04214_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_217_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15821_ net2163 _13198_ _14236_ VGND VGND VPWR VPWR _14242_ sky130_fd_sc_hd__mux2_1
X_27807_ _10598_ _12345_ _12260_ VGND VGND VPWR VPWR _12346_ sky130_fd_sc_hd__a21oi_1
X_28787_ _12766_ net2787 _12887_ VGND VGND VPWR VPWR _12895_ sky130_fd_sc_hd__mux2_1
X_25999_ net14 _11317_ VGND VGND VPWR VPWR _11324_ sky130_fd_sc_hd__or2_1
XFILLER_0_126_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18540_ _05626_ _05621_ _05622_ _05574_ _05682_ _05579_ VGND VGND VPWR VPWR _05901_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_172_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27738_ _12308_ VGND VGND VPWR VPWR _03719_ sky130_fd_sc_hd__clkbuf_1
X_15752_ _14141_ net3082 _14199_ VGND VGND VPWR VPWR _14205_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1190 datamem.data_ram\[42\]\[22\] VGND VGND VPWR VPWR net2340 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14703_ rvcpu.dp.plmw.ALUResultW\[5\] rvcpu.dp.plmw.ReadDataW\[5\] rvcpu.dp.plmw.PCPlus4W\[5\]
+ rvcpu.dp.plmw.lAuiPCW\[5\] _13192_ _13193_ VGND VGND VPWR VPWR _13262_ sky130_fd_sc_hd__mux4_2
XFILLER_0_169_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18471_ _05363_ _05830_ _05833_ _05781_ VGND VGND VPWR VPWR _05834_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_197_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27669_ _12271_ VGND VGND VPWR VPWR _03687_ sky130_fd_sc_hd__clkbuf_1
X_15683_ _14159_ VGND VGND VPWR VPWR _02174_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_330 _14457_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_197_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_414 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_341 _14468_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_352 rvcpu.ALUResultE\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29408_ clknet_leaf_290_clk _01143_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD2E\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_17422_ _04977_ VGND VGND VPWR VPWR _01329_ sky130_fd_sc_hd__clkbuf_1
X_24018__550 clknet_1_0__leaf__10242_ VGND VGND VPWR VPWR net676 sky130_fd_sc_hd__inv_2
XANTENNA_363 rvcpu.dp.SrcBFW_Mux.y\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14634_ _13209_ VGND VGND VPWR VPWR _13210_ sky130_fd_sc_hd__buf_4
X_30680_ clknet_leaf_96_clk _02415_ VGND VGND VPWR VPWR datamem.data_ram\[4\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_374 rvcpu.dp.plem.ALUResultM\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23498__144 clknet_1_1__leaf__10160_ VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_215_5645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_215_5656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_385 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_215_5667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_396 _05886_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17353_ _14135_ net3223 _04938_ VGND VGND VPWR VPWR _04941_ sky130_fd_sc_hd__mux2_1
X_29339_ clknet_leaf_174_clk _01074_ VGND VGND VPWR VPWR datamem.data_ram\[62\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_222_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16304_ net2599 _14470_ _14511_ VGND VGND VPWR VPWR _14515_ sky130_fd_sc_hd__mux2_1
X_32350_ clknet_leaf_82_clk _03772_ VGND VGND VPWR VPWR datamem.data_ram\[30\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_222_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17284_ _04904_ VGND VGND VPWR VPWR _01402_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31301_ clknet_leaf_48_clk _03004_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCPlus4E\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_19023_ _06354_ rvcpu.dp.plde.ImmExtE\[0\] _06355_ VGND VGND VPWR VPWR _06356_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16235_ _14475_ VGND VGND VPWR VPWR _01922_ sky130_fd_sc_hd__clkbuf_1
X_32281_ clknet_leaf_241_clk _03703_ VGND VGND VPWR VPWR datamem.data_ram\[33\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload305 clknet_1_0__leaf__10198_ VGND VGND VPWR VPWR clkload305/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload13 clknet_5_15__leaf_clk VGND VGND VPWR VPWR clkload13/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_141_826 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload316 clknet_1_0__leaf__10176_ VGND VGND VPWR VPWR clkload316/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_144_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload24 clknet_5_29__leaf_clk VGND VGND VPWR VPWR clkload24/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_125_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload327 clknet_1_0__leaf__10267_ VGND VGND VPWR VPWR clkload327/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload35 clknet_leaf_18_clk VGND VGND VPWR VPWR clkload35/Y sky130_fd_sc_hd__clkinv_1
XFILLER_0_144_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload338 clknet_1_0__leaf__10108_ VGND VGND VPWR VPWR clkload338/X sky130_fd_sc_hd__clkbuf_8
X_31232_ clknet_leaf_42_clk _02935_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCD\[21\] sky130_fd_sc_hd__dfxtp_1
Xclkload46 clknet_leaf_8_clk VGND VGND VPWR VPWR clkload46/Y sky130_fd_sc_hd__inv_6
Xclkload349 clknet_1_0__leaf__10102_ VGND VGND VPWR VPWR clkload349/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_23_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16166_ net2254 _14428_ _14422_ VGND VGND VPWR VPWR _14429_ sky130_fd_sc_hd__mux2_1
Xclkload57 clknet_leaf_3_clk VGND VGND VPWR VPWR clkload57/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_51_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_224_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload68 clknet_leaf_66_clk VGND VGND VPWR VPWR clkload68/Y sky130_fd_sc_hd__clkinvlp_2
Xclkload79 clknet_leaf_41_clk VGND VGND VPWR VPWR clkload79/Y sky130_fd_sc_hd__inv_8
X_15117_ _13646_ _13653_ _13655_ _13661_ VGND VGND VPWR VPWR _13662_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_71_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31163_ clknet_leaf_28_clk rvcpu.ALUResultE\[22\] VGND VGND VPWR VPWR rvcpu.dp.plem.ALUResultM\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16097_ _14390_ VGND VGND VPWR VPWR _01975_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_166_4475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30114_ net476 _01849_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[10\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_15048_ _13588_ _13591_ _13594_ VGND VGND VPWR VPWR _13595_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_166_4486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19925_ datamem.data_ram\[48\]\[17\] _06807_ _06789_ datamem.data_ram\[49\]\[17\]
+ VGND VGND VPWR VPWR _07220_ sky130_fd_sc_hd__o22a_1
XFILLER_0_55_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31094_ clknet_leaf_273_clk _02829_ VGND VGND VPWR VPWR datamem.data_ram\[9\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2808 rvcpu.dp.rf.reg_file_arr\[29\]\[27\] VGND VGND VPWR VPWR net3958 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_167_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2819 datamem.data_ram\[40\]\[19\] VGND VGND VPWR VPWR net3969 sky130_fd_sc_hd__dlygate4sd3_1
X_19856_ datamem.data_ram\[63\]\[1\] _07125_ _07147_ _07150_ VGND VGND VPWR VPWR _07151_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_208_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30045_ net407 _01780_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[12\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_177_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_179_4803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18807_ _05504_ _06134_ _06153_ _05568_ VGND VGND VPWR VPWR _06154_ sky130_fd_sc_hd__o211a_1
X_19787_ datamem.data_ram\[47\]\[9\] _06672_ _07080_ _07081_ VGND VGND VPWR VPWR _07082_
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_30_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16999_ net2293 _14482_ _04742_ VGND VGND VPWR VPWR _04752_ sky130_fd_sc_hd__mux2_1
XFILLER_0_207_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18738_ _05610_ _05330_ VGND VGND VPWR VPWR _06089_ sky130_fd_sc_hd__nor2_1
XFILLER_0_222_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31996_ clknet_leaf_128_clk _03418_ VGND VGND VPWR VPWR datamem.data_ram\[31\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_125_3493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30947_ clknet_leaf_86_clk _02682_ VGND VGND VPWR VPWR datamem.data_ram\[3\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_18669_ _05990_ _05824_ _05829_ _06022_ _06023_ VGND VGND VPWR VPWR _06024_ sky130_fd_sc_hd__o221a_1
XFILLER_0_149_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20700_ datamem.data_ram\[6\]\[5\] _07127_ _07989_ _07990_ VGND VGND VPWR VPWR _07991_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_153_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21680_ rvcpu.dp.rf.reg_file_arr\[4\]\[15\] rvcpu.dp.rf.reg_file_arr\[5\]\[15\] rvcpu.dp.rf.reg_file_arr\[6\]\[15\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[15\] _08687_ _08856_ VGND VGND VPWR VPWR _08927_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_138_3810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30878_ clknet_leaf_281_clk _02613_ VGND VGND VPWR VPWR datamem.data_ram\[42\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_175_255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32617_ clknet_leaf_251_clk _04039_ VGND VGND VPWR VPWR datamem.data_ram\[20\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_20631_ datamem.data_ram\[2\]\[29\] _06612_ _06779_ datamem.data_ram\[0\]\[29\] _07921_
+ VGND VGND VPWR VPWR _07922_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_28_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_3707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_1277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_178_Right_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_134_3718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20562_ _06603_ _07848_ _07852_ VGND VGND VPWR VPWR _07853_ sky130_fd_sc_hd__and3_1
XFILLER_0_149_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32548_ clknet_leaf_253_clk _03970_ VGND VGND VPWR VPWR datamem.data_ram\[23\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload7 clknet_5_8__leaf_clk VGND VGND VPWR VPWR clkload7/Y sky130_fd_sc_hd__inv_8
XFILLER_0_132_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22301_ _09465_ VGND VGND VPWR VPWR _09466_ sky130_fd_sc_hd__buf_4
XFILLER_0_190_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23281_ clknet_1_0__leaf__10130_ VGND VGND VPWR VPWR _10131_ sky130_fd_sc_hd__buf_1
XFILLER_0_73_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20493_ _06915_ _07781_ _07646_ _07277_ VGND VGND VPWR VPWR _07785_ sky130_fd_sc_hd__o22a_1
X_32479_ clknet_leaf_274_clk _03901_ VGND VGND VPWR VPWR datamem.data_ram\[26\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25020_ _10733_ net3792 net100 VGND VGND VPWR VPWR _10734_ sky130_fd_sc_hd__mux2_1
X_22232_ rvcpu.dp.plfd.InstrD\[22\] VGND VGND VPWR VPWR _09398_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_95_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22163_ _09298_ net2916 _09352_ VGND VGND VPWR VPWR _09353_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21114_ datamem.data_ram\[30\]\[7\] _06950_ _06923_ datamem.data_ram\[31\]\[7\] _08402_
+ VGND VGND VPWR VPWR _08403_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_58_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26971_ _11863_ net1521 _11865_ _11869_ VGND VGND VPWR VPWR _03391_ sky130_fd_sc_hd__a31o_1
X_22094_ _09306_ net2300 _09302_ VGND VGND VPWR VPWR _09307_ sky130_fd_sc_hd__mux2_1
X_28710_ _12694_ net2988 _12850_ VGND VGND VPWR VPWR _12854_ sky130_fd_sc_hd__mux2_1
X_25922_ net1291 _11279_ VGND VGND VPWR VPWR _11281_ sky130_fd_sc_hd__or2_1
X_21045_ datamem.data_ram\[2\]\[31\] datamem.data_ram\[3\]\[31\] _06933_ VGND VGND
+ VPWR VPWR _08334_ sky130_fd_sc_hd__mux2_1
X_29690_ net1036 _01425_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[23\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_54_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28641_ _12817_ VGND VGND VPWR VPWR _04113_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_214_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25853_ rvcpu.dp.pcreg.q\[27\] rvcpu.dp.pcreg.q\[26\] _11226_ VGND VGND VPWR VPWR
+ _11234_ sky130_fd_sc_hd__and3_1
X_23405__1020 clknet_1_1__leaf__10140_ VGND VGND VPWR VPWR net1146 sky130_fd_sc_hd__inv_2
XFILLER_0_214_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24804_ _10615_ VGND VGND VPWR VPWR _02478_ sky130_fd_sc_hd__clkbuf_1
X_28572_ _12780_ VGND VGND VPWR VPWR _04081_ sky130_fd_sc_hd__clkbuf_1
X_25784_ _11178_ _11179_ _11149_ VGND VGND VPWR VPWR _11180_ sky130_fd_sc_hd__o21ai_1
X_27523_ _12193_ VGND VGND VPWR VPWR _03619_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24735_ _10576_ VGND VGND VPWR VPWR _02448_ sky130_fd_sc_hd__clkbuf_1
X_21947_ rvcpu.dp.rf.reg_file_arr\[20\]\[30\] rvcpu.dp.rf.reg_file_arr\[21\]\[30\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[30\] rvcpu.dp.rf.reg_file_arr\[23\]\[30\] _08535_
+ _08533_ VGND VGND VPWR VPWR _09179_ sky130_fd_sc_hd__mux4_1
XFILLER_0_16_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27454_ _09287_ VGND VGND VPWR VPWR _12155_ sky130_fd_sc_hd__clkbuf_2
X_24666_ _10416_ _10532_ VGND VGND VPWR VPWR _10539_ sky130_fd_sc_hd__and2_1
X_21878_ rvcpu.dp.rf.reg_file_arr\[24\]\[26\] rvcpu.dp.rf.reg_file_arr\[25\]\[26\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[26\] rvcpu.dp.rf.reg_file_arr\[27\]\[26\] _08536_
+ _08693_ VGND VGND VPWR VPWR _09114_ sky130_fd_sc_hd__mux4_1
XFILLER_0_139_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26405_ _06404_ _11522_ _11526_ _11167_ _11546_ VGND VGND VPWR VPWR _11547_ sky130_fd_sc_hd__a221o_1
XFILLER_0_65_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20829_ datamem.data_ram\[8\]\[30\] _06647_ _06782_ datamem.data_ram\[9\]\[30\] VGND
+ VGND VPWR VPWR _08119_ sky130_fd_sc_hd__o22a_1
X_27385_ _10733_ net3863 net86 VGND VGND VPWR VPWR _12112_ sky130_fd_sc_hd__mux2_1
X_24597_ _10499_ VGND VGND VPWR VPWR _02387_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_194_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29124_ _09235_ net4129 _13076_ VGND VGND VPWR VPWR _13078_ sky130_fd_sc_hd__mux2_1
X_26336_ _11501_ net1724 _11496_ _11503_ VGND VGND VPWR VPWR _03122_ sky130_fd_sc_hd__a31o_1
XFILLER_0_167_1328 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_145_Right_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_210_5531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_210_5542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29055_ _13041_ VGND VGND VPWR VPWR _04303_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26267_ _11465_ VGND VGND VPWR VPWR _03091_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_190_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28006_ _12355_ net4255 net97 VGND VGND VPWR VPWR _12465_ sky130_fd_sc_hd__mux2_1
X_23651__251 clknet_1_1__leaf__10181_ VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__inv_2
X_16020_ net2150 _13173_ _14349_ VGND VGND VPWR VPWR _14350_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25218_ _10838_ _10630_ _10828_ VGND VGND VPWR VPWR _10848_ sky130_fd_sc_hd__a21oi_4
X_26198_ rvcpu.c.ad.opb5 _11436_ _11377_ VGND VGND VPWR VPWR _11437_ sky130_fd_sc_hd__and3_1
XFILLER_0_66_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24048__576 clknet_1_1__leaf__10246_ VGND VGND VPWR VPWR net702 sky130_fd_sc_hd__inv_2
X_25149_ _10760_ net3999 _10802_ VGND VGND VPWR VPWR _10807_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17971_ rvcpu.dp.plde.RD1E\[7\] _05292_ _05341_ VGND VGND VPWR VPWR _05342_ sky130_fd_sc_hd__o21a_2
X_29957_ net327 _01692_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[15\]\[16\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_208_5482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22976__684 clknet_1_0__leaf__10082_ VGND VGND VPWR VPWR net810 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_208_5493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19710_ datamem.data_ram\[22\]\[0\] _06951_ _06936_ datamem.data_ram\[16\]\[0\] _06741_
+ VGND VGND VPWR VPWR _07006_ sky130_fd_sc_hd__a221o_1
XFILLER_0_218_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16922_ _04711_ VGND VGND VPWR VPWR _01579_ sky130_fd_sc_hd__clkbuf_1
X_28908_ _09350_ _10997_ _12886_ VGND VGND VPWR VPWR _12959_ sky130_fd_sc_hd__a21oi_4
X_29888_ net266 _01623_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[17\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_161_4350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19641_ _06936_ VGND VGND VPWR VPWR _06937_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_161_4361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28839_ _12922_ VGND VGND VPWR VPWR _04206_ sky130_fd_sc_hd__clkbuf_1
X_16853_ net2179 _14472_ _04670_ VGND VGND VPWR VPWR _04675_ sky130_fd_sc_hd__mux2_1
X_23420__73 clknet_1_0__leaf__10153_ VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__inv_2
XFILLER_0_102_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15804_ _14193_ net3314 _14198_ VGND VGND VPWR VPWR _14232_ sky130_fd_sc_hd__mux2_1
X_31850_ clknet_leaf_110_clk _03304_ VGND VGND VPWR VPWR datamem.data_ram\[61\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_19572_ datamem.data_ram\[2\]\[8\] _06804_ _06837_ datamem.data_ram\[0\]\[8\] _06867_
+ VGND VGND VPWR VPWR _06868_ sky130_fd_sc_hd__o221a_1
X_16784_ _04638_ VGND VGND VPWR VPWR _01652_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_217_5707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18523_ _05584_ _05582_ _05583_ VGND VGND VPWR VPWR _05884_ sky130_fd_sc_hd__or3_1
X_30801_ clknet_leaf_220_clk _02536_ VGND VGND VPWR VPWR datamem.data_ram\[45\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23506__151 clknet_1_0__leaf__10161_ VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__inv_2
X_15735_ _14194_ VGND VGND VPWR VPWR _02157_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31781_ clknet_leaf_278_clk _03235_ VGND VGND VPWR VPWR datamem.data_ram\[6\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_201_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18454_ _05389_ _05729_ _05808_ _05396_ _05816_ VGND VGND VPWR VPWR _05817_ sky130_fd_sc_hd__a221o_1
X_30732_ clknet_leaf_199_clk _02467_ VGND VGND VPWR VPWR datamem.data_ram\[48\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15666_ _14147_ net4124 _14131_ VGND VGND VPWR VPWR _14148_ sky130_fd_sc_hd__mux2_1
XANTENNA_160 _08549_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_171 _08744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_201_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17405_ _14187_ net3872 _04960_ VGND VGND VPWR VPWR _04968_ sky130_fd_sc_hd__mux2_1
XANTENNA_182 _09024_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14617_ rvcpu.dp.plmw.ALUResultW\[26\] rvcpu.dp.plmw.ReadDataW\[26\] rvcpu.dp.plmw.PCPlus4W\[26\]
+ rvcpu.dp.plmw.lAuiPCW\[26\] _13192_ _13193_ VGND VGND VPWR VPWR _13197_ sky130_fd_sc_hd__mux4_2
XANTENNA_193 _09309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18385_ _05748_ VGND VGND VPWR VPWR _05749_ sky130_fd_sc_hd__clkbuf_4
X_30663_ clknet_leaf_149_clk _02398_ VGND VGND VPWR VPWR datamem.data_ram\[50\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15597_ _14106_ VGND VGND VPWR VPWR _02207_ sky130_fd_sc_hd__clkbuf_1
X_32402_ clknet_leaf_286_clk _03824_ VGND VGND VPWR VPWR datamem.data_ram\[29\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17336_ _04931_ VGND VGND VPWR VPWR _01377_ sky130_fd_sc_hd__clkbuf_1
X_30594_ clknet_leaf_118_clk _02329_ VGND VGND VPWR VPWR datamem.data_ram\[53\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_112_Right_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32333_ clknet_leaf_249_clk _03755_ VGND VGND VPWR VPWR datamem.data_ram\[31\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_17267_ _04894_ VGND VGND VPWR VPWR _01409_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload102 clknet_leaf_88_clk VGND VGND VPWR VPWR clkload102/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload113 clknet_leaf_103_clk VGND VGND VPWR VPWR clkload113/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_12_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19006_ _05290_ _05647_ _06055_ VGND VGND VPWR VPWR _06340_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_12_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload124 clknet_leaf_251_clk VGND VGND VPWR VPWR clkload124/Y sky130_fd_sc_hd__clkinv_4
X_16218_ _14421_ VGND VGND VPWR VPWR _14464_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_168_4526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23849__413 clknet_1_1__leaf__10208_ VGND VGND VPWR VPWR net539 sky130_fd_sc_hd__inv_2
Xclkload135 clknet_leaf_239_clk VGND VGND VPWR VPWR clkload135/Y sky130_fd_sc_hd__bufinv_16
X_32264_ clknet_leaf_275_clk _03686_ VGND VGND VPWR VPWR datamem.data_ram\[34\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_168_4537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17198_ _14185_ net2956 _04851_ VGND VGND VPWR VPWR _04858_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload146 clknet_leaf_259_clk VGND VGND VPWR VPWR clkload146/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_144_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload157 clknet_leaf_284_clk VGND VGND VPWR VPWR clkload157/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_144_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload168 clknet_leaf_269_clk VGND VGND VPWR VPWR clkload168/Y sky130_fd_sc_hd__clkinv_4
X_31215_ clknet_leaf_37_clk _02918_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCD\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16149_ _14417_ VGND VGND VPWR VPWR _01950_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload179 clknet_leaf_235_clk VGND VGND VPWR VPWR clkload179/Y sky130_fd_sc_hd__inv_6
XFILLER_0_11_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32195_ clknet_leaf_210_clk _03617_ VGND VGND VPWR VPWR datamem.data_ram\[36\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_90_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31146_ clknet_leaf_63_clk rvcpu.ALUResultE\[5\] VGND VGND VPWR VPWR rvcpu.dp.plem.ALUResultM\[5\]
+ sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_90_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2605 rvcpu.dp.rf.reg_file_arr\[2\]\[15\] VGND VGND VPWR VPWR net3755 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2616 rvcpu.dp.rf.reg_file_arr\[14\]\[7\] VGND VGND VPWR VPWR net3766 sky130_fd_sc_hd__dlygate4sd3_1
X_19908_ _07023_ VGND VGND VPWR VPWR _07203_ sky130_fd_sc_hd__clkbuf_8
X_31077_ clknet_leaf_101_clk _02812_ VGND VGND VPWR VPWR datamem.data_ram\[20\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold19 rvcpu.dp.plem.lAuiPCM\[4\] VGND VGND VPWR VPWR net1169 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_127_3533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2627 rvcpu.dp.rf.reg_file_arr\[15\]\[22\] VGND VGND VPWR VPWR net3777 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_127_3544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2638 datamem.data_ram\[36\]\[26\] VGND VGND VPWR VPWR net3788 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1904 datamem.data_ram\[43\]\[15\] VGND VGND VPWR VPWR net3054 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2649 datamem.data_ram\[44\]\[10\] VGND VGND VPWR VPWR net3799 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_127_3555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1915 datamem.data_ram\[32\]\[29\] VGND VGND VPWR VPWR net3065 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30028_ net390 _01763_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[13\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19839_ datamem.data_ram\[47\]\[1\] _06993_ _06976_ datamem.data_ram\[44\]\[1\] VGND
+ VGND VPWR VPWR _07134_ sky130_fd_sc_hd__a22o_1
Xhold1926 datamem.data_ram\[24\]\[15\] VGND VGND VPWR VPWR net3076 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1937 datamem.data_ram\[36\]\[10\] VGND VGND VPWR VPWR net3087 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1948 datamem.data_ram\[49\]\[19\] VGND VGND VPWR VPWR net3098 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1959 rvcpu.dp.rf.reg_file_arr\[28\]\[6\] VGND VGND VPWR VPWR net3109 sky130_fd_sc_hd__dlygate4sd3_1
X_22850_ rvcpu.dp.rf.reg_file_arr\[16\]\[29\] rvcpu.dp.rf.reg_file_arr\[17\]\[29\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[29\] rvcpu.dp.rf.reg_file_arr\[19\]\[29\] _09517_
+ _09513_ VGND VGND VPWR VPWR _09987_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_190_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21801_ rvcpu.dp.rf.reg_file_arr\[20\]\[22\] rvcpu.dp.rf.reg_file_arr\[21\]\[22\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[22\] rvcpu.dp.rf.reg_file_arr\[23\]\[22\] _08516_
+ _08518_ VGND VGND VPWR VPWR _09041_ sky130_fd_sc_hd__mux4_1
XFILLER_0_91_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22781_ rvcpu.dp.rf.reg_file_arr\[24\]\[25\] rvcpu.dp.rf.reg_file_arr\[25\]\[25\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[25\] rvcpu.dp.rf.reg_file_arr\[27\]\[25\] _09463_
+ _09637_ VGND VGND VPWR VPWR _09922_ sky130_fd_sc_hd__mux4_1
XFILLER_0_155_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31979_ clknet_leaf_151_clk _03401_ VGND VGND VPWR VPWR datamem.data_ram\[53\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24520_ _10454_ datamem.data_ram\[52\]\[23\] _10440_ VGND VGND VPWR VPWR _10455_
+ sky130_fd_sc_hd__mux2_1
X_21732_ _08795_ _08971_ _08973_ _08975_ VGND VGND VPWR VPWR _08976_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_91_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24451_ _10413_ _10406_ VGND VGND VPWR VPWR _10414_ sky130_fd_sc_hd__and2_1
XFILLER_0_164_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21663_ _08692_ _08908_ _08910_ VGND VGND VPWR VPWR _08911_ sky130_fd_sc_hd__a21o_1
XFILLER_0_143_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20614_ datamem.data_ram\[26\]\[13\] _06802_ _06661_ datamem.data_ram\[29\]\[13\]
+ VGND VGND VPWR VPWR _07905_ sky130_fd_sc_hd__o22a_1
X_27170_ _11918_ VGND VGND VPWR VPWR _11991_ sky130_fd_sc_hd__buf_2
X_24382_ _09240_ net4291 _10367_ VGND VGND VPWR VPWR _10370_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21594_ _08833_ _08838_ _08845_ _08625_ VGND VGND VPWR VPWR _01038_ sky130_fd_sc_hd__o31a_1
XFILLER_0_47_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26121_ net1650 _11386_ VGND VGND VPWR VPWR _11396_ sky130_fd_sc_hd__and2_1
XFILLER_0_145_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20545_ _07835_ VGND VGND VPWR VPWR _07836_ sky130_fd_sc_hd__buf_8
XFILLER_0_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_140_clk clknet_5_31__leaf_clk VGND VGND VPWR VPWR clknet_leaf_140_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_145_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_104_Left_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_229_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26052_ _11083_ _11351_ VGND VGND VPWR VPWR _11355_ sky130_fd_sc_hd__and2_1
XFILLER_0_132_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20476_ datamem.data_ram\[32\]\[20\] _06779_ _07764_ _07767_ VGND VGND VPWR VPWR
+ _07768_ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25003_ _10722_ VGND VGND VPWR VPWR _02570_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_1247 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22215_ _08595_ VGND VGND VPWR VPWR _09381_ sky130_fd_sc_hd__buf_4
X_23195_ _10118_ VGND VGND VPWR VPWR _01366_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29811_ net1149 _01546_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[1\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_22146_ _09273_ net2215 net62 VGND VGND VPWR VPWR _09343_ sky130_fd_sc_hd__mux2_1
X_29742_ net1088 _01477_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[21\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26954_ _11803_ _11854_ VGND VGND VPWR VPWR _11859_ sky130_fd_sc_hd__and2_1
X_22077_ _09291_ net1875 _09270_ VGND VGND VPWR VPWR _09292_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_1023 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25905_ net1852 _11263_ VGND VGND VPWR VPWR _11271_ sky130_fd_sc_hd__or2_1
X_21028_ datamem.data_ram\[26\]\[31\] _06802_ _08312_ _08316_ VGND VGND VPWR VPWR
+ _08317_ sky130_fd_sc_hd__o211a_1
XFILLER_0_195_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29673_ net1019 _01408_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[23\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_26885_ _11684_ _11810_ VGND VGND VPWR VPWR _11815_ sky130_fd_sc_hd__and2_1
XFILLER_0_214_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_113_Left_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23681__277 clknet_1_0__leaf__10194_ VGND VGND VPWR VPWR net403 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_76_Right_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28624_ _12808_ VGND VGND VPWR VPWR _04105_ sky130_fd_sc_hd__clkbuf_1
X_25836_ _11220_ VGND VGND VPWR VPWR _02905_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_214_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_214_Right_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_198_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28555_ _12771_ VGND VGND VPWR VPWR _04073_ sky130_fd_sc_hd__clkbuf_1
X_25767_ _11165_ _11166_ _11157_ VGND VGND VPWR VPWR _11167_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_195_5180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15520_ _13504_ _13831_ _13577_ _13538_ VGND VGND VPWR VPWR _14047_ sky130_fd_sc_hd__a31o_1
X_27506_ _12184_ VGND VGND VPWR VPWR _03611_ sky130_fd_sc_hd__clkbuf_1
X_24718_ _10476_ net3197 net59 VGND VGND VPWR VPWR _10567_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_201_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28486_ _06587_ VGND VGND VPWR VPWR _12727_ sky130_fd_sc_hd__buf_2
XFILLER_0_70_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25698_ _11104_ VGND VGND VPWR VPWR _11121_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_191_5077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_191_5088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15451_ _13308_ _13565_ _13832_ VGND VGND VPWR VPWR _13981_ sky130_fd_sc_hd__o21ai_1
X_27437_ _12142_ net3521 net84 VGND VGND VPWR VPWR _12144_ sky130_fd_sc_hd__mux2_1
X_24649_ _10528_ VGND VGND VPWR VPWR _02410_ sky130_fd_sc_hd__clkbuf_1
X_31748__125 VGND VGND VPWR VPWR _31748__125/HI net125 sky130_fd_sc_hd__conb_1
XFILLER_0_38_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18170_ _05533_ _05534_ VGND VGND VPWR VPWR _05535_ sky130_fd_sc_hd__and2_1
X_15382_ _13412_ _13483_ _13912_ _13913_ _13915_ VGND VGND VPWR VPWR _13916_ sky130_fd_sc_hd__o311a_1
X_27368_ _12102_ VGND VGND VPWR VPWR _03555_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_122_Left_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17121_ _04817_ VGND VGND VPWR VPWR _01478_ sky130_fd_sc_hd__clkbuf_1
X_29107_ _09272_ net3133 _13067_ VGND VGND VPWR VPWR _13069_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_85_Right_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26319_ _11492_ VGND VGND VPWR VPWR _03116_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27299_ _11980_ _12054_ VGND VGND VPWR VPWR _12063_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_131_clk clknet_5_30__leaf_clk VGND VGND VPWR VPWR clknet_leaf_131_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_52_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29038_ _13018_ net1615 _13030_ _13032_ VGND VGND VPWR VPWR _04295_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_150_4084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17052_ net2425 _14466_ _04779_ VGND VGND VPWR VPWR _04781_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_4095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16003_ _14339_ VGND VGND VPWR VPWR _02026_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_204_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31000_ clknet_leaf_100_clk _02735_ VGND VGND VPWR VPWR datamem.data_ram\[22\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_163_4401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_4412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17954_ rvcpu.dp.plem.ALUResultM\[12\] _05268_ VGND VGND VPWR VPWR _05326_ sky130_fd_sc_hd__and2_1
XFILLER_0_206_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_131_Left_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_94_Right_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16905_ _04702_ VGND VGND VPWR VPWR _01587_ sky130_fd_sc_hd__clkbuf_1
X_32951_ clknet_leaf_187_clk _04373_ VGND VGND VPWR VPWR datamem.data_ram\[6\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_1276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17885_ _13178_ _05254_ _05255_ _05256_ _05257_ VGND VGND VPWR VPWR _05258_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_79_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_198_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_198_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_217_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31902_ _04444_ net121 VGND VGND VPWR VPWR datamem.rd_data_mem\[7\] sky130_fd_sc_hd__dlxtn_1
X_19624_ _06919_ VGND VGND VPWR VPWR _06920_ sky130_fd_sc_hd__buf_4
XFILLER_0_206_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16836_ net3147 _14455_ _04659_ VGND VGND VPWR VPWR _04666_ sky130_fd_sc_hd__mux2_1
X_32882_ clknet_leaf_273_clk _04304_ VGND VGND VPWR VPWR datamem.data_ram\[10\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_122_3430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26489__43 clknet_1_1__leaf__10267_ VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__inv_2
XFILLER_0_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_220_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_205_487 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19555_ _06599_ VGND VGND VPWR VPWR _06851_ sky130_fd_sc_hd__buf_8
X_31833_ clknet_leaf_211_clk _03287_ VGND VGND VPWR VPWR datamem.data_ram\[3\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_16767_ _04629_ VGND VGND VPWR VPWR _01660_ sky130_fd_sc_hd__clkbuf_1
X_18506_ _05704_ _05382_ _05784_ VGND VGND VPWR VPWR _05868_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_220_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15718_ _13259_ VGND VGND VPWR VPWR _14183_ sky130_fd_sc_hd__clkbuf_8
X_31764_ clknet_leaf_108_clk _03218_ VGND VGND VPWR VPWR datamem.data_ram\[18\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_840 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19486_ _06781_ VGND VGND VPWR VPWR _06782_ sky130_fd_sc_hd__buf_8
X_16698_ _14162_ net3764 _04587_ VGND VGND VPWR VPWR _04593_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30715_ clknet_leaf_136_clk _02450_ VGND VGND VPWR VPWR datamem.data_ram\[49\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_18437_ _05421_ _05342_ _05349_ _05358_ _05769_ _05689_ VGND VGND VPWR VPWR _05800_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_111_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15649_ _14136_ VGND VGND VPWR VPWR _02185_ sky130_fd_sc_hd__clkbuf_1
X_23658__257 clknet_1_1__leaf__10191_ VGND VGND VPWR VPWR net383 sky130_fd_sc_hd__inv_2
X_31695_ clknet_leaf_50_clk _03153_ VGND VGND VPWR VPWR rvcpu.dp.pcreg.q\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_185_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_140_Left_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18368_ rvcpu.dp.plde.ALUControlE\[0\] rvcpu.dp.plde.ALUControlE\[1\] rvcpu.dp.plde.ALUControlE\[3\]
+ rvcpu.dp.plde.ALUControlE\[2\] VGND VGND VPWR VPWR _05733_ sky130_fd_sc_hd__and4_2
X_30646_ clknet_leaf_190_clk _02381_ VGND VGND VPWR VPWR datamem.data_ram\[51\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17319_ _04922_ VGND VGND VPWR VPWR _01385_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_122_clk clknet_5_27__leaf_clk VGND VGND VPWR VPWR clknet_leaf_122_clk
+ sky130_fd_sc_hd__clkbuf_8
X_18299_ _05663_ VGND VGND VPWR VPWR _05664_ sky130_fd_sc_hd__clkbuf_4
X_30577_ clknet_leaf_179_clk _02312_ VGND VGND VPWR VPWR datamem.data_ram\[54\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_116_3278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20330_ datamem.data_ram\[45\]\[4\] _06921_ _06993_ datamem.data_ram\[47\]\[4\] VGND
+ VGND VPWR VPWR _07622_ sky130_fd_sc_hd__a22o_1
X_32316_ clknet_leaf_232_clk _03738_ VGND VGND VPWR VPWR datamem.data_ram\[31\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_187_4979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20261_ datamem.data_ram\[54\]\[19\] _06683_ _07023_ datamem.data_ram\[50\]\[19\]
+ _07553_ VGND VGND VPWR VPWR _07554_ sky130_fd_sc_hd__o221a_1
X_32247_ clknet_leaf_187_clk _03669_ VGND VGND VPWR VPWR datamem.data_ram\[34\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24144__648 clknet_1_0__leaf__10262_ VGND VGND VPWR VPWR net774 sky130_fd_sc_hd__inv_2
X_22000_ _06591_ VGND VGND VPWR VPWR _09230_ sky130_fd_sc_hd__buf_8
XFILLER_0_228_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3103 rvcpu.dp.rf.reg_file_arr\[19\]\[7\] VGND VGND VPWR VPWR net4253 sky130_fd_sc_hd__dlygate4sd3_1
X_32178_ clknet_leaf_160_clk _03600_ VGND VGND VPWR VPWR datamem.data_ram\[37\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_20192_ datamem.data_ram\[42\]\[11\] _06728_ _06656_ datamem.data_ram\[41\]\[11\]
+ _07484_ VGND VGND VPWR VPWR _07485_ sky130_fd_sc_hd__o221a_1
Xhold3114 datamem.data_ram\[28\]\[28\] VGND VGND VPWR VPWR net4264 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold3125 rvcpu.dp.rf.reg_file_arr\[24\]\[17\] VGND VGND VPWR VPWR net4275 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold3136 datamem.data_ram\[13\]\[12\] VGND VGND VPWR VPWR net4286 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31129_ clknet_leaf_125_clk _02864_ VGND VGND VPWR VPWR datamem.data_ram\[25\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3147 datamem.data_ram\[51\]\[26\] VGND VGND VPWR VPWR net4297 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2402 rvcpu.dp.rf.reg_file_arr\[31\]\[18\] VGND VGND VPWR VPWR net3552 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3158 datamem.data_ram\[55\]\[21\] VGND VGND VPWR VPWR net4308 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2413 datamem.data_ram\[17\]\[27\] VGND VGND VPWR VPWR net3563 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23823__405 clknet_1_0__leaf__10208_ VGND VGND VPWR VPWR net531 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_51_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2424 rvcpu.dp.rf.reg_file_arr\[22\]\[30\] VGND VGND VPWR VPWR net3574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3169 rvcpu.dp.rf.reg_file_arr\[31\]\[25\] VGND VGND VPWR VPWR net4319 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2435 datamem.data_ram\[59\]\[30\] VGND VGND VPWR VPWR net3585 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2446 datamem.data_ram\[40\]\[28\] VGND VGND VPWR VPWR net3596 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1701 rvcpu.dp.rf.reg_file_arr\[7\]\[12\] VGND VGND VPWR VPWR net2851 sky130_fd_sc_hd__dlygate4sd3_1
X_23951_ _10209_ _09229_ _09361_ VGND VGND VPWR VPWR _10229_ sky130_fd_sc_hd__a21oi_4
Xhold1712 datamem.data_ram\[1\]\[24\] VGND VGND VPWR VPWR net2862 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2457 datamem.data_ram\[22\]\[9\] VGND VGND VPWR VPWR net3607 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1723 rvcpu.dp.rf.reg_file_arr\[8\]\[15\] VGND VGND VPWR VPWR net2873 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2468 rvcpu.dp.rf.reg_file_arr\[25\]\[13\] VGND VGND VPWR VPWR net3618 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_189_clk clknet_5_22__leaf_clk VGND VGND VPWR VPWR clknet_leaf_189_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_192_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1734 datamem.data_ram\[46\]\[21\] VGND VGND VPWR VPWR net2884 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_146_3997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2479 rvcpu.dp.rf.reg_file_arr\[15\]\[13\] VGND VGND VPWR VPWR net3629 sky130_fd_sc_hd__dlygate4sd3_1
X_22902_ rvcpu.dp.rf.reg_file_arr\[12\]\[31\] rvcpu.dp.rf.reg_file_arr\[13\]\[31\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[31\] rvcpu.dp.rf.reg_file_arr\[15\]\[31\] _09462_
+ _09465_ VGND VGND VPWR VPWR _10037_ sky130_fd_sc_hd__mux4_1
Xhold1745 datamem.data_ram\[4\]\[26\] VGND VGND VPWR VPWR net2895 sky130_fd_sc_hd__dlygate4sd3_1
X_23903__462 clknet_1_1__leaf__10223_ VGND VGND VPWR VPWR net588 sky130_fd_sc_hd__inv_2
X_26670_ _11683_ net1699 _11675_ _11686_ VGND VGND VPWR VPWR _03273_ sky130_fd_sc_hd__a31o_1
Xhold1756 datamem.data_ram\[59\]\[9\] VGND VGND VPWR VPWR net2906 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1767 datamem.data_ram\[5\]\[26\] VGND VGND VPWR VPWR net2917 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1778 datamem.data_ram\[19\]\[8\] VGND VGND VPWR VPWR net2928 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1789 datamem.data_ram\[47\]\[19\] VGND VGND VPWR VPWR net2939 sky130_fd_sc_hd__dlygate4sd3_1
X_25621_ _10141_ _10051_ VGND VGND VPWR VPWR _11075_ sky130_fd_sc_hd__nand2_8
XFILLER_0_93_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22833_ rvcpu.dp.rf.reg_file_arr\[20\]\[28\] rvcpu.dp.rf.reg_file_arr\[21\]\[28\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[28\] rvcpu.dp.rf.reg_file_arr\[23\]\[28\] _09434_
+ _09558_ VGND VGND VPWR VPWR _09971_ sky130_fd_sc_hd__mux4_1
XFILLER_0_155_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_224_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28340_ _12644_ VGND VGND VPWR VPWR _03985_ sky130_fd_sc_hd__clkbuf_1
X_25552_ _11034_ VGND VGND VPWR VPWR _02807_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_49_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22764_ rvcpu.dp.rf.reg_file_arr\[16\]\[24\] rvcpu.dp.rf.reg_file_arr\[17\]\[24\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[24\] rvcpu.dp.rf.reg_file_arr\[19\]\[24\] _09406_
+ _09408_ VGND VGND VPWR VPWR _09906_ sky130_fd_sc_hd__mux4_1
XFILLER_0_211_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_195_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24503_ _10443_ VGND VGND VPWR VPWR _02349_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28271_ _12363_ net3338 _12603_ VGND VGND VPWR VPWR _12607_ sky130_fd_sc_hd__mux2_1
X_21715_ _08510_ _08959_ VGND VGND VPWR VPWR _08960_ sky130_fd_sc_hd__nor2_1
X_25483_ _10782_ net35 _10996_ net1313 VGND VGND VPWR VPWR _02776_ sky130_fd_sc_hd__a22o_1
X_22695_ rvcpu.dp.rf.reg_file_arr\[0\]\[20\] rvcpu.dp.rf.reg_file_arr\[1\]\[20\] rvcpu.dp.rf.reg_file_arr\[2\]\[20\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[20\] _09714_ _09383_ VGND VGND VPWR VPWR _09841_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_82_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23717__310 clknet_1_0__leaf__10197_ VGND VGND VPWR VPWR net436 sky130_fd_sc_hd__inv_2
X_27222_ _11970_ _12019_ VGND VGND VPWR VPWR _12023_ sky130_fd_sc_hd__and2_1
X_24434_ _10400_ net4438 _10386_ VGND VGND VPWR VPWR _10401_ sky130_fd_sc_hd__mux2_1
X_21646_ rvcpu.dp.rf.reg_file_arr\[8\]\[13\] rvcpu.dp.rf.reg_file_arr\[10\]\[13\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[13\] rvcpu.dp.rf.reg_file_arr\[11\]\[13\] _08693_
+ _08818_ VGND VGND VPWR VPWR _08895_ sky130_fd_sc_hd__mux4_1
XFILLER_0_192_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_882 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27153_ _11980_ _11966_ VGND VGND VPWR VPWR _11981_ sky130_fd_sc_hd__and2_1
XFILLER_0_164_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_113_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_113_clk
+ sky130_fd_sc_hd__clkbuf_8
X_24365_ _10360_ VGND VGND VPWR VPWR _02294_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21577_ _08725_ _08828_ VGND VGND VPWR VPWR _08829_ sky130_fd_sc_hd__nor2_1
XANTENNA_60 _06718_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_71 _06769_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26104_ _11387_ VGND VGND VPWR VPWR _03005_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_82 _06782_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_93 _06810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20528_ _06640_ VGND VGND VPWR VPWR _07819_ sky130_fd_sc_hd__clkbuf_8
X_27084_ rvcpu.ALUResultE\[1\] _06358_ _11598_ VGND VGND VPWR VPWR _11936_ sky130_fd_sc_hd__mux2_1
X_24296_ _10321_ VGND VGND VPWR VPWR _02264_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26035_ _11121_ net1526 _11339_ _11344_ VGND VGND VPWR VPWR _02980_ sky130_fd_sc_hd__a31o_1
X_20459_ datamem.data_ram\[29\]\[20\] _06663_ _07749_ _07750_ VGND VGND VPWR VPWR
+ _07751_ sky130_fd_sc_hd__o211a_1
X_23247_ clknet_1_0__leaf__10108_ VGND VGND VPWR VPWR _10127_ sky130_fd_sc_hd__buf_1
XFILLER_0_123_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22129_ _09236_ net4266 _09332_ VGND VGND VPWR VPWR _09334_ sky130_fd_sc_hd__mux2_1
X_27986_ _12451_ VGND VGND VPWR VPWR _03824_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_201_5316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23763__352 clknet_1_1__leaf__10201_ VGND VGND VPWR VPWR net478 sky130_fd_sc_hd__inv_2
X_29725_ net1071 _01460_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[22\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_201_5327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14951_ _13386_ _13491_ _13497_ _13498_ _13499_ VGND VGND VPWR VPWR _13500_ sky130_fd_sc_hd__a41o_1
X_26937_ _11831_ net1424 _11841_ _11848_ VGND VGND VPWR VPWR _03378_ sky130_fd_sc_hd__a31o_1
XFILLER_0_101_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_197_5220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_197_5231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2980 datamem.data_ram\[5\]\[18\] VGND VGND VPWR VPWR net4130 sky130_fd_sc_hd__dlygate4sd3_1
X_29656_ net1002 _01391_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[24\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_17670_ _05108_ VGND VGND VPWR VPWR _01204_ sky130_fd_sc_hd__clkbuf_1
X_14882_ _13433_ VGND VGND VPWR VPWR _13434_ sky130_fd_sc_hd__clkbuf_4
X_26868_ _11795_ net1540 _11797_ _11804_ VGND VGND VPWR VPWR _03353_ sky130_fd_sc_hd__a31o_1
Xhold2991 rvcpu.dp.rf.reg_file_arr\[29\]\[22\] VGND VGND VPWR VPWR net4141 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_193_5117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_193_5128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16621_ _04552_ VGND VGND VPWR VPWR _01729_ sky130_fd_sc_hd__clkbuf_1
X_28607_ _12799_ VGND VGND VPWR VPWR _04097_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_193_5139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25819_ _08620_ VGND VGND VPWR VPWR _11206_ sky130_fd_sc_hd__clkbuf_2
X_29587_ net941 _01322_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[26\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_26799_ _11753_ net1568 _11761_ _11763_ VGND VGND VPWR VPWR _03325_ sky130_fd_sc_hd__a31o_1
Xmax_cap40 _13058_ VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__buf_4
XFILLER_0_199_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap51 _12270_ VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__buf_4
X_19340_ _06635_ VGND VGND VPWR VPWR _06636_ sky130_fd_sc_hd__buf_6
X_28538_ _12760_ net3315 _12752_ VGND VGND VPWR VPWR _12761_ sky130_fd_sc_hd__mux2_1
X_16552_ _04515_ VGND VGND VPWR VPWR _01769_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap73 _12537_ VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__buf_4
XFILLER_0_43_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap84 _12143_ VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__buf_4
Xmax_cap95 _12650_ VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__buf_4
X_15503_ _13458_ _13360_ _14029_ _13357_ _14030_ VGND VGND VPWR VPWR _14031_ sky130_fd_sc_hd__o221a_1
XFILLER_0_174_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19271_ _06570_ rvcpu.dp.plfd.InstrD\[13\] rvcpu.dp.plfd.InstrD\[12\] rvcpu.dp.plfd.InstrD\[14\]
+ VGND VGND VPWR VPWR _06571_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28469_ _12454_ net3576 _12713_ VGND VGND VPWR VPWR _12717_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16483_ net2693 _14442_ _04478_ VGND VGND VPWR VPWR _04479_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18222_ _05358_ VGND VGND VPWR VPWR _05587_ sky130_fd_sc_hd__inv_2
X_30500_ clknet_leaf_146_clk _02235_ VGND VGND VPWR VPWR datamem.data_ram\[57\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15434_ _13509_ _13565_ VGND VGND VPWR VPWR _13965_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_152_4135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31480_ clknet_leaf_64_clk rvcpu.dp.lAuiPCE\[6\] VGND VGND VPWR VPWR rvcpu.dp.plem.lAuiPCM\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_152_4146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18153_ _05486_ _05494_ _05517_ _05487_ VGND VGND VPWR VPWR _05518_ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30431_ net769 _02166_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[29\]\[10\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_104_clk clknet_5_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_104_clk
+ sky130_fd_sc_hd__clkbuf_8
X_15365_ _13472_ _13589_ _13417_ VGND VGND VPWR VPWR _13900_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_26_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17104_ _04808_ VGND VGND VPWR VPWR _01486_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18084_ _05451_ _05440_ VGND VGND VPWR VPWR _05452_ sky130_fd_sc_hd__and2_1
XFILLER_0_41_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30362_ net708 _02097_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[3\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_15296_ _13547_ _13833_ _13385_ VGND VGND VPWR VPWR _13834_ sky130_fd_sc_hd__and3b_1
XFILLER_0_0_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32101_ clknet_leaf_114_clk _03523_ VGND VGND VPWR VPWR datamem.data_ram\[23\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold308 datamem.data_ram\[6\]\[5\] VGND VGND VPWR VPWR net1458 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold319 datamem.data_ram\[60\]\[3\] VGND VGND VPWR VPWR net1469 sky130_fd_sc_hd__dlygate4sd3_1
X_17035_ net2222 _14449_ _04768_ VGND VGND VPWR VPWR _04772_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30293_ net639 _02028_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[5\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_229_5986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_229_5997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32032_ clknet_leaf_128_clk _03454_ VGND VGND VPWR VPWR datamem.data_ram\[26\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_659 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_221_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_182_4854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_4865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_225_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_209_Left_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18986_ _05302_ _06320_ _05561_ VGND VGND VPWR VPWR _06321_ sky130_fd_sc_hd__or3_1
X_23091__771 clknet_1_1__leaf__10102_ VGND VGND VPWR VPWR net897 sky130_fd_sc_hd__inv_2
Xhold1008 rvcpu.dp.rf.reg_file_arr\[30\]\[18\] VGND VGND VPWR VPWR net2158 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17937_ _05309_ VGND VGND VPWR VPWR rvcpu.dp.SrcBFW_Mux.y\[14\] sky130_fd_sc_hd__dlymetal6s2s_1
X_23013__717 clknet_1_0__leaf__10086_ VGND VGND VPWR VPWR net843 sky130_fd_sc_hd__inv_2
Xhold1019 rvcpu.dp.rf.reg_file_arr\[25\]\[21\] VGND VGND VPWR VPWR net2169 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_175_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32934_ clknet_leaf_134_clk _04356_ VGND VGND VPWR VPWR datamem.data_ram\[7\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_17868_ rvcpu.dp.plde.Rs1E\[0\] VGND VGND VPWR VPWR _05241_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_1_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_85_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_1081 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19607_ datamem.data_ram\[29\]\[8\] _06823_ _06807_ datamem.data_ram\[24\]\[8\] _06902_
+ VGND VGND VPWR VPWR _06903_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_85_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16819_ net2636 _14438_ _04648_ VGND VGND VPWR VPWR _04657_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_141_3872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17799_ rvcpu.dp.plem.ALUResultM\[4\] _05175_ _05191_ _05192_ VGND VGND VPWR VPWR
+ _05193_ sky130_fd_sc_hd__o22a_1
X_32865_ clknet_leaf_254_clk _04287_ VGND VGND VPWR VPWR datamem.data_ram\[11\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_141_3883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31816_ clknet_leaf_104_clk _03270_ VGND VGND VPWR VPWR datamem.data_ram\[9\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19538_ datamem.data_ram\[35\]\[24\] _06829_ _06830_ _06833_ VGND VGND VPWR VPWR
+ _06834_ sky130_fd_sc_hd__o211a_1
XFILLER_0_48_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_81_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32796_ clknet_leaf_233_clk _04218_ VGND VGND VPWR VPWR datamem.data_ram\[13\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_79 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31747_ _04448_ net124 VGND VGND VPWR VPWR rvcpu.ALUControl\[1\] sky130_fd_sc_hd__dlxtn_1
X_19469_ _06684_ VGND VGND VPWR VPWR _06765_ sky130_fd_sc_hd__buf_6
XFILLER_0_174_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_218_Left_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_118_3318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21500_ rvcpu.dp.rf.reg_file_arr\[4\]\[6\] rvcpu.dp.rf.reg_file_arr\[5\]\[6\] rvcpu.dp.rf.reg_file_arr\[6\]\[6\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[6\] _08567_ _08570_ VGND VGND VPWR VPWR _08756_ sky130_fd_sc_hd__mux4_1
XFILLER_0_158_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_118_3329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22480_ _09395_ VGND VGND VPWR VPWR _09637_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_44_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31678_ clknet_leaf_9_clk net1275 VGND VGND VPWR VPWR rvcpu.dp.plmw.ALUResultW\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_44_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23933__488 clknet_1_0__leaf__10227_ VGND VGND VPWR VPWR net614 sky130_fd_sc_hd__inv_2
X_21431_ _08686_ _08688_ _08689_ VGND VGND VPWR VPWR _08690_ sky130_fd_sc_hd__a21o_1
XFILLER_0_90_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30629_ clknet_leaf_217_clk _02364_ VGND VGND VPWR VPWR datamem.data_ram\[51\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21362_ _08623_ VGND VGND VPWR VPWR _08624_ sky130_fd_sc_hd__buf_2
XFILLER_0_140_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23448__98 clknet_1_0__leaf__10156_ VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__inv_2
XFILLER_0_32_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20313_ datamem.data_ram\[10\]\[4\] _07000_ _07133_ datamem.data_ram\[9\]\[4\] VGND
+ VGND VPWR VPWR _07605_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24081_ _10252_ VGND VGND VPWR VPWR _02118_ sky130_fd_sc_hd__clkbuf_1
X_21293_ _08554_ VGND VGND VPWR VPWR _08555_ sky130_fd_sc_hd__buf_4
Xhold820 datamem.data_ram\[50\]\[31\] VGND VGND VPWR VPWR net1970 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_800 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold831 rvcpu.dp.rf.reg_file_arr\[9\]\[19\] VGND VGND VPWR VPWR net1981 sky130_fd_sc_hd__dlygate4sd3_1
Xhold842 rvcpu.dp.rf.reg_file_arr\[17\]\[5\] VGND VGND VPWR VPWR net1992 sky130_fd_sc_hd__dlygate4sd3_1
X_20244_ datamem.data_ram\[59\]\[3\] _06961_ _06948_ datamem.data_ram\[57\]\[3\] VGND
+ VGND VPWR VPWR _07537_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold853 datamem.data_ram\[18\]\[31\] VGND VGND VPWR VPWR net2003 sky130_fd_sc_hd__dlygate4sd3_1
Xhold864 rvcpu.dp.rf.reg_file_arr\[2\]\[19\] VGND VGND VPWR VPWR net2014 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_227_Left_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold875 rvcpu.dp.rf.reg_file_arr\[7\]\[2\] VGND VGND VPWR VPWR net2025 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold886 datamem.data_ram\[53\]\[0\] VGND VGND VPWR VPWR net2036 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27840_ _12366_ VGND VGND VPWR VPWR _03763_ sky130_fd_sc_hd__clkbuf_1
Xhold897 rvcpu.dp.rf.reg_file_arr\[3\]\[2\] VGND VGND VPWR VPWR net2047 sky130_fd_sc_hd__dlygate4sd3_1
X_20175_ datamem.data_ram\[21\]\[11\] _06768_ _06726_ datamem.data_ram\[23\]\[11\]
+ VGND VGND VPWR VPWR _07468_ sky130_fd_sc_hd__o22a_1
XFILLER_0_216_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23215__865 clknet_1_1__leaf__10124_ VGND VGND VPWR VPWR net991 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_38_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2210 datamem.data_ram\[57\]\[13\] VGND VGND VPWR VPWR net3360 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2221 datamem.data_ram\[37\]\[8\] VGND VGND VPWR VPWR net3371 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2232 datamem.data_ram\[31\]\[10\] VGND VGND VPWR VPWR net3382 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2243 datamem.data_ram\[29\]\[28\] VGND VGND VPWR VPWR net3393 sky130_fd_sc_hd__dlygate4sd3_1
X_27771_ _10598_ _12325_ _12260_ VGND VGND VPWR VPWR _12326_ sky130_fd_sc_hd__a21oi_4
X_24983_ _10476_ net2832 net101 VGND VGND VPWR VPWR _10712_ sky130_fd_sc_hd__mux2_1
Xhold2254 datamem.data_ram\[56\]\[11\] VGND VGND VPWR VPWR net3404 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2265 datamem.data_ram\[8\]\[18\] VGND VGND VPWR VPWR net3415 sky130_fd_sc_hd__dlygate4sd3_1
X_29510_ net872 _01245_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[28\]\[17\] sky130_fd_sc_hd__dfxtp_1
Xhold1520 datamem.data_ram\[44\]\[26\] VGND VGND VPWR VPWR net2670 sky130_fd_sc_hd__dlygate4sd3_1
X_26722_ _10756_ net3415 _11714_ VGND VGND VPWR VPWR _11717_ sky130_fd_sc_hd__mux2_1
Xhold1531 rvcpu.dp.rf.reg_file_arr\[18\]\[29\] VGND VGND VPWR VPWR net2681 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2276 datamem.data_ram\[29\]\[9\] VGND VGND VPWR VPWR net3426 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2287 rvcpu.dp.rf.reg_file_arr\[1\]\[23\] VGND VGND VPWR VPWR net3437 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1542 rvcpu.dp.rf.reg_file_arr\[29\]\[1\] VGND VGND VPWR VPWR net2692 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1553 rvcpu.dp.rf.reg_file_arr\[2\]\[8\] VGND VGND VPWR VPWR net2703 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2298 datamem.data_ram\[51\]\[14\] VGND VGND VPWR VPWR net3448 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23526__154 clknet_1_1__leaf__10161_ VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__inv_2
XFILLER_0_58_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1564 rvcpu.dp.rf.reg_file_arr\[2\]\[14\] VGND VGND VPWR VPWR net2714 sky130_fd_sc_hd__dlygate4sd3_1
X_29441_ net803 _01176_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[30\]\[12\] sky130_fd_sc_hd__dfxtp_1
Xhold1575 rvcpu.dp.rf.reg_file_arr\[31\]\[10\] VGND VGND VPWR VPWR net2725 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f__10222_ clknet_0__10222_ VGND VGND VPWR VPWR clknet_1_1__leaf__10222_
+ sky130_fd_sc_hd__clkbuf_16
X_26653_ _07808_ _10932_ _11494_ VGND VGND VPWR VPWR _11674_ sky130_fd_sc_hd__or3_1
Xhold1586 datamem.data_ram\[6\]\[11\] VGND VGND VPWR VPWR net2736 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1597 datamem.data_ram\[20\]\[10\] VGND VGND VPWR VPWR net2747 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25604_ _10570_ _11020_ _10998_ VGND VGND VPWR VPWR _11066_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_169_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__10153_ clknet_0__10153_ VGND VGND VPWR VPWR clknet_1_1__leaf__10153_
+ sky130_fd_sc_hd__clkbuf_16
X_29372_ clknet_leaf_202_clk _01107_ VGND VGND VPWR VPWR datamem.data_ram\[60\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_22816_ rvcpu.dp.rf.reg_file_arr\[28\]\[27\] rvcpu.dp.rf.reg_file_arr\[30\]\[27\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[27\] rvcpu.dp.rf.reg_file_arr\[31\]\[27\] _09446_
+ _09402_ VGND VGND VPWR VPWR _09955_ sky130_fd_sc_hd__mux4_1
X_26584_ _11637_ VGND VGND VPWR VPWR _03236_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28323_ _12635_ VGND VGND VPWR VPWR _03977_ sky130_fd_sc_hd__clkbuf_1
X_25535_ _11025_ VGND VGND VPWR VPWR _02799_ sky130_fd_sc_hd__clkbuf_1
X_22747_ _09390_ _09889_ VGND VGND VPWR VPWR _09890_ sky130_fd_sc_hd__or2_1
Xclkbuf_1_1__f__10084_ clknet_0__10084_ VGND VGND VPWR VPWR clknet_1_1__leaf__10084_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_211_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23793__378 clknet_1_0__leaf__10205_ VGND VGND VPWR VPWR net504 sky130_fd_sc_hd__inv_2
XFILLER_0_109_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28254_ _12456_ net3706 net44 VGND VGND VPWR VPWR _12597_ sky130_fd_sc_hd__mux2_1
X_25466_ _10413_ _10985_ VGND VGND VPWR VPWR _10989_ sky130_fd_sc_hd__and2_1
X_22678_ _09433_ _09824_ _09789_ VGND VGND VPWR VPWR _09825_ sky130_fd_sc_hd__a21o_1
X_27205_ _12005_ net1401 _12007_ _12012_ VGND VGND VPWR VPWR _03482_ sky130_fd_sc_hd__a31o_1
XFILLER_0_180_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24417_ _10389_ VGND VGND VPWR VPWR _02317_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28185_ _12439_ net3357 _12555_ VGND VGND VPWR VPWR _12560_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21629_ _08686_ _08878_ _08689_ VGND VGND VPWR VPWR _08879_ sky130_fd_sc_hd__a21o_1
X_25397_ _10410_ _10950_ VGND VGND VPWR VPWR _10953_ sky130_fd_sc_hd__and2_1
XFILLER_0_152_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15150_ _13291_ _13319_ VGND VGND VPWR VPWR _13694_ sky130_fd_sc_hd__nand2_1
X_27136_ _11956_ net1486 _11964_ _11969_ VGND VGND VPWR VPWR _03456_ sky130_fd_sc_hd__a31o_1
XFILLER_0_35_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24348_ _10351_ VGND VGND VPWR VPWR _02286_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27067_ _11919_ net1727 _11923_ _11926_ VGND VGND VPWR VPWR _03430_ sky130_fd_sc_hd__a31o_1
X_15081_ _13517_ _13625_ _13626_ _13326_ VGND VGND VPWR VPWR _13627_ sky130_fd_sc_hd__o211a_1
X_24279_ _10312_ VGND VGND VPWR VPWR _02256_ sky130_fd_sc_hd__clkbuf_1
X_26018_ net1176 _11329_ _11325_ _11334_ VGND VGND VPWR VPWR _02973_ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18840_ _05700_ _05672_ _05677_ VGND VGND VPWR VPWR _06185_ sky130_fd_sc_hd__mux2_1
X_23687__283 clknet_1_1__leaf__10194_ VGND VGND VPWR VPWR net409 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_224_5861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_224_5872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_224_5883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18771_ _06055_ _06104_ _06105_ _06120_ VGND VGND VPWR VPWR rvcpu.ALUResultE\[14\]
+ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_8_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27969_ _12439_ net3785 _12431_ VGND VGND VPWR VPWR _12440_ sky130_fd_sc_hd__mux2_1
X_15983_ net2030 _13232_ _14322_ VGND VGND VPWR VPWR _14329_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_220_5769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17722_ _13232_ net2098 _05129_ VGND VGND VPWR VPWR _05136_ sky130_fd_sc_hd__mux2_1
X_14934_ _13482_ VGND VGND VPWR VPWR _13483_ sky130_fd_sc_hd__clkbuf_4
X_29708_ net1054 _01443_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[22\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_30980_ clknet_leaf_162_clk _02715_ VGND VGND VPWR VPWR datamem.data_ram\[39\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17653_ _05099_ VGND VGND VPWR VPWR _01212_ sky130_fd_sc_hd__clkbuf_1
X_14865_ _13332_ _13416_ VGND VGND VPWR VPWR _13417_ sky130_fd_sc_hd__or2_1
X_29639_ net985 _01374_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[24\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16604_ _04543_ VGND VGND VPWR VPWR _01737_ sky130_fd_sc_hd__clkbuf_1
X_32650_ clknet_leaf_239_clk _04072_ VGND VGND VPWR VPWR datamem.data_ram\[19\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17584_ _13229_ net2240 _05057_ VGND VGND VPWR VPWR _05063_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14796_ _13346_ _13348_ VGND VGND VPWR VPWR _13349_ sky130_fd_sc_hd__nand2_2
XFILLER_0_202_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_212_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31601_ clknet_leaf_68_clk net1225 VGND VGND VPWR VPWR rvcpu.dp.plmw.PCPlus4W\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19323_ _06618_ VGND VGND VPWR VPWR _06619_ sky130_fd_sc_hd__buf_6
XFILLER_0_97_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_175_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16535_ _04506_ VGND VGND VPWR VPWR _01777_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_670 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32581_ clknet_leaf_233_clk _04003_ VGND VGND VPWR VPWR datamem.data_ram\[21\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_174_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_175_4691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19254_ _06548_ _06556_ VGND VGND VPWR VPWR _06557_ sky130_fd_sc_hd__nand2_1
X_31532_ clknet_leaf_26_clk net1196 VGND VGND VPWR VPWR rvcpu.dp.plem.PCPlus4M\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_16466_ net2085 _14426_ _04467_ VGND VGND VPWR VPWR _04470_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18205_ rvcpu.dp.plde.RD1E\[18\] _05564_ _05489_ VGND VGND VPWR VPWR _05570_ sky130_fd_sc_hd__o21ai_2
X_15417_ _13305_ _13349_ VGND VGND VPWR VPWR _13949_ sky130_fd_sc_hd__and2_1
X_23320__960 clknet_1_0__leaf__10134_ VGND VGND VPWR VPWR net1086 sky130_fd_sc_hd__inv_2
XFILLER_0_72_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19185_ _06495_ _06496_ VGND VGND VPWR VPWR _06497_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_171_4588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31463_ clknet_leaf_75_clk rvcpu.dp.SrcBFW_Mux.y\[21\] VGND VGND VPWR VPWR rvcpu.dp.plem.WriteDataM\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_171_4599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16397_ _14564_ VGND VGND VPWR VPWR _01841_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_3204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18136_ _05500_ _05501_ VGND VGND VPWR VPWR _05502_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_113_3215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30414_ net752 _02149_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[31\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_15348_ _13422_ _13465_ _13622_ _13883_ VGND VGND VPWR VPWR _13884_ sky130_fd_sc_hd__o31a_1
X_31394_ clknet_leaf_38_clk _03097_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCE\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__10242_ clknet_0__10242_ VGND VGND VPWR VPWR clknet_1_0__leaf__10242_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_130_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_184_4905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18067_ _05331_ _05434_ VGND VGND VPWR VPWR _05435_ sky130_fd_sc_hd__and2b_1
Xhold105 rvcpu.dp.plem.ALUResultM\[28\] VGND VGND VPWR VPWR net1255 sky130_fd_sc_hd__dlygate4sd3_1
X_30345_ net691 _02080_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[4\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_15279_ _13328_ _13692_ _13414_ _13366_ VGND VGND VPWR VPWR _13818_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_184_4916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold116 rvcpu.dp.plem.ALUResultM\[12\] VGND VGND VPWR VPWR net1266 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_145_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold127 rvcpu.dp.plde.PCE\[0\] VGND VGND VPWR VPWR net1277 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 rvcpu.dp.plde.PCE\[1\] VGND VGND VPWR VPWR net1288 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__10173_ clknet_0__10173_ VGND VGND VPWR VPWR clknet_1_0__leaf__10173_
+ sky130_fd_sc_hd__clkbuf_16
Xhold149 datamem.data_ram\[42\]\[3\] VGND VGND VPWR VPWR net1299 sky130_fd_sc_hd__dlygate4sd3_1
X_17018_ net3818 _14432_ _04757_ VGND VGND VPWR VPWR _04763_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_74_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30276_ net630 _02011_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[6\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32015_ clknet_leaf_42_clk _03437_ VGND VGND VPWR VPWR rvcpu.dp.pcreg.q\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_226_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_225_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18969_ _06294_ _06305_ VGND VGND VPWR VPWR _06306_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_143_3923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_3934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21980_ rvcpu.dp.plfd.InstrD\[19\] _09202_ _09206_ _09210_ VGND VGND VPWR VPWR _09211_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_217_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_193_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20931_ datamem.data_ram\[35\]\[22\] _07831_ VGND VGND VPWR VPWR _08221_ sky130_fd_sc_hd__or2_1
X_32917_ clknet_leaf_153_clk _04339_ VGND VGND VPWR VPWR datamem.data_ram\[0\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20862_ _08148_ _08149_ _08150_ _08151_ VGND VGND VPWR VPWR _08152_ sky130_fd_sc_hd__a31o_1
XFILLER_0_194_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_191_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32848_ clknet_leaf_85_clk _04270_ VGND VGND VPWR VPWR datamem.data_ram\[7\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_221_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22601_ rvcpu.dp.rf.reg_file_arr\[4\]\[15\] rvcpu.dp.rf.reg_file_arr\[5\]\[15\] rvcpu.dp.rf.reg_file_arr\[6\]\[15\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[15\] _09604_ _09716_ VGND VGND VPWR VPWR _09752_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_102_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20793_ datamem.data_ram\[34\]\[30\] datamem.data_ram\[35\]\[30\] _07849_ VGND VGND
+ VPWR VPWR _08083_ sky130_fd_sc_hd__mux2_1
X_32779_ clknet_leaf_165_clk _04201_ VGND VGND VPWR VPWR datamem.data_ram\[14\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25320_ _10822_ net3714 _10899_ VGND VGND VPWR VPWR _10905_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22532_ _09476_ _09684_ _09686_ _09489_ VGND VGND VPWR VPWR _09687_ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_627 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25251_ _10865_ VGND VGND VPWR VPWR _02675_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22463_ _09615_ _09617_ _09620_ _09412_ _09413_ VGND VGND VPWR VPWR _09621_ sky130_fd_sc_hd__a221o_1
XFILLER_0_151_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24202_ _10271_ VGND VGND VPWR VPWR _02220_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21414_ rvcpu.dp.plfd.InstrD\[17\] VGND VGND VPWR VPWR _08673_ sky130_fd_sc_hd__buf_4
X_25182_ _10500_ VGND VGND VPWR VPWR _10828_ sky130_fd_sc_hd__buf_8
X_22394_ _09389_ _09546_ _09550_ _09555_ VGND VGND VPWR VPWR _09556_ sky130_fd_sc_hd__and4_1
XFILLER_0_17_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23098__777 clknet_1_0__leaf__10103_ VGND VGND VPWR VPWR net903 sky130_fd_sc_hd__inv_2
X_21345_ _06122_ _06130_ rvcpu.ALUResultE\[24\] _08606_ VGND VGND VPWR VPWR _08607_
+ sky130_fd_sc_hd__or4_1
X_29990_ net360 _01725_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[14\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_1194 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28941_ _12976_ VGND VGND VPWR VPWR _04254_ sky130_fd_sc_hd__clkbuf_1
X_21276_ rvcpu.dp.rf.reg_file_arr\[28\]\[0\] rvcpu.dp.rf.reg_file_arr\[30\]\[0\] rvcpu.dp.rf.reg_file_arr\[29\]\[0\]
+ rvcpu.dp.rf.reg_file_arr\[31\]\[0\] _08534_ _08537_ VGND VGND VPWR VPWR _08538_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_103_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold650 datamem.data_ram\[7\]\[5\] VGND VGND VPWR VPWR net1800 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold661 datamem.data_ram\[15\]\[6\] VGND VGND VPWR VPWR net1811 sky130_fd_sc_hd__dlygate4sd3_1
Xhold672 datamem.data_ram\[17\]\[4\] VGND VGND VPWR VPWR net1822 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold683 datamem.data_ram\[18\]\[6\] VGND VGND VPWR VPWR net1833 sky130_fd_sc_hd__dlygate4sd3_1
X_20227_ datamem.data_ram\[13\]\[3\] _06919_ _06925_ datamem.data_ram\[15\]\[3\] _07519_
+ VGND VGND VPWR VPWR _07520_ sky130_fd_sc_hd__a221o_1
Xhold694 rvcpu.dp.plfd.PCPlus4D\[24\] VGND VGND VPWR VPWR net1844 sky130_fd_sc_hd__dlygate4sd3_1
X_28872_ _12702_ net2126 _12932_ VGND VGND VPWR VPWR _12940_ sky130_fd_sc_hd__mux2_1
XFILLER_0_229_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27823_ _12354_ VGND VGND VPWR VPWR _03758_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20158_ datamem.data_ram\[26\]\[27\] _06690_ _06730_ datamem.data_ram\[27\]\[27\]
+ VGND VGND VPWR VPWR _07451_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_5_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2040 datamem.data_ram\[42\]\[8\] VGND VGND VPWR VPWR net3190 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2051 datamem.data_ram\[7\]\[27\] VGND VGND VPWR VPWR net3201 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2062 datamem.data_ram\[22\]\[19\] VGND VGND VPWR VPWR net3212 sky130_fd_sc_hd__dlygate4sd3_1
X_27754_ _12142_ net2492 net48 VGND VGND VPWR VPWR _12317_ sky130_fd_sc_hd__mux2_1
Xhold2073 rvcpu.dp.rf.reg_file_arr\[25\]\[29\] VGND VGND VPWR VPWR net3223 sky130_fd_sc_hd__dlygate4sd3_1
X_20089_ datamem.data_ram\[51\]\[10\] _06829_ _07379_ _07382_ VGND VGND VPWR VPWR
+ _07383_ sky130_fd_sc_hd__o211a_1
X_24966_ _10702_ VGND VGND VPWR VPWR _02553_ sky130_fd_sc_hd__clkbuf_1
Xhold2084 rvcpu.dp.rf.reg_file_arr\[12\]\[23\] VGND VGND VPWR VPWR net3234 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1350 rvcpu.dp.rf.reg_file_arr\[20\]\[25\] VGND VGND VPWR VPWR net2500 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2095 datamem.data_ram\[43\]\[13\] VGND VGND VPWR VPWR net3245 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1361 rvcpu.dp.rf.reg_file_arr\[19\]\[28\] VGND VGND VPWR VPWR net2511 sky130_fd_sc_hd__dlygate4sd3_1
X_26705_ _11707_ VGND VGND VPWR VPWR _03287_ sky130_fd_sc_hd__clkbuf_1
Xhold1372 datamem.data_ram\[44\]\[21\] VGND VGND VPWR VPWR net2522 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27685_ _12279_ _10908_ _12260_ VGND VGND VPWR VPWR _12280_ sky130_fd_sc_hd__a21oi_4
X_24897_ _10665_ VGND VGND VPWR VPWR _02521_ sky130_fd_sc_hd__clkbuf_1
Xhold1383 rvcpu.dp.rf.reg_file_arr\[8\]\[25\] VGND VGND VPWR VPWR net2533 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1394 datamem.data_ram\[48\]\[23\] VGND VGND VPWR VPWR net2544 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_501 _11603_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29424_ clknet_leaf_98_clk _01159_ VGND VGND VPWR VPWR datamem.data_ram\[5\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_512 _13222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26636_ _11618_ net1717 _11662_ _11664_ VGND VGND VPWR VPWR _03261_ sky130_fd_sc_hd__a31o_1
XFILLER_0_197_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14650_ rvcpu.dp.plmw.ALUResultW\[18\] rvcpu.dp.plmw.ReadDataW\[18\] rvcpu.dp.plmw.PCPlus4W\[18\]
+ rvcpu.dp.plmw.lAuiPCW\[18\] _13192_ _13193_ VGND VGND VPWR VPWR _13222_ sky130_fd_sc_hd__mux4_2
XANTENNA_523 _13257_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_1_1__f__10205_ clknet_0__10205_ VGND VGND VPWR VPWR clknet_1_1__leaf__10205_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_19_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_574 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_534 rvcpu.dp.plmw.ReadDataW\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23801__385 clknet_1_1__leaf__10206_ VGND VGND VPWR VPWR net511 sky130_fd_sc_hd__inv_2
XFILLER_0_196_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_545 _06753_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_556 _07845_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_567 rvcpu.dp.plmw.ReadDataW\[24\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29355_ clknet_leaf_141_clk _01090_ VGND VGND VPWR VPWR datamem.data_ram\[61\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__10136_ clknet_0__10136_ VGND VGND VPWR VPWR clknet_1_1__leaf__10136_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_67_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26567_ _11628_ VGND VGND VPWR VPWR _03228_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_200_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28306_ _12626_ VGND VGND VPWR VPWR _03969_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16320_ net2558 _14486_ _14488_ VGND VGND VPWR VPWR _14523_ sky130_fd_sc_hd__mux2_1
X_25518_ _10991_ net1550 _11009_ _11015_ VGND VGND VPWR VPWR _02792_ sky130_fd_sc_hd__a31o_1
XFILLER_0_138_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29286_ _13164_ VGND VGND VPWR VPWR _04411_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_211_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_188_5005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_188_5016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28237_ _12439_ net2843 _12583_ VGND VGND VPWR VPWR _12588_ sky130_fd_sc_hd__mux2_1
X_16251_ _13277_ VGND VGND VPWR VPWR _14486_ sky130_fd_sc_hd__buf_4
X_25449_ _10048_ _10981_ _10982_ net1337 VGND VGND VPWR VPWR _02756_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23042__743 clknet_1_0__leaf__10089_ VGND VGND VPWR VPWR net869 sky130_fd_sc_hd__inv_2
XFILLER_0_36_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15202_ _13526_ _13541_ VGND VGND VPWR VPWR _13744_ sky130_fd_sc_hd__nand2_1
XFILLER_0_180_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28168_ _12365_ net3249 _12546_ VGND VGND VPWR VPWR _12551_ sky130_fd_sc_hd__mux2_1
X_16182_ _14439_ VGND VGND VPWR VPWR _01939_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_535 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15133_ _13607_ _13553_ VGND VGND VPWR VPWR _13678_ sky130_fd_sc_hd__nor2_1
X_27119_ _11956_ net1816 _11952_ _11958_ VGND VGND VPWR VPWR _03450_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_226_5912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23157__830 clknet_1_1__leaf__10109_ VGND VGND VPWR VPWR net956 sky130_fd_sc_hd__inv_2
X_28099_ _12514_ VGND VGND VPWR VPWR _03874_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_226_5923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23427__79 clknet_1_0__leaf__10154_ VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_147_4012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30130_ net492 _01865_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[10\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_15064_ _13364_ _13610_ _13410_ VGND VGND VPWR VPWR _13611_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_147_4023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19941_ datamem.data_ram\[45\]\[18\] _06664_ _06783_ datamem.data_ram\[41\]\[18\]
+ VGND VGND VPWR VPWR _07235_ sky130_fd_sc_hd__o22a_1
XFILLER_0_107_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_147_4034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30061_ net423 _01796_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[12\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_19872_ datamem.data_ram\[26\]\[1\] _06989_ _06973_ datamem.data_ram\[24\]\[1\] VGND
+ VGND VPWR VPWR _07167_ sky130_fd_sc_hd__a22o_1
X_18823_ _05497_ _06168_ VGND VGND VPWR VPWR _06169_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18754_ _05611_ _06091_ _05311_ VGND VGND VPWR VPWR _06104_ sky130_fd_sc_hd__a21o_1
X_15966_ net1922 _13207_ _14311_ VGND VGND VPWR VPWR _14320_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_106_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_106_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_216_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14917_ _13466_ _13423_ VGND VGND VPWR VPWR _13467_ sky130_fd_sc_hd__nor2_1
X_17705_ _13207_ net1976 _05118_ VGND VGND VPWR VPWR _05127_ sky130_fd_sc_hd__mux2_1
X_30963_ clknet_leaf_157_clk _02698_ VGND VGND VPWR VPWR datamem.data_ram\[3\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_18685_ _05599_ _05601_ _05605_ VGND VGND VPWR VPWR _06039_ sky130_fd_sc_hd__a21boi_1
X_15897_ _14283_ VGND VGND VPWR VPWR _02076_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_159_Right_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_188_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_177_4742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32702_ clknet_leaf_244_clk _04124_ VGND VGND VPWR VPWR datamem.data_ram\[17\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_14848_ _13400_ VGND VGND VPWR VPWR _13401_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_177_4753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17636_ _05090_ VGND VGND VPWR VPWR _01220_ sky130_fd_sc_hd__clkbuf_1
X_30894_ clknet_leaf_137_clk _02629_ VGND VGND VPWR VPWR datamem.data_ram\[41\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_67_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32633_ clknet_leaf_255_clk _04055_ VGND VGND VPWR VPWR datamem.data_ram\[1\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_17567_ _13204_ net2440 _05046_ VGND VGND VPWR VPWR _05054_ sky130_fd_sc_hd__mux2_1
X_14779_ _13331_ VGND VGND VPWR VPWR _13332_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_173_4639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19306_ _06601_ VGND VGND VPWR VPWR _06602_ sky130_fd_sc_hd__clkbuf_8
X_16518_ net2963 _14478_ _04489_ VGND VGND VPWR VPWR _04497_ sky130_fd_sc_hd__mux2_1
X_32564_ clknet_leaf_80_clk _03986_ VGND VGND VPWR VPWR datamem.data_ram\[22\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17498_ _05017_ VGND VGND VPWR VPWR _01293_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31515_ clknet_leaf_52_clk net1186 VGND VGND VPWR VPWR rvcpu.dp.plem.PCPlus4M\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19237_ _06540_ _06541_ VGND VGND VPWR VPWR _06542_ sky130_fd_sc_hd__nor2_1
XFILLER_0_143_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23475__123 clknet_1_1__leaf__10158_ VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__inv_2
X_16449_ _04459_ VGND VGND VPWR VPWR _01816_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_171_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32495_ clknet_leaf_74_clk _03917_ VGND VGND VPWR VPWR datamem.data_ram\[25\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_136_3760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_3771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19168_ _06480_ _06481_ VGND VGND VPWR VPWR _06482_ sky130_fd_sc_hd__or2b_1
X_31446_ clknet_leaf_76_clk rvcpu.dp.SrcBFW_Mux.y\[4\] VGND VGND VPWR VPWR rvcpu.dp.plem.WriteDataM\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_76_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_3657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18119_ _05484_ _05485_ VGND VGND VPWR VPWR _05486_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_132_3668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19099_ rvcpu.dp.plde.ImmExtE\[11\] rvcpu.dp.plde.PCE\[11\] VGND VGND VPWR VPWR _06421_
+ sky130_fd_sc_hd__or2_1
X_31377_ clknet_leaf_22_clk _03080_ VGND VGND VPWR VPWR rvcpu.dp.plde.ImmExtE\[26\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_170_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__10225_ clknet_0__10225_ VGND VGND VPWR VPWR clknet_1_0__leaf__10225_
+ sky130_fd_sc_hd__clkbuf_16
X_21130_ _07820_ _08416_ _08418_ _07867_ VGND VGND VPWR VPWR _08419_ sky130_fd_sc_hd__o211a_1
X_30328_ net674 _02063_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[4\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__10156_ clknet_0__10156_ VGND VGND VPWR VPWR clknet_1_0__leaf__10156_
+ sky130_fd_sc_hd__clkbuf_16
X_23019__723 clknet_1_1__leaf__10086_ VGND VGND VPWR VPWR net849 sky130_fd_sc_hd__inv_2
XFILLER_0_1_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21061_ _07859_ _08348_ _08349_ _07866_ VGND VGND VPWR VPWR _08350_ sky130_fd_sc_hd__o22a_1
X_30259_ net613 _01994_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[6\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_35_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20012_ datamem.data_ram\[54\]\[2\] _06950_ _06930_ datamem.data_ram\[50\]\[2\] VGND
+ VGND VPWR VPWR _07306_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_35_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__10087_ clknet_0__10087_ VGND VGND VPWR VPWR clknet_1_0__leaf__10087_
+ sky130_fd_sc_hd__clkbuf_16
X_24820_ _10390_ net3419 _10621_ VGND VGND VPWR VPWR _10624_ sky130_fd_sc_hd__mux2_1
XFILLER_0_213_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24751_ _10394_ net2935 _10580_ VGND VGND VPWR VPWR _10585_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21963_ _09194_ VGND VGND VPWR VPWR _01058_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_193_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_93_clk clknet_5_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_93_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_154_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_126_Right_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20914_ datamem.data_ram\[30\]\[22\] datamem.data_ram\[31\]\[22\] _07836_ VGND VGND
+ VPWR VPWR _08204_ sky130_fd_sc_hd__mux2_1
X_27470_ _12164_ VGND VGND VPWR VPWR _03595_ sky130_fd_sc_hd__clkbuf_1
X_23327__966 clknet_1_1__leaf__10135_ VGND VGND VPWR VPWR net1092 sky130_fd_sc_hd__inv_2
X_24682_ _10394_ net3840 _10543_ VGND VGND VPWR VPWR _10548_ sky130_fd_sc_hd__mux2_1
XFILLER_0_178_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21894_ _08522_ _09128_ VGND VGND VPWR VPWR _09129_ sky130_fd_sc_hd__or2_1
X_26421_ _11545_ rvcpu.ALUResultE\[13\] VGND VGND VPWR VPWR _11558_ sky130_fd_sc_hd__and2_1
XFILLER_0_178_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_169_Left_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23633_ _09267_ net3178 _10182_ VGND VGND VPWR VPWR _10183_ sky130_fd_sc_hd__mux2_1
XFILLER_0_221_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_193_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23939__494 clknet_1_1__leaf__10227_ VGND VGND VPWR VPWR net620 sky130_fd_sc_hd__inv_2
X_20845_ _07867_ _08134_ VGND VGND VPWR VPWR _08135_ sky130_fd_sc_hd__or2_1
XFILLER_0_194_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29140_ _13086_ VGND VGND VPWR VPWR _04343_ sky130_fd_sc_hd__clkbuf_1
X_26352_ _10783_ _11507_ _11508_ net1331 VGND VGND VPWR VPWR _03133_ sky130_fd_sc_hd__a22o_1
X_20776_ _06681_ _07872_ VGND VGND VPWR VPWR _08066_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25303_ _10894_ VGND VGND VPWR VPWR _02698_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29071_ _12751_ net3593 _13049_ VGND VGND VPWR VPWR _13050_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22515_ _09662_ _09666_ _09670_ _09491_ VGND VGND VPWR VPWR _01134_ sky130_fd_sc_hd__o31a_1
X_26283_ net1821 _11467_ VGND VGND VPWR VPWR _11474_ sky130_fd_sc_hd__and2_1
XFILLER_0_119_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28022_ _09350_ _12335_ _12356_ VGND VGND VPWR VPWR _12473_ sky130_fd_sc_hd__a21oi_4
X_25234_ _10856_ VGND VGND VPWR VPWR _02667_ sky130_fd_sc_hd__clkbuf_1
X_22446_ rvcpu.dp.rf.reg_file_arr\[4\]\[7\] rvcpu.dp.rf.reg_file_arr\[5\]\[7\] rvcpu.dp.rf.reg_file_arr\[6\]\[7\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[7\] _09604_ _09424_ VGND VGND VPWR VPWR _09605_ sky130_fd_sc_hd__mux4_1
XFILLER_0_161_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25165_ _10816_ net3669 net58 VGND VGND VPWR VPWR _10817_ sky130_fd_sc_hd__mux2_1
X_22377_ rvcpu.dp.rf.reg_file_arr\[24\]\[4\] rvcpu.dp.rf.reg_file_arr\[25\]\[4\] rvcpu.dp.rf.reg_file_arr\[26\]\[4\]
+ rvcpu.dp.rf.reg_file_arr\[27\]\[4\] _09393_ _09395_ VGND VGND VPWR VPWR _09539_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_206_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21328_ rvcpu.dp.plfd.InstrD\[22\] rvcpu.dp.plde.RdE\[2\] VGND VGND VPWR VPWR _08590_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_60_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25096_ _10048_ _10779_ _10781_ net1323 VGND VGND VPWR VPWR _02604_ sky130_fd_sc_hd__a22o_1
X_29973_ net343 _01708_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[14\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21259_ _08515_ _08520_ VGND VGND VPWR VPWR _08521_ sky130_fd_sc_hd__nor2_1
X_28924_ _12967_ VGND VGND VPWR VPWR _04246_ sky130_fd_sc_hd__clkbuf_1
Xhold480 datamem.data_ram\[33\]\[2\] VGND VGND VPWR VPWR net1630 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold491 datamem.data_ram\[22\]\[1\] VGND VGND VPWR VPWR net1641 sky130_fd_sc_hd__dlygate4sd3_1
X_28855_ _12749_ net2267 _12923_ VGND VGND VPWR VPWR _12931_ sky130_fd_sc_hd__mux2_1
X_15820_ _14241_ VGND VGND VPWR VPWR _02111_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_176_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27806_ _08125_ _09268_ VGND VGND VPWR VPWR _12345_ sky130_fd_sc_hd__nor2_2
XFILLER_0_99_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_205_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28786_ _12894_ VGND VGND VPWR VPWR _04181_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_216_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25998_ rvcpu.dp.plfd.InstrD\[19\] _11315_ _11312_ _11323_ VGND VGND VPWR VPWR _02964_
+ sky130_fd_sc_hd__o211a_1
X_27737_ _12125_ net2423 _12307_ VGND VGND VPWR VPWR _12308_ sky130_fd_sc_hd__mux2_1
X_15751_ _14204_ VGND VGND VPWR VPWR _02151_ sky130_fd_sc_hd__clkbuf_1
X_24949_ _10693_ VGND VGND VPWR VPWR _02545_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_220_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_84_clk clknet_5_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_84_clk sky130_fd_sc_hd__clkbuf_8
Xhold1180 datamem.data_ram\[0\]\[24\] VGND VGND VPWR VPWR net2330 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14702_ _13261_ VGND VGND VPWR VPWR _03178_ sky130_fd_sc_hd__clkbuf_1
Xhold1191 datamem.data_ram\[62\]\[27\] VGND VGND VPWR VPWR net2341 sky130_fd_sc_hd__dlygate4sd3_1
X_18470_ _05831_ _05832_ _05674_ VGND VGND VPWR VPWR _05833_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23799__384 clknet_1_1__leaf__10205_ VGND VGND VPWR VPWR net510 sky130_fd_sc_hd__inv_2
X_27668_ _12080_ net2741 net51 VGND VGND VPWR VPWR _12271_ sky130_fd_sc_hd__mux2_1
X_15682_ _14158_ net2673 _14152_ VGND VGND VPWR VPWR _14159_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_320 _14428_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_219_5760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_331 _14457_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17421_ _14135_ net2574 _04974_ VGND VGND VPWR VPWR _04977_ sky130_fd_sc_hd__mux2_1
XANTENNA_342 _14468_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_212_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14633_ rvcpu.dp.plmw.ALUResultW\[22\] rvcpu.dp.plmw.ReadDataW\[22\] rvcpu.dp.plmw.PCPlus4W\[22\]
+ rvcpu.dp.plmw.lAuiPCW\[22\] _13169_ _13171_ VGND VGND VPWR VPWR _13209_ sky130_fd_sc_hd__mux4_2
X_29407_ clknet_leaf_0_clk _01142_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD2E\[18\] sky130_fd_sc_hd__dfxtp_1
X_26619_ _11657_ VGND VGND VPWR VPWR _03251_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_200_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_353 rvcpu.ALUResultE\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_364 rvcpu.dp.SrcBFW_Mux.y\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27599_ _12142_ net4061 net81 VGND VGND VPWR VPWR _12234_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_215_5646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_375 rvcpu.dp.plem.ALUResultM\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_386 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_0__10219_ _10219_ VGND VGND VPWR VPWR clknet_0__10219_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_56_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_215_5657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_397 _06096_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17352_ _04940_ VGND VGND VPWR VPWR _01362_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29338_ clknet_leaf_269_clk _01073_ VGND VGND VPWR VPWR datamem.data_ram\[62\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16303_ _14514_ VGND VGND VPWR VPWR _01885_ sky130_fd_sc_hd__clkbuf_1
X_17283_ net2783 _13183_ _04902_ VGND VGND VPWR VPWR _04904_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29269_ _13155_ VGND VGND VPWR VPWR _04403_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_183_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31300_ clknet_leaf_48_clk _03003_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCPlus4E\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_19022_ rvcpu.dp.plde.luiE VGND VGND VPWR VPWR _06355_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16234_ net1971 _14474_ _14464_ VGND VGND VPWR VPWR _14475_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32280_ clknet_leaf_168_clk _03702_ VGND VGND VPWR VPWR datamem.data_ram\[33\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_805 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload306 clknet_1_1__leaf__10197_ VGND VGND VPWR VPWR clkload306/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_67_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_183_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload14 clknet_5_16__leaf_clk VGND VGND VPWR VPWR clkload14/X sky130_fd_sc_hd__clkbuf_8
Xclkload317 clknet_1_1__leaf__10152_ VGND VGND VPWR VPWR clkload317/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_152_164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31231_ clknet_leaf_42_clk _02934_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCD\[20\] sky130_fd_sc_hd__dfxtp_1
Xclkload25 clknet_5_30__leaf_clk VGND VGND VPWR VPWR clkload25/Y sky130_fd_sc_hd__inv_6
XFILLER_0_141_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload328 clknet_1_0__leaf__10266_ VGND VGND VPWR VPWR clkload328/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload36 clknet_leaf_24_clk VGND VGND VPWR VPWR clkload36/Y sky130_fd_sc_hd__clkinv_1
Xclkload339 clknet_1_1__leaf__10129_ VGND VGND VPWR VPWR clkload339/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_51_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16165_ _13189_ VGND VGND VPWR VPWR _14428_ sky130_fd_sc_hd__clkbuf_4
Xclkload47 clknet_leaf_29_clk VGND VGND VPWR VPWR clkload47/Y sky130_fd_sc_hd__clkinv_1
XFILLER_0_24_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload58 clknet_leaf_4_clk VGND VGND VPWR VPWR clkload58/Y sky130_fd_sc_hd__inv_6
XFILLER_0_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload69 clknet_leaf_67_clk VGND VGND VPWR VPWR clkload69/Y sky130_fd_sc_hd__clkinvlp_2
X_15116_ _13307_ _13393_ _13598_ _13429_ _13660_ VGND VGND VPWR VPWR _13661_ sky130_fd_sc_hd__a41o_1
XFILLER_0_224_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31162_ clknet_leaf_69_clk rvcpu.ALUResultE\[21\] VGND VGND VPWR VPWR rvcpu.dp.plem.ALUResultM\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_71_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16096_ net4416 _13195_ _14385_ VGND VGND VPWR VPWR _14390_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30113_ net475 _01848_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[10\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_15047_ _13353_ _13593_ _13438_ VGND VGND VPWR VPWR _13594_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_166_4476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19924_ datamem.data_ram\[54\]\[17\] _06683_ _06664_ datamem.data_ram\[53\]\[17\]
+ VGND VGND VPWR VPWR _07219_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_228_Right_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31093_ clknet_leaf_254_clk _02828_ VGND VGND VPWR VPWR datamem.data_ram\[9\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_166_4487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2809 datamem.data_ram\[40\]\[24\] VGND VGND VPWR VPWR net3959 sky130_fd_sc_hd__dlygate4sd3_1
X_30044_ net406 _01779_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[13\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_19855_ datamem.data_ram\[60\]\[1\] _06977_ _07148_ _07149_ VGND VGND VPWR VPWR _07150_
+ sky130_fd_sc_hd__a211o_1
X_18806_ _05504_ _05567_ _06134_ _05655_ VGND VGND VPWR VPWR _06153_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_207_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19786_ _06602_ VGND VGND VPWR VPWR _07081_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_30_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16998_ _04751_ VGND VGND VPWR VPWR _01543_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_69_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18737_ _06085_ _06086_ _05886_ VGND VGND VPWR VPWR _06088_ sky130_fd_sc_hd__a21oi_1
X_15949_ _14310_ VGND VGND VPWR VPWR _14311_ sky130_fd_sc_hd__clkbuf_4
X_31995_ clknet_leaf_128_clk _03417_ VGND VGND VPWR VPWR datamem.data_ram\[31\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_75_clk clknet_5_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_75_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_125_3494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30946_ clknet_leaf_96_clk _02681_ VGND VGND VPWR VPWR datamem.data_ram\[3\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_18668_ _05775_ _05833_ VGND VGND VPWR VPWR _06023_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23049__749 clknet_1_1__leaf__10090_ VGND VGND VPWR VPWR net875 sky130_fd_sc_hd__inv_2
XFILLER_0_114_1111 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17619_ _14234_ _14347_ VGND VGND VPWR VPWR _05081_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_138_3800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18599_ _05354_ _05355_ VGND VGND VPWR VPWR _05957_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_138_3811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30877_ clknet_leaf_264_clk _02612_ VGND VGND VPWR VPWR datamem.data_ram\[42\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32616_ clknet_leaf_171_clk _04038_ VGND VGND VPWR VPWR datamem.data_ram\[20\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_20630_ datamem.data_ram\[5\]\[29\] _06663_ _06784_ datamem.data_ram\[7\]\[29\] VGND
+ VGND VPWR VPWR _07921_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_28_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24071__597 clknet_1_1__leaf__10248_ VGND VGND VPWR VPWR net723 sky130_fd_sc_hd__inv_2
XFILLER_0_191_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_134_3708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20561_ datamem.data_ram\[13\]\[21\] _06664_ _07850_ _07851_ VGND VGND VPWR VPWR
+ _07852_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_134_3719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32547_ clknet_leaf_248_clk _03969_ VGND VGND VPWR VPWR datamem.data_ram\[23\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload8 clknet_5_9__leaf_clk VGND VGND VPWR VPWR clkload8/Y sky130_fd_sc_hd__inv_12
XFILLER_0_144_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22300_ _09381_ VGND VGND VPWR VPWR _09465_ sky130_fd_sc_hd__buf_4
XFILLER_0_171_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20492_ _06589_ _07646_ _07783_ _06583_ VGND VGND VPWR VPWR _07784_ sky130_fd_sc_hd__a211o_1
XFILLER_0_15_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23280_ clknet_1_0__leaf__10079_ VGND VGND VPWR VPWR _10130_ sky130_fd_sc_hd__buf_1
X_32478_ clknet_leaf_249_clk _03900_ VGND VGND VPWR VPWR datamem.data_ram\[26\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_225_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22231_ _09391_ _09396_ VGND VGND VPWR VPWR _09397_ sky130_fd_sc_hd__or2_1
X_31429_ clknet_leaf_97_clk _03132_ VGND VGND VPWR VPWR datamem.data_ram\[44\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22162_ _09351_ _09301_ _09231_ VGND VGND VPWR VPWR _09352_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_160_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__10208_ clknet_0__10208_ VGND VGND VPWR VPWR clknet_1_0__leaf__10208_
+ sky130_fd_sc_hd__clkbuf_16
X_21113_ datamem.data_ram\[28\]\[7\] _06652_ _08401_ _06615_ VGND VGND VPWR VPWR _08402_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_112_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_58_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26970_ _11827_ _11866_ VGND VGND VPWR VPWR _11869_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22093_ _09305_ VGND VGND VPWR VPWR _09306_ sky130_fd_sc_hd__buf_2
XFILLER_0_100_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__10139_ clknet_0__10139_ VGND VGND VPWR VPWR clknet_1_0__leaf__10139_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_100_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25921_ net1362 _11275_ _11273_ _11280_ VGND VGND VPWR VPWR _02930_ sky130_fd_sc_hd__o211a_1
X_21044_ datamem.data_ram\[0\]\[31\] datamem.data_ram\[1\]\[31\] _06933_ VGND VGND
+ VPWR VPWR _08333_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_227_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28640_ _12739_ net2840 net71 VGND VGND VPWR VPWR _12817_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_54_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25852_ _11233_ VGND VGND VPWR VPWR _02908_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_199_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24803_ _10444_ net4035 _10612_ VGND VGND VPWR VPWR _10615_ sky130_fd_sc_hd__mux2_1
XFILLER_0_199_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28571_ _12756_ net3039 _12777_ VGND VGND VPWR VPWR _12780_ sky130_fd_sc_hd__mux2_1
X_25783_ rvcpu.dp.pcreg.q\[11\] _11171_ rvcpu.dp.pcreg.q\[12\] VGND VGND VPWR VPWR
+ _11179_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_158_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_66_clk clknet_5_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_66_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_213_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_177_Left_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27522_ _12089_ net2978 net99 VGND VGND VPWR VPWR _12193_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24734_ _10448_ net3151 _10571_ VGND VGND VPWR VPWR _10576_ sky130_fd_sc_hd__mux2_1
X_21946_ rvcpu.dp.rf.reg_file_arr\[16\]\[30\] rvcpu.dp.rf.reg_file_arr\[17\]\[30\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[30\] rvcpu.dp.rf.reg_file_arr\[19\]\[30\] _08516_
+ _08518_ VGND VGND VPWR VPWR _09178_ sky130_fd_sc_hd__mux4_1
XFILLER_0_16_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27453_ _12154_ VGND VGND VPWR VPWR _03588_ sky130_fd_sc_hd__clkbuf_1
X_24665_ _10055_ VGND VGND VPWR VPWR _10538_ sky130_fd_sc_hd__buf_2
XFILLER_0_179_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23260__906 clknet_1_0__leaf__10128_ VGND VGND VPWR VPWR net1032 sky130_fd_sc_hd__inv_2
X_21877_ _08725_ _09112_ VGND VGND VPWR VPWR _09113_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26404_ _11545_ rvcpu.ALUResultE\[8\] VGND VGND VPWR VPWR _11546_ sky130_fd_sc_hd__and2_1
X_23616_ clknet_1_1__leaf__10172_ VGND VGND VPWR VPWR _10180_ sky130_fd_sc_hd__buf_1
X_23872__434 clknet_1_0__leaf__10220_ VGND VGND VPWR VPWR net560 sky130_fd_sc_hd__inv_2
XFILLER_0_166_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27384_ _12111_ VGND VGND VPWR VPWR _03562_ sky130_fd_sc_hd__clkbuf_1
X_20828_ datamem.data_ram\[15\]\[30\] _06706_ _06595_ _08117_ VGND VGND VPWR VPWR
+ _08118_ sky130_fd_sc_hd__o211a_1
X_24596_ _10400_ net2601 _10491_ VGND VGND VPWR VPWR _10499_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29123_ _13077_ VGND VGND VPWR VPWR _04335_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26335_ _11047_ _11497_ VGND VGND VPWR VPWR _11503_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20759_ datamem.data_ram\[3\]\[6\] _07832_ VGND VGND VPWR VPWR _08049_ sky130_fd_sc_hd__or2_1
XFILLER_0_53_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_210_5532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_210_5543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29054_ _09266_ net3425 net65 VGND VGND VPWR VPWR _13041_ sky130_fd_sc_hd__mux2_1
X_26266_ net1884 _11432_ VGND VGND VPWR VPWR _11465_ sky130_fd_sc_hd__and2_1
XFILLER_0_208_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28005_ _10542_ _12325_ _12356_ VGND VGND VPWR VPWR _12464_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_186_Left_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25217_ _10847_ VGND VGND VPWR VPWR _02659_ sky130_fd_sc_hd__clkbuf_1
X_22429_ _09415_ _09586_ _09588_ VGND VGND VPWR VPWR _09589_ sky130_fd_sc_hd__a21o_1
XFILLER_0_208_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26197_ _11413_ VGND VGND VPWR VPWR _11436_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_122_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25148_ _10806_ VGND VGND VPWR VPWR _02631_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17970_ rvcpu.dp.plem.ALUResultM\[7\] _05339_ _05340_ _13256_ VGND VGND VPWR VPWR
+ _05341_ sky130_fd_sc_hd__o22a_1
XFILLER_0_130_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29956_ net326 _01691_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[15\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_25079_ _10729_ net3923 net89 VGND VGND VPWR VPWR _10771_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_208_5483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_208_5494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16921_ net2092 _14472_ _04706_ VGND VGND VPWR VPWR _04711_ sky130_fd_sc_hd__mux2_1
X_28907_ _12958_ VGND VGND VPWR VPWR _04238_ sky130_fd_sc_hd__clkbuf_1
X_29887_ net265 _01622_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[17\]\[18\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_161_4351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19640_ _06935_ VGND VGND VPWR VPWR _06936_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_161_4362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28838_ _12766_ net2038 _12914_ VGND VGND VPWR VPWR _12922_ sky130_fd_sc_hd__mux2_1
X_16852_ _04674_ VGND VGND VPWR VPWR _01612_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_205_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23807__391 clknet_1_0__leaf__10206_ VGND VGND VPWR VPWR net517 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_195_Left_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15803_ _14231_ VGND VGND VPWR VPWR _02126_ sky130_fd_sc_hd__clkbuf_1
X_16783_ net2304 _14470_ _04634_ VGND VGND VPWR VPWR _04638_ sky130_fd_sc_hd__mux2_1
X_19571_ datamem.data_ram\[6\]\[8\] _06718_ _06789_ datamem.data_ram\[1\]\[8\] VGND
+ VGND VPWR VPWR _06867_ sky130_fd_sc_hd__o22a_1
XFILLER_0_189_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28769_ _12702_ net2678 _12877_ VGND VGND VPWR VPWR _12885_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_57_clk clknet_5_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_57_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_172_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_217_5708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18522_ _05375_ _05702_ _05878_ _05882_ VGND VGND VPWR VPWR _05883_ sky130_fd_sc_hd__a31o_1
X_26504__56 clknet_1_1__leaf__11602_ VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__inv_2
X_30800_ clknet_leaf_224_clk _02535_ VGND VGND VPWR VPWR datamem.data_ram\[45\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15734_ _14193_ net2692 _14130_ VGND VGND VPWR VPWR _14194_ sky130_fd_sc_hd__mux2_1
X_31780_ clknet_leaf_180_clk _03234_ VGND VGND VPWR VPWR datamem.data_ram\[6\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18453_ _05577_ _05809_ _05811_ _05815_ VGND VGND VPWR VPWR _05816_ sky130_fd_sc_hd__a31o_1
X_30731_ clknet_leaf_195_clk _02466_ VGND VGND VPWR VPWR datamem.data_ram\[48\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_15665_ _13206_ VGND VGND VPWR VPWR _14147_ sky130_fd_sc_hd__clkbuf_8
XANTENNA_150 _07874_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_120_3380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_161 _08568_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_213_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17404_ _04967_ VGND VGND VPWR VPWR _01337_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14616_ _13196_ VGND VGND VPWR VPWR _03199_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_172 _08744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_200_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30662_ clknet_leaf_142_clk _02397_ VGND VGND VPWR VPWR datamem.data_ram\[50\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_18384_ _05724_ _05733_ VGND VGND VPWR VPWR _05748_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_183 _09041_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15596_ net3432 _13220_ _14103_ VGND VGND VPWR VPWR _14106_ sky130_fd_sc_hd__mux2_1
XANTENNA_194 _09313_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17335_ net4413 _13262_ _04924_ VGND VGND VPWR VPWR _04931_ sky130_fd_sc_hd__mux2_1
X_32401_ clknet_leaf_247_clk _03823_ VGND VGND VPWR VPWR datamem.data_ram\[29\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_30593_ clknet_leaf_118_clk _02328_ VGND VGND VPWR VPWR datamem.data_ram\[53\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17266_ _14185_ net3319 _04887_ VGND VGND VPWR VPWR _04894_ sky130_fd_sc_hd__mux2_1
X_32332_ clknet_leaf_254_clk _03754_ VGND VGND VPWR VPWR datamem.data_ram\[31\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload103 clknet_leaf_89_clk VGND VGND VPWR VPWR clkload103/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_153_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload114 clknet_leaf_104_clk VGND VGND VPWR VPWR clkload114/Y sky130_fd_sc_hd__bufinv_16
X_19005_ _05290_ _05647_ VGND VGND VPWR VPWR _06339_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_12_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16217_ _13243_ VGND VGND VPWR VPWR _14463_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_168_4516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload125 clknet_leaf_252_clk VGND VGND VPWR VPWR clkload125/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_12_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32263_ clknet_leaf_270_clk _03685_ VGND VGND VPWR VPWR datamem.data_ram\[34\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_168_4527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17197_ _04857_ VGND VGND VPWR VPWR _01442_ sky130_fd_sc_hd__clkbuf_1
Xclkload136 clknet_leaf_241_clk VGND VGND VPWR VPWR clkload136/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_168_4538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload147 clknet_leaf_260_clk VGND VGND VPWR VPWR clkload147/Y sky130_fd_sc_hd__clkinv_4
X_31214_ clknet_leaf_33_clk _02917_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCD\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload158 clknet_leaf_285_clk VGND VGND VPWR VPWR clkload158/Y sky130_fd_sc_hd__clkinvlp_4
X_16148_ net2025 _13272_ _14407_ VGND VGND VPWR VPWR _14417_ sky130_fd_sc_hd__mux2_1
Xclkload169 clknet_leaf_270_clk VGND VGND VPWR VPWR clkload169/Y sky130_fd_sc_hd__clkinv_8
X_32194_ clknet_leaf_230_clk _03616_ VGND VGND VPWR VPWR datamem.data_ram\[36\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31145_ clknet_leaf_62_clk rvcpu.ALUResultE\[4\] VGND VGND VPWR VPWR rvcpu.dp.plem.ALUResultM\[4\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_41_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_90_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16079_ _14380_ VGND VGND VPWR VPWR _01983_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_227_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19907_ _07196_ _07201_ _06596_ VGND VGND VPWR VPWR _07202_ sky130_fd_sc_hd__o21a_1
Xhold2606 datamem.data_ram\[26\]\[8\] VGND VGND VPWR VPWR net3756 sky130_fd_sc_hd__dlygate4sd3_1
X_31076_ clknet_leaf_152_clk _02811_ VGND VGND VPWR VPWR datamem.data_ram\[9\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2617 datamem.data_ram\[5\]\[13\] VGND VGND VPWR VPWR net3767 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_3534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2628 datamem.data_ram\[29\]\[15\] VGND VGND VPWR VPWR net3778 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_127_3545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2639 datamem.data_ram\[56\]\[10\] VGND VGND VPWR VPWR net3789 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1905 datamem.data_ram\[10\]\[19\] VGND VGND VPWR VPWR net3055 sky130_fd_sc_hd__dlygate4sd3_1
X_30027_ net389 _01762_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[13\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_19838_ _06948_ VGND VGND VPWR VPWR _07133_ sky130_fd_sc_hd__clkbuf_8
Xhold1916 rvcpu.dp.rf.reg_file_arr\[0\]\[24\] VGND VGND VPWR VPWR net3066 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1927 rvcpu.dp.rf.reg_file_arr\[8\]\[1\] VGND VGND VPWR VPWR net3077 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1938 datamem.data_ram\[18\]\[8\] VGND VGND VPWR VPWR net3088 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1949 datamem.data_ram\[13\]\[30\] VGND VGND VPWR VPWR net3099 sky130_fd_sc_hd__dlygate4sd3_1
Xinput1 reset VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_4
X_19769_ datamem.data_ram\[24\]\[25\] _06697_ _06657_ datamem.data_ram\[25\]\[25\]
+ _07063_ VGND VGND VPWR VPWR _07064_ sky130_fd_sc_hd__o221a_1
XFILLER_0_79_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_48_clk clknet_5_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_48_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_155_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_88_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21800_ _08514_ _09039_ VGND VGND VPWR VPWR _09040_ sky130_fd_sc_hd__or2_1
XFILLER_0_211_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22780_ _09919_ _09920_ _09449_ VGND VGND VPWR VPWR _09921_ sky130_fd_sc_hd__mux2_2
XFILLER_0_210_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31978_ clknet_leaf_155_clk _03400_ VGND VGND VPWR VPWR datamem.data_ram\[53\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21731_ _08686_ _08974_ _08748_ VGND VGND VPWR VPWR _08975_ sky130_fd_sc_hd__o21ai_1
X_30929_ clknet_leaf_151_clk _02664_ VGND VGND VPWR VPWR datamem.data_ram\[40\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24450_ _10063_ VGND VGND VPWR VPWR _10413_ sky130_fd_sc_hd__buf_2
XFILLER_0_137_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21662_ _08813_ _08909_ _08689_ VGND VGND VPWR VPWR _08910_ sky130_fd_sc_hd__a21o_1
XFILLER_0_47_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_191_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23401_ _10151_ VGND VGND VPWR VPWR _01539_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20613_ _07900_ _07901_ _07902_ _07903_ VGND VGND VPWR VPWR _07904_ sky130_fd_sc_hd__a31o_1
X_24381_ _10369_ VGND VGND VPWR VPWR _02301_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21593_ _08565_ _08841_ _08844_ _08652_ VGND VGND VPWR VPWR _08845_ sky130_fd_sc_hd__o211a_1
XFILLER_0_7_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26120_ _11395_ VGND VGND VPWR VPWR _03013_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20544_ _07826_ VGND VGND VPWR VPWR _07835_ sky130_fd_sc_hd__buf_6
XFILLER_0_132_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26051_ _11353_ net1878 _11350_ _11354_ VGND VGND VPWR VPWR _02986_ sky130_fd_sc_hd__a31o_1
XFILLER_0_131_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20475_ datamem.data_ram\[39\]\[20\] _06706_ _07765_ _07766_ VGND VGND VPWR VPWR
+ _07767_ sky130_fd_sc_hd__o211a_1
XFILLER_0_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25002_ _10452_ net2820 _10715_ VGND VGND VPWR VPWR _10722_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22214_ rvcpu.dp.plfd.InstrD\[22\] VGND VGND VPWR VPWR _09380_ sky130_fd_sc_hd__buf_4
XFILLER_0_162_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23194_ _09240_ net4130 _10115_ VGND VGND VPWR VPWR _10118_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29810_ net1148 _01545_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[1\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22145_ _09342_ VGND VGND VPWR VPWR _01092_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_218_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24121__627 clknet_1_0__leaf__10260_ VGND VGND VPWR VPWR net753 sky130_fd_sc_hd__inv_2
X_29741_ net1087 _01476_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[21\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_26953_ _11849_ net1487 _11853_ _11858_ VGND VGND VPWR VPWR _03384_ sky130_fd_sc_hd__a31o_1
XFILLER_0_203_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22076_ _09290_ VGND VGND VPWR VPWR _09291_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_199_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25904_ net1627 _11181_ _11258_ _11270_ VGND VGND VPWR VPWR _02923_ sky130_fd_sc_hd__o211a_1
X_21027_ datamem.data_ram\[24\]\[31\] _06644_ _08313_ _07859_ _08315_ VGND VGND VPWR
+ VPWR _08316_ sky130_fd_sc_hd__o221a_1
X_26884_ _11813_ net1504 _11809_ _11814_ VGND VGND VPWR VPWR _03359_ sky130_fd_sc_hd__a31o_1
XFILLER_0_22_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29672_ net1018 _01407_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[23\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25835_ _11206_ _11207_ _11219_ VGND VGND VPWR VPWR _11220_ sky130_fd_sc_hd__and3_1
X_28623_ _12756_ net3324 _12805_ VGND VGND VPWR VPWR _12808_ sky130_fd_sc_hd__mux2_1
XFILLER_0_214_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_39_clk clknet_5_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_39_clk sky130_fd_sc_hd__clkbuf_8
X_25766_ _13463_ _13301_ _13294_ _13439_ VGND VGND VPWR VPWR _11166_ sky130_fd_sc_hd__a31o_1
XFILLER_0_198_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_195_5170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28554_ _12692_ net2649 _12768_ VGND VGND VPWR VPWR _12771_ sky130_fd_sc_hd__mux2_1
XFILLER_0_186_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_195_5181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27505_ _12151_ net2861 _12179_ VGND VGND VPWR VPWR _12184_ sky130_fd_sc_hd__mux2_1
X_24717_ _10566_ VGND VGND VPWR VPWR _02440_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28485_ _12391_ net1695 _12723_ _12726_ VGND VGND VPWR VPWR _04048_ sky130_fd_sc_hd__a31o_1
X_21929_ rvcpu.dp.rf.reg_file_arr\[20\]\[29\] rvcpu.dp.rf.reg_file_arr\[21\]\[29\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[29\] rvcpu.dp.rf.reg_file_arr\[23\]\[29\] _08778_
+ _08825_ VGND VGND VPWR VPWR _09162_ sky130_fd_sc_hd__mux4_1
X_25697_ _11105_ net1841 _11111_ _11120_ VGND VGND VPWR VPWR _02866_ sky130_fd_sc_hd__a31o_1
XFILLER_0_84_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_210_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15450_ _13553_ _13597_ _13564_ VGND VGND VPWR VPWR _13980_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_191_5078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27436_ _10668_ _12106_ _11713_ VGND VGND VPWR VPWR _12143_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_191_5089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24648_ _10398_ net1920 _10521_ VGND VGND VPWR VPWR _10528_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15381_ _13382_ _13319_ _13349_ _13914_ VGND VGND VPWR VPWR _13915_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_167_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27367_ _12089_ net4023 _12097_ VGND VGND VPWR VPWR _12102_ sky130_fd_sc_hd__mux2_1
X_24579_ _10454_ net3297 _10482_ VGND VGND VPWR VPWR _10490_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17120_ _14175_ net4040 _04815_ VGND VGND VPWR VPWR _04817_ sky130_fd_sc_hd__mux2_1
X_26318_ net2022 _11436_ VGND VGND VPWR VPWR _11492_ sky130_fd_sc_hd__and2_1
X_29106_ _13068_ VGND VGND VPWR VPWR _04327_ sky130_fd_sc_hd__clkbuf_1
X_27298_ _12061_ net1628 _12053_ _12062_ VGND VGND VPWR VPWR _03525_ sky130_fd_sc_hd__a31o_1
XFILLER_0_37_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_208_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29037_ _10047_ _13031_ VGND VGND VPWR VPWR _13032_ sky130_fd_sc_hd__and2_1
XFILLER_0_135_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17051_ _04780_ VGND VGND VPWR VPWR _01511_ sky130_fd_sc_hd__clkbuf_1
X_26249_ _11438_ _11458_ _11459_ net1296 VGND VGND VPWR VPWR _03079_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_150_4085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_4096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16002_ net2054 _13260_ _14333_ VGND VGND VPWR VPWR _14339_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_4402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_4413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17953_ _05324_ VGND VGND VPWR VPWR _05325_ sky130_fd_sc_hd__inv_2
X_29939_ net309 _01674_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[16\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_225_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16904_ net2489 _14455_ _04695_ VGND VGND VPWR VPWR _04702_ sky130_fd_sc_hd__mux2_1
X_32950_ clknet_leaf_214_clk _04372_ VGND VGND VPWR VPWR datamem.data_ram\[6\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_17884_ rvcpu.dp.plde.Rs1E\[2\] _13174_ VGND VGND VPWR VPWR _05257_ sky130_fd_sc_hd__and2b_1
XFILLER_0_228_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_1288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31901_ _04443_ net121 VGND VGND VPWR VPWR datamem.rd_data_mem\[6\] sky130_fd_sc_hd__dlxtn_1
X_19623_ _06918_ VGND VGND VPWR VPWR _06919_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_164_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16835_ _04665_ VGND VGND VPWR VPWR _01620_ sky130_fd_sc_hd__clkbuf_1
X_32881_ clknet_leaf_254_clk _04303_ VGND VGND VPWR VPWR datamem.data_ram\[10\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_122_3420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23740__331 clknet_1_1__leaf__10199_ VGND VGND VPWR VPWR net457 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_122_3431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19554_ datamem.data_ram\[8\]\[24\] _06820_ _06669_ datamem.data_ram\[15\]\[24\]
+ _06849_ VGND VGND VPWR VPWR _06850_ sky130_fd_sc_hd__o221a_1
X_31832_ clknet_leaf_213_clk _03286_ VGND VGND VPWR VPWR datamem.data_ram\[3\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16766_ net2362 _14453_ _04623_ VGND VGND VPWR VPWR _04629_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_177_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18505_ _05866_ _05692_ _05719_ _05733_ VGND VGND VPWR VPWR _05867_ sky130_fd_sc_hd__and4_1
X_15717_ _14182_ VGND VGND VPWR VPWR _02163_ sky130_fd_sc_hd__clkbuf_1
X_31763_ clknet_leaf_106_clk _03217_ VGND VGND VPWR VPWR datamem.data_ram\[18\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_16697_ _04592_ VGND VGND VPWR VPWR _01693_ sky130_fd_sc_hd__clkbuf_1
X_19485_ _06780_ VGND VGND VPWR VPWR _06781_ sky130_fd_sc_hd__buf_6
XFILLER_0_220_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_83_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30714_ clknet_leaf_136_clk _02449_ VGND VGND VPWR VPWR datamem.data_ram\[49\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_18436_ _05704_ VGND VGND VPWR VPWR _05799_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_200_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15648_ _14135_ net4083 _14131_ VGND VGND VPWR VPWR _14136_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31694_ clknet_leaf_39_clk _03152_ VGND VGND VPWR VPWR rvcpu.dp.pcreg.q\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18367_ _05731_ VGND VGND VPWR VPWR _05732_ sky130_fd_sc_hd__clkbuf_4
X_15579_ net2694 _13195_ _14092_ VGND VGND VPWR VPWR _14097_ sky130_fd_sc_hd__mux2_1
X_30645_ clknet_leaf_181_clk _02380_ VGND VGND VPWR VPWR datamem.data_ram\[51\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17318_ net3026 _13237_ _04913_ VGND VGND VPWR VPWR _04922_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30576_ clknet_leaf_188_clk _02311_ VGND VGND VPWR VPWR datamem.data_ram\[54\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18298_ _05662_ VGND VGND VPWR VPWR _05663_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_126_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_3279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32315_ clknet_leaf_240_clk _03737_ VGND VGND VPWR VPWR datamem.data_ram\[31\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17249_ _14168_ net3834 _04876_ VGND VGND VPWR VPWR _04885_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_92_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20260_ datamem.data_ram\[51\]\[19\] _06635_ _06620_ datamem.data_ram\[52\]\[19\]
+ VGND VGND VPWR VPWR _07553_ sky130_fd_sc_hd__o22a_1
XFILLER_0_222_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32246_ clknet_leaf_229_clk _03668_ VGND VGND VPWR VPWR datamem.data_ram\[34\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32177_ clknet_leaf_168_clk _03599_ VGND VGND VPWR VPWR datamem.data_ram\[37\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_20191_ datamem.data_ram\[46\]\[11\] _06717_ _06730_ datamem.data_ram\[43\]\[11\]
+ VGND VGND VPWR VPWR _07484_ sky130_fd_sc_hd__o22a_1
Xhold3104 rvcpu.dp.rf.reg_file_arr\[28\]\[27\] VGND VGND VPWR VPWR net4254 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3115 datamem.data_ram\[10\]\[27\] VGND VGND VPWR VPWR net4265 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3126 rvcpu.dp.rf.reg_file_arr\[0\]\[28\] VGND VGND VPWR VPWR net4276 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1300 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31128_ clknet_leaf_125_clk _02863_ VGND VGND VPWR VPWR datamem.data_ram\[25\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3137 rvcpu.dp.rf.reg_file_arr\[22\]\[22\] VGND VGND VPWR VPWR net4287 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3148 datamem.data_ram\[56\]\[19\] VGND VGND VPWR VPWR net4298 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2403 rvcpu.dp.rf.reg_file_arr\[25\]\[22\] VGND VGND VPWR VPWR net3553 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold3159 datamem.data_ram\[54\]\[26\] VGND VGND VPWR VPWR net4309 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2414 datamem.data_ram\[31\]\[9\] VGND VGND VPWR VPWR net3564 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2425 rvcpu.dp.rf.reg_file_arr\[30\]\[2\] VGND VGND VPWR VPWR net3575 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2436 datamem.data_ram\[62\]\[13\] VGND VGND VPWR VPWR net3586 sky130_fd_sc_hd__dlygate4sd3_1
X_31059_ clknet_leaf_91_clk _02794_ VGND VGND VPWR VPWR datamem.data_ram\[38\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1702 datamem.data_ram\[20\]\[26\] VGND VGND VPWR VPWR net2852 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2447 datamem.data_ram\[8\]\[16\] VGND VGND VPWR VPWR net3597 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1713 rvcpu.dp.rf.reg_file_arr\[13\]\[3\] VGND VGND VPWR VPWR net2863 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2458 rvcpu.dp.rf.reg_file_arr\[31\]\[6\] VGND VGND VPWR VPWR net3608 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_3998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1724 rvcpu.dp.rf.reg_file_arr\[18\]\[3\] VGND VGND VPWR VPWR net2874 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2469 datamem.data_ram\[28\]\[13\] VGND VGND VPWR VPWR net3619 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1735 rvcpu.dp.rf.reg_file_arr\[18\]\[26\] VGND VGND VPWR VPWR net2885 sky130_fd_sc_hd__dlygate4sd3_1
X_22901_ rvcpu.dp.rf.reg_file_arr\[8\]\[31\] rvcpu.dp.rf.reg_file_arr\[10\]\[31\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[31\] rvcpu.dp.rf.reg_file_arr\[11\]\[31\] _09483_
+ _09656_ VGND VGND VPWR VPWR _10036_ sky130_fd_sc_hd__mux4_1
Xhold1746 rvcpu.dp.rf.reg_file_arr\[20\]\[17\] VGND VGND VPWR VPWR net2896 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1757 datamem.data_ram\[9\]\[31\] VGND VGND VPWR VPWR net2907 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1768 rvcpu.dp.rf.reg_file_arr\[21\]\[1\] VGND VGND VPWR VPWR net2918 sky130_fd_sc_hd__dlygate4sd3_1
X_25620_ _11074_ VGND VGND VPWR VPWR _02835_ sky130_fd_sc_hd__clkbuf_1
Xhold1779 datamem.data_ram\[45\]\[11\] VGND VGND VPWR VPWR net2929 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22832_ rvcpu.dp.rf.reg_file_arr\[16\]\[28\] rvcpu.dp.rf.reg_file_arr\[17\]\[28\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[28\] rvcpu.dp.rf.reg_file_arr\[19\]\[28\] _09445_
+ _09447_ VGND VGND VPWR VPWR _09970_ sky130_fd_sc_hd__mux4_1
XFILLER_0_79_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25551_ _10758_ net2610 _11030_ VGND VGND VPWR VPWR _11034_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22763_ _09451_ _09904_ _09404_ VGND VGND VPWR VPWR _09905_ sky130_fd_sc_hd__o21a_1
XFILLER_0_195_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24502_ _10442_ datamem.data_ram\[52\]\[17\] _10440_ VGND VGND VPWR VPWR _10443_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_220_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28270_ _12606_ VGND VGND VPWR VPWR _03953_ sky130_fd_sc_hd__clkbuf_1
X_21714_ _08627_ _08954_ _08956_ _08958_ VGND VGND VPWR VPWR _08959_ sky130_fd_sc_hd__o2bb2a_1
X_25482_ _10064_ net35 _10996_ net1332 VGND VGND VPWR VPWR _02775_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22694_ _09510_ _09833_ _09835_ _09839_ _09525_ VGND VGND VPWR VPWR _09840_ sky130_fd_sc_hd__a311o_1
XFILLER_0_30_1300 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27221_ _11918_ VGND VGND VPWR VPWR _12022_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_137_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24433_ _09290_ VGND VGND VPWR VPWR _10400_ sky130_fd_sc_hd__buf_2
XFILLER_0_176_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21645_ _08692_ _08891_ _08893_ VGND VGND VPWR VPWR _08894_ sky130_fd_sc_hd__a21o_1
XFILLER_0_164_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27152_ _10075_ VGND VGND VPWR VPWR _11980_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_117_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24364_ _09310_ net4309 _10357_ VGND VGND VPWR VPWR _10360_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21576_ rvcpu.dp.rf.reg_file_arr\[28\]\[10\] rvcpu.dp.rf.reg_file_arr\[30\]\[10\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[10\] rvcpu.dp.rf.reg_file_arr\[31\]\[10\] _08629_
+ _08637_ VGND VGND VPWR VPWR _08828_ sky130_fd_sc_hd__mux4_1
XANTENNA_50 _06684_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_61 _06726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26103_ net1776 _11386_ VGND VGND VPWR VPWR _11387_ sky130_fd_sc_hd__and2_1
XANTENNA_72 _06776_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27083_ net1679 _11933_ _11935_ _10041_ VGND VGND VPWR VPWR _03437_ sky130_fd_sc_hd__o211a_1
X_20527_ datamem.data_ram\[18\]\[21\] _07203_ _07814_ _07817_ VGND VGND VPWR VPWR
+ _07818_ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_83 _06784_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_94 _06810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24295_ _09282_ net3428 _10316_ VGND VGND VPWR VPWR _10321_ sky130_fd_sc_hd__mux2_1
X_23910__467 clknet_1_0__leaf__10225_ VGND VGND VPWR VPWR net593 sky130_fd_sc_hd__inv_2
XFILLER_0_166_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26034_ _11086_ _11340_ VGND VGND VPWR VPWR _11344_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20458_ datamem.data_ram\[26\]\[20\] _06690_ _06633_ datamem.data_ram\[27\]\[20\]
+ _06600_ VGND VGND VPWR VPWR _07750_ sky130_fd_sc_hd__o221a_1
XFILLER_0_30_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_219_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20389_ datamem.data_ram\[21\]\[28\] _06768_ _06737_ datamem.data_ram\[19\]\[28\]
+ _07680_ VGND VGND VPWR VPWR _07681_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_205_5420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22128_ _09333_ VGND VGND VPWR VPWR _01084_ sky130_fd_sc_hd__clkbuf_1
X_24179__20 clknet_1_1__leaf__10265_ VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__inv_2
XFILLER_0_98_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27985_ _12450_ net3426 net76 VGND VGND VPWR VPWR _12451_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_201_5317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14950_ rvcpu.dp.pcreg.q\[9\] _13438_ VGND VGND VPWR VPWR _13499_ sky130_fd_sc_hd__nand2_2
X_29724_ net1070 _01459_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[22\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_201_5328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26936_ _11833_ _11842_ VGND VGND VPWR VPWR _11848_ sky130_fd_sc_hd__and2_1
X_22059_ rvcpu.dp.plem.WriteDataM\[3\] _09264_ _09265_ rvcpu.dp.plem.WriteDataM\[11\]
+ VGND VGND VPWR VPWR _09278_ sky130_fd_sc_hd__a22o_4
XTAP_TAPCELL_ROW_197_5221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_197_5232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2970 rvcpu.dp.rf.reg_file_arr\[3\]\[23\] VGND VGND VPWR VPWR net4120 sky130_fd_sc_hd__dlygate4sd3_1
X_14881_ rvcpu.dp.pcreg.q\[5\] _13280_ VGND VGND VPWR VPWR _13433_ sky130_fd_sc_hd__or2_1
Xhold2981 rvcpu.dp.rf.reg_file_arr\[16\]\[28\] VGND VGND VPWR VPWR net4131 sky130_fd_sc_hd__dlygate4sd3_1
X_24194__34 clknet_1_1__leaf__10266_ VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__inv_2
XFILLER_0_89_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29655_ net1001 _01390_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[24\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_26867_ _11803_ _11798_ VGND VGND VPWR VPWR _11804_ sky130_fd_sc_hd__and2_1
X_23266__912 clknet_1_1__leaf__10128_ VGND VGND VPWR VPWR net1038 sky130_fd_sc_hd__inv_2
Xhold2992 datamem.data_ram\[19\]\[9\] VGND VGND VPWR VPWR net4142 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_193_5118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_193_5129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16620_ _14151_ net3030 _04551_ VGND VGND VPWR VPWR _04552_ sky130_fd_sc_hd__mux2_1
X_28606_ _12692_ net3296 _12796_ VGND VGND VPWR VPWR _12799_ sky130_fd_sc_hd__mux2_1
X_25818_ net1761 _11181_ _11177_ _11205_ VGND VGND VPWR VPWR _02902_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_3_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26798_ _11676_ _11762_ VGND VGND VPWR VPWR _11763_ sky130_fd_sc_hd__and2_1
X_29586_ net940 _01321_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[26\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap52 _12041_ VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__buf_2
X_16551_ _14151_ net4114 _04514_ VGND VGND VPWR VPWR _04515_ sky130_fd_sc_hd__mux2_1
X_25749_ _11152_ VGND VGND VPWR VPWR _11153_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_134_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28537_ _09247_ VGND VGND VPWR VPWR _12760_ sky130_fd_sc_hd__buf_2
Xmax_cap63 _13103_ VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_4
XFILLER_0_85_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap74 _12519_ VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__buf_4
XFILLER_0_186_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap85 _12116_ VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__buf_4
Xmax_cap96 _12483_ VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__buf_4
XFILLER_0_214_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15502_ _13381_ _13876_ _13504_ VGND VGND VPWR VPWR _14030_ sky130_fd_sc_hd__o21ai_1
X_19270_ rvcpu.c.ad.funct7b5 VGND VGND VPWR VPWR _06570_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_156_4250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16482_ _04466_ VGND VGND VPWR VPWR _04478_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_85_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28468_ _12716_ VGND VGND VPWR VPWR _04041_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_5_0__f_clk clknet_2_0_0_clk VGND VGND VPWR VPWR clknet_5_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_73_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_210_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15433_ _13785_ _13962_ _13963_ _13458_ VGND VGND VPWR VPWR _13964_ sky130_fd_sc_hd__a31o_1
X_18221_ _05375_ _05373_ VGND VGND VPWR VPWR _05586_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_14_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27419_ _12131_ VGND VGND VPWR VPWR _03577_ sky130_fd_sc_hd__clkbuf_1
X_28399_ _12443_ net4328 _12669_ VGND VGND VPWR VPWR _12676_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_152_4136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_4147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30430_ net768 _02165_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[29\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_15364_ _13638_ _13537_ VGND VGND VPWR VPWR _13899_ sky130_fd_sc_hd__nor2_1
X_18152_ _05498_ _05516_ VGND VGND VPWR VPWR _05517_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17103_ _14158_ net2200 _04804_ VGND VGND VPWR VPWR _04808_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18083_ _05410_ _05419_ _05445_ _05450_ VGND VGND VPWR VPWR _05451_ sky130_fd_sc_hd__a31o_1
X_30361_ net707 _02096_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[3\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_15295_ _13430_ _13375_ _13348_ _13614_ VGND VGND VPWR VPWR _13833_ sky130_fd_sc_hd__a31o_1
XFILLER_0_68_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32100_ clknet_leaf_107_clk _03522_ VGND VGND VPWR VPWR datamem.data_ram\[23\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_17034_ _04771_ VGND VGND VPWR VPWR _01519_ sky130_fd_sc_hd__clkbuf_1
Xhold309 datamem.data_ram\[33\]\[6\] VGND VGND VPWR VPWR net1459 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30292_ net638 _02027_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[5\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_229_5987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32031_ clknet_leaf_128_clk _03453_ VGND VGND VPWR VPWR datamem.data_ram\[26\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_111_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_229_5998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_182_4855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23584__205 clknet_1_0__leaf__10177_ VGND VGND VPWR VPWR net331 sky130_fd_sc_hd__inv_2
XFILLER_0_42_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_182_4866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18985_ _05305_ _05555_ VGND VGND VPWR VPWR _06320_ sky130_fd_sc_hd__nor2_1
XFILLER_0_225_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17936_ rvcpu.dp.plem.ALUResultM\[14\] _05308_ _05176_ VGND VGND VPWR VPWR _05309_
+ sky130_fd_sc_hd__mux2_1
Xhold1009 rvcpu.dp.rf.reg_file_arr\[9\]\[30\] VGND VGND VPWR VPWR net2159 sky130_fd_sc_hd__dlygate4sd3_1
X_32933_ clknet_leaf_150_clk _04355_ VGND VGND VPWR VPWR datamem.data_ram\[7\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17867_ _05239_ VGND VGND VPWR VPWR _05240_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_75_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_1_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19606_ datamem.data_ram\[26\]\[8\] _06802_ _06669_ datamem.data_ram\[31\]\[8\] VGND
+ VGND VPWR VPWR _06902_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_1_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16818_ _04656_ VGND VGND VPWR VPWR _01628_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_85_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32864_ clknet_leaf_55_clk _04286_ VGND VGND VPWR VPWR datamem.data_ram\[11\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_141_3873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17798_ _13265_ _05179_ _05180_ net114 VGND VGND VPWR VPWR _05192_ sky130_fd_sc_hd__a31o_1
XFILLER_0_89_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_141_3884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31815_ clknet_leaf_104_clk _03269_ VGND VGND VPWR VPWR datamem.data_ram\[9\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19537_ datamem.data_ram\[37\]\[24\] _06823_ _06733_ _06832_ VGND VGND VPWR VPWR
+ _06833_ sky130_fd_sc_hd__o211a_1
XFILLER_0_159_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22989__695 clknet_1_0__leaf__10084_ VGND VGND VPWR VPWR net821 sky130_fd_sc_hd__inv_2
X_16749_ net3356 _14436_ _04612_ VGND VGND VPWR VPWR _04620_ sky130_fd_sc_hd__mux2_1
X_32795_ clknet_leaf_212_clk _04217_ VGND VGND VPWR VPWR datamem.data_ram\[13\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31746_ _04447_ net123 VGND VGND VPWR VPWR rvcpu.ALUControl\[0\] sky130_fd_sc_hd__dlxtn_1
XFILLER_0_14_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19468_ _06763_ VGND VGND VPWR VPWR _06764_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_186_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18419_ _05236_ _05659_ VGND VGND VPWR VPWR _05783_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31677_ clknet_leaf_9_clk net1267 VGND VGND VPWR VPWR rvcpu.dp.plmw.ALUResultW\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_19399_ _06645_ VGND VGND VPWR VPWR _06695_ sky130_fd_sc_hd__buf_6
XFILLER_0_5_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21430_ _08579_ VGND VGND VPWR VPWR _08689_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_100_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30628_ clknet_leaf_191_clk _02363_ VGND VGND VPWR VPWR datamem.data_ram\[52\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21361_ _08514_ _08569_ _08578_ _08579_ _08622_ VGND VGND VPWR VPWR _08623_ sky130_fd_sc_hd__o41a_1
X_30559_ clknet_leaf_197_clk _02294_ VGND VGND VPWR VPWR datamem.data_ram\[54\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_20312_ datamem.data_ram\[5\]\[4\] _07132_ _07600_ _07603_ VGND VGND VPWR VPWR _07604_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_163_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24080_ _09276_ net3996 _10249_ VGND VGND VPWR VPWR _10252_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21292_ _08553_ VGND VGND VPWR VPWR _08554_ sky130_fd_sc_hd__clkbuf_4
Xhold810 datamem.data_ram\[32\]\[31\] VGND VGND VPWR VPWR net1960 sky130_fd_sc_hd__dlygate4sd3_1
Xhold821 rvcpu.dp.rf.reg_file_arr\[8\]\[6\] VGND VGND VPWR VPWR net1971 sky130_fd_sc_hd__dlygate4sd3_1
X_23100__779 clknet_1_1__leaf__10103_ VGND VGND VPWR VPWR net905 sky130_fd_sc_hd__inv_2
Xhold832 rvcpu.dp.rf.reg_file_arr\[4\]\[21\] VGND VGND VPWR VPWR net1982 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold843 datamem.data_ram\[36\]\[30\] VGND VGND VPWR VPWR net1993 sky130_fd_sc_hd__dlygate4sd3_1
X_20243_ datamem.data_ram\[56\]\[3\] _06937_ _06926_ datamem.data_ram\[63\]\[3\] VGND
+ VGND VPWR VPWR _07536_ sky130_fd_sc_hd__a22o_1
X_32229_ clknet_leaf_170_clk _03651_ VGND VGND VPWR VPWR datamem.data_ram\[35\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold854 datamem.data_ram\[6\]\[30\] VGND VGND VPWR VPWR net2004 sky130_fd_sc_hd__dlygate4sd3_1
Xhold865 rvcpu.dp.rf.reg_file_arr\[5\]\[16\] VGND VGND VPWR VPWR net2015 sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 rvcpu.dp.rf.reg_file_arr\[3\]\[18\] VGND VGND VPWR VPWR net2026 sky130_fd_sc_hd__dlygate4sd3_1
Xhold887 rvcpu.dp.plfd.PCPlus4D\[21\] VGND VGND VPWR VPWR net2037 sky130_fd_sc_hd__dlygate4sd3_1
X_23747__337 clknet_1_0__leaf__10200_ VGND VGND VPWR VPWR net463 sky130_fd_sc_hd__inv_2
XFILLER_0_228_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20174_ datamem.data_ram\[16\]\[11\] _06837_ _06687_ datamem.data_ram\[20\]\[11\]
+ _07466_ VGND VGND VPWR VPWR _07467_ sky130_fd_sc_hd__o221a_1
Xhold898 datamem.data_ram\[36\]\[13\] VGND VGND VPWR VPWR net2048 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2200 datamem.data_ram\[17\]\[18\] VGND VGND VPWR VPWR net3350 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2211 datamem.data_ram\[54\]\[20\] VGND VGND VPWR VPWR net3361 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2222 datamem.data_ram\[28\]\[19\] VGND VGND VPWR VPWR net3372 sky130_fd_sc_hd__dlygate4sd3_1
X_24982_ _10711_ VGND VGND VPWR VPWR _02560_ sky130_fd_sc_hd__clkbuf_1
X_27770_ _08125_ net111 VGND VGND VPWR VPWR _12325_ sky130_fd_sc_hd__nor2_8
Xhold2233 datamem.data_ram\[8\]\[13\] VGND VGND VPWR VPWR net3383 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2244 datamem.data_ram\[23\]\[29\] VGND VGND VPWR VPWR net3394 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2255 datamem.data_ram\[39\]\[18\] VGND VGND VPWR VPWR net3405 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1510 datamem.data_ram\[54\]\[27\] VGND VGND VPWR VPWR net2660 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1521 rvcpu.dp.rf.reg_file_arr\[20\]\[9\] VGND VGND VPWR VPWR net2671 sky130_fd_sc_hd__dlygate4sd3_1
X_26721_ _11716_ VGND VGND VPWR VPWR _03294_ sky130_fd_sc_hd__clkbuf_1
Xhold2266 datamem.data_ram\[22\]\[29\] VGND VGND VPWR VPWR net3416 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2277 rvcpu.dp.rf.reg_file_arr\[19\]\[22\] VGND VGND VPWR VPWR net3427 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1532 datamem.data_ram\[4\]\[30\] VGND VGND VPWR VPWR net2682 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2288 datamem.data_ram\[24\]\[8\] VGND VGND VPWR VPWR net3438 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1543 rvcpu.dp.rf.reg_file_arr\[12\]\[21\] VGND VGND VPWR VPWR net2693 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2299 datamem.data_ram\[11\]\[12\] VGND VGND VPWR VPWR net3449 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1554 datamem.data_ram\[57\]\[29\] VGND VGND VPWR VPWR net2704 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1565 datamem.data_ram\[57\]\[11\] VGND VGND VPWR VPWR net2715 sky130_fd_sc_hd__dlygate4sd3_1
X_26652_ _11665_ net1456 _11662_ _11673_ VGND VGND VPWR VPWR _03268_ sky130_fd_sc_hd__a31o_1
XFILLER_0_165_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1576 rvcpu.dp.rf.reg_file_arr\[14\]\[31\] VGND VGND VPWR VPWR net2726 sky130_fd_sc_hd__dlygate4sd3_1
X_29440_ net802 _01175_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[30\]\[11\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__10221_ clknet_0__10221_ VGND VGND VPWR VPWR clknet_1_1__leaf__10221_
+ sky130_fd_sc_hd__clkbuf_16
Xhold1587 datamem.data_ram\[34\]\[22\] VGND VGND VPWR VPWR net2737 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1598 datamem.data_ram\[3\]\[18\] VGND VGND VPWR VPWR net2748 sky130_fd_sc_hd__dlygate4sd3_1
X_25603_ _11057_ net1479 _11053_ _11065_ VGND VGND VPWR VPWR _02827_ sky130_fd_sc_hd__a31o_1
XFILLER_0_196_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22815_ _09511_ _09953_ VGND VGND VPWR VPWR _09954_ sky130_fd_sc_hd__or2_1
X_29371_ clknet_leaf_195_clk _01106_ VGND VGND VPWR VPWR datamem.data_ram\[60\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__10152_ clknet_0__10152_ VGND VGND VPWR VPWR clknet_1_1__leaf__10152_
+ sky130_fd_sc_hd__clkbuf_16
X_26583_ _10739_ net2505 _11629_ VGND VGND VPWR VPWR _11637_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25534_ _10731_ net3649 net54 VGND VGND VPWR VPWR _11025_ sky130_fd_sc_hd__mux2_1
X_28322_ _12361_ net2780 _12632_ VGND VGND VPWR VPWR _12635_ sky130_fd_sc_hd__mux2_1
X_22746_ rvcpu.dp.rf.reg_file_arr\[24\]\[23\] rvcpu.dp.rf.reg_file_arr\[25\]\[23\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[23\] rvcpu.dp.rf.reg_file_arr\[27\]\[23\] _09392_
+ _09394_ VGND VGND VPWR VPWR _09889_ sky130_fd_sc_hd__mux4_1
XFILLER_0_94_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__10083_ clknet_0__10083_ VGND VGND VPWR VPWR clknet_1_1__leaf__10083_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_39_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28253_ _12596_ VGND VGND VPWR VPWR _03946_ sky130_fd_sc_hd__clkbuf_1
X_25465_ _10954_ net1388 _10984_ _10988_ VGND VGND VPWR VPWR _02766_ sky130_fd_sc_hd__a31o_1
XFILLER_0_176_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22677_ rvcpu.dp.rf.reg_file_arr\[4\]\[19\] rvcpu.dp.rf.reg_file_arr\[5\]\[19\] rvcpu.dp.rf.reg_file_arr\[6\]\[19\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[19\] _09604_ _09716_ VGND VGND VPWR VPWR _09824_
+ sky130_fd_sc_hd__mux4_1
X_27204_ _11972_ _12008_ VGND VGND VPWR VPWR _12012_ sky130_fd_sc_hd__and2_1
XFILLER_0_165_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24416_ _10388_ net4423 _10386_ VGND VGND VPWR VPWR _10389_ sky130_fd_sc_hd__mux2_1
XFILLER_0_191_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28184_ _12559_ VGND VGND VPWR VPWR _03914_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21628_ rvcpu.dp.rf.reg_file_arr\[4\]\[12\] rvcpu.dp.rf.reg_file_arr\[5\]\[12\] rvcpu.dp.rf.reg_file_arr\[6\]\[12\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[12\] _08687_ _08649_ VGND VGND VPWR VPWR _08878_
+ sky130_fd_sc_hd__mux4_1
X_25396_ _10938_ net1641 _10949_ _10952_ VGND VGND VPWR VPWR _02733_ sky130_fd_sc_hd__a31o_1
X_23296__938 clknet_1_0__leaf__10132_ VGND VGND VPWR VPWR net1064 sky130_fd_sc_hd__inv_2
XFILLER_0_180_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27135_ _11968_ _11966_ VGND VGND VPWR VPWR _11969_ sky130_fd_sc_hd__and2_1
XFILLER_0_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24347_ _09276_ net3389 _10348_ VGND VGND VPWR VPWR _10351_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21559_ rvcpu.dp.rf.reg_file_arr\[0\]\[9\] rvcpu.dp.rf.reg_file_arr\[1\]\[9\] rvcpu.dp.rf.reg_file_arr\[2\]\[9\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[9\] _08810_ _08811_ VGND VGND VPWR VPWR _08812_ sky130_fd_sc_hd__mux4_1
XFILLER_0_90_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27066_ _11825_ _11924_ VGND VGND VPWR VPWR _11926_ sky130_fd_sc_hd__and2_1
X_15080_ _13358_ _13607_ _13465_ _13493_ VGND VGND VPWR VPWR _13626_ sky130_fd_sc_hd__or4_1
X_24127__633 clknet_1_1__leaf__10260_ VGND VGND VPWR VPWR net759 sky130_fd_sc_hd__inv_2
XFILLER_0_205_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24278_ _09248_ net3362 _10307_ VGND VGND VPWR VPWR _10312_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26017_ net22 _11152_ VGND VGND VPWR VPWR _11334_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_224_5862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_224_5873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_270_clk clknet_5_19__leaf_clk VGND VGND VPWR VPWR clknet_leaf_270_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_209_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18770_ _05886_ _06107_ _06119_ VGND VGND VPWR VPWR _06120_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_8_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27968_ _09247_ VGND VGND VPWR VPWR _12439_ sky130_fd_sc_hd__clkbuf_2
X_15982_ _14328_ VGND VGND VPWR VPWR _02036_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29707_ net1053 _01442_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[22\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_17721_ _05135_ VGND VGND VPWR VPWR _01180_ sky130_fd_sc_hd__clkbuf_1
X_14933_ _13313_ _13283_ VGND VGND VPWR VPWR _13482_ sky130_fd_sc_hd__or2_1
X_26919_ _10075_ VGND VGND VPWR VPWR _11837_ sky130_fd_sc_hd__clkbuf_4
X_27899_ _12391_ net1559 _12393_ _12400_ VGND VGND VPWR VPWR _03788_ sky130_fd_sc_hd__a31o_1
XFILLER_0_215_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29638_ net984 _01373_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[24\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_17652_ net2061 _13228_ _05093_ VGND VGND VPWR VPWR _05099_ sky130_fd_sc_hd__mux2_1
X_14864_ _13369_ _13415_ VGND VGND VPWR VPWR _13416_ sky130_fd_sc_hd__nor2_2
XFILLER_0_188_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_225_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_19_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16603_ _14135_ net2535 _04540_ VGND VGND VPWR VPWR _04543_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_19_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14795_ _13347_ VGND VGND VPWR VPWR _13348_ sky130_fd_sc_hd__buf_4
XFILLER_0_159_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29569_ net923 _01304_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[26\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_17583_ _05062_ VGND VGND VPWR VPWR _01245_ sky130_fd_sc_hd__clkbuf_1
X_31600_ clknet_leaf_68_clk net1151 VGND VGND VPWR VPWR rvcpu.dp.plmw.PCPlus4W\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_19322_ _06617_ VGND VGND VPWR VPWR _06618_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16534_ _14135_ net3762 _04503_ VGND VGND VPWR VPWR _04506_ sky130_fd_sc_hd__mux2_1
X_32580_ clknet_leaf_232_clk _04002_ VGND VGND VPWR VPWR datamem.data_ram\[21\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_682 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_175_4692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31531_ clknet_leaf_27_clk net1200 VGND VGND VPWR VPWR rvcpu.dp.plem.PCPlus4M\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_19253_ _06547_ _06549_ VGND VGND VPWR VPWR _06556_ sky130_fd_sc_hd__or2b_1
XFILLER_0_112_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16465_ _04469_ VGND VGND VPWR VPWR _01810_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18204_ _05565_ _05501_ _05568_ VGND VGND VPWR VPWR _05569_ sky130_fd_sc_hd__o21a_1
XFILLER_0_26_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15416_ _13533_ _13640_ _13853_ _13947_ VGND VGND VPWR VPWR _13948_ sky130_fd_sc_hd__o31ai_1
X_19184_ rvcpu.dp.plde.ImmExtE\[21\] rvcpu.dp.plde.PCE\[21\] VGND VGND VPWR VPWR _06496_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_171_4589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31462_ clknet_leaf_5_clk rvcpu.dp.SrcBFW_Mux.y\[20\] VGND VGND VPWR VPWR rvcpu.dp.plem.WriteDataM\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16396_ net2313 _14426_ _14561_ VGND VGND VPWR VPWR _14564_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15347_ _13291_ _13343_ _13352_ _13759_ VGND VGND VPWR VPWR _13883_ sky130_fd_sc_hd__a211o_1
X_18135_ rvcpu.dp.plde.ImmExtE\[17\] rvcpu.dp.SrcBFW_Mux.y\[17\] _05278_ VGND VGND
+ VPWR VPWR _05501_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_113_3205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30413_ net751 _02148_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[31\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_31393_ clknet_leaf_40_clk _03096_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCE\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__10241_ clknet_0__10241_ VGND VGND VPWR VPWR clknet_1_0__leaf__10241_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_78_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15278_ _13599_ _13536_ _13802_ VGND VGND VPWR VPWR _13817_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_184_4906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18066_ _05327_ _05330_ VGND VGND VPWR VPWR _05434_ sky130_fd_sc_hd__or2_1
Xhold106 rvcpu.dp.plem.RdM\[1\] VGND VGND VPWR VPWR net1256 sky130_fd_sc_hd__dlygate4sd3_1
X_30344_ net690 _02079_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[4\]\[27\] sky130_fd_sc_hd__dfxtp_1
Xhold117 rvcpu.dp.plem.ALUResultM\[25\] VGND VGND VPWR VPWR net1267 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_184_4917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__10172_ clknet_0__10172_ VGND VGND VPWR VPWR clknet_1_0__leaf__10172_
+ sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold128 rvcpu.dp.plde.RdE\[2\] VGND VGND VPWR VPWR net1278 sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 rvcpu.dp.hu.ResultSrcE0 VGND VGND VPWR VPWR net1289 sky130_fd_sc_hd__dlygate4sd3_1
X_17017_ _04762_ VGND VGND VPWR VPWR _01527_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_74_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30275_ net629 _02010_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[6\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32014_ clknet_leaf_128_clk _03436_ VGND VGND VPWR VPWR datamem.data_ram\[27\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_261_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_261_clk
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_107_Right_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18968_ _06055_ _06296_ _06304_ VGND VGND VPWR VPWR _06305_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_143_3924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17919_ _05291_ VGND VGND VPWR VPWR _05292_ sky130_fd_sc_hd__clkbuf_4
X_18899_ _05627_ _06228_ _05461_ VGND VGND VPWR VPWR _06240_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_33_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20930_ _08218_ _08219_ _07839_ VGND VGND VPWR VPWR _08220_ sky130_fd_sc_hd__mux2_1
X_32916_ clknet_leaf_154_clk _04338_ VGND VGND VPWR VPWR datamem.data_ram\[0\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_221_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32847_ clknet_leaf_85_clk _04269_ VGND VGND VPWR VPWR datamem.data_ram\[7\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_20861_ _06967_ _06595_ VGND VGND VPWR VPWR _08151_ sky130_fd_sc_hd__nand2_4
XFILLER_0_49_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22600_ rvcpu.dp.rf.reg_file_arr\[0\]\[15\] rvcpu.dp.rf.reg_file_arr\[1\]\[15\] rvcpu.dp.rf.reg_file_arr\[2\]\[15\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[15\] _09714_ _09585_ VGND VGND VPWR VPWR _09751_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_18_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32778_ clknet_leaf_159_clk _04200_ VGND VGND VPWR VPWR datamem.data_ram\[14\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_102_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20792_ _06753_ _08072_ _08074_ _08081_ VGND VGND VPWR VPWR _08082_ sky130_fd_sc_hd__a31o_1
XFILLER_0_77_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22531_ _09482_ _09685_ VGND VGND VPWR VPWR _09686_ sky130_fd_sc_hd__or2_1
X_23180__851 clknet_1_0__leaf__10111_ VGND VGND VPWR VPWR net977 sky130_fd_sc_hd__inv_2
X_31729_ net178 _03187_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[9\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25250_ _10739_ net2334 _10857_ VGND VGND VPWR VPWR _10865_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22462_ _09618_ _09619_ _09380_ VGND VGND VPWR VPWR _09620_ sky130_fd_sc_hd__mux2_2
XFILLER_0_106_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24201_ _09298_ net2515 _10270_ VGND VGND VPWR VPWR _10271_ sky130_fd_sc_hd__mux2_1
X_21413_ _08623_ VGND VGND VPWR VPWR _08672_ sky130_fd_sc_hd__buf_2
X_25181_ _10827_ VGND VGND VPWR VPWR _02643_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22393_ _09429_ _09551_ _09554_ _09438_ VGND VGND VPWR VPWR _09555_ sky130_fd_sc_hd__a211o_1
X_23452__102 clknet_1_0__leaf__10156_ VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__inv_2
X_21344_ _05239_ _06195_ _06209_ rvcpu.ALUResultE\[18\] VGND VGND VPWR VPWR _08606_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_170_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28940_ _12766_ net1954 _12968_ VGND VGND VPWR VPWR _12976_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23981__516 clknet_1_1__leaf__10239_ VGND VGND VPWR VPWR net642 sky130_fd_sc_hd__inv_2
Xhold640 datamem.data_ram\[0\]\[6\] VGND VGND VPWR VPWR net1790 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21275_ _08536_ VGND VGND VPWR VPWR _08537_ sky130_fd_sc_hd__clkbuf_8
Xhold651 rvcpu.dp.plfd.PCD\[4\] VGND VGND VPWR VPWR net1801 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold662 datamem.data_ram\[10\]\[1\] VGND VGND VPWR VPWR net1812 sky130_fd_sc_hd__dlygate4sd3_1
X_20226_ datamem.data_ram\[8\]\[3\] _06935_ _06946_ datamem.data_ram\[9\]\[3\] VGND
+ VGND VPWR VPWR _07519_ sky130_fd_sc_hd__a22o_1
Xhold673 rvcpu.dp.pcreg.q\[30\] VGND VGND VPWR VPWR net1823 sky130_fd_sc_hd__dlygate4sd3_1
Xhold684 datamem.data_ram\[9\]\[0\] VGND VGND VPWR VPWR net1834 sky130_fd_sc_hd__dlygate4sd3_1
X_28871_ _12939_ VGND VGND VPWR VPWR _04221_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_228_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold695 datamem.data_ram\[61\]\[4\] VGND VGND VPWR VPWR net1845 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_252_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_252_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_5_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27822_ _12157_ net2418 net78 VGND VGND VPWR VPWR _12354_ sky130_fd_sc_hd__mux2_1
XFILLER_0_229_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20157_ datamem.data_ram\[31\]\[27\] _06671_ _06687_ datamem.data_ram\[28\]\[27\]
+ VGND VGND VPWR VPWR _07450_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_5_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2030 rvcpu.dp.rf.reg_file_arr\[14\]\[6\] VGND VGND VPWR VPWR net3180 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2041 rvcpu.dp.rf.reg_file_arr\[31\]\[9\] VGND VGND VPWR VPWR net3191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2052 datamem.data_ram\[51\]\[16\] VGND VGND VPWR VPWR net3202 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2063 datamem.data_ram\[2\]\[26\] VGND VGND VPWR VPWR net3213 sky130_fd_sc_hd__dlygate4sd3_1
X_27753_ _10838_ _12106_ _12260_ VGND VGND VPWR VPWR _12316_ sky130_fd_sc_hd__a21oi_4
X_24965_ _10396_ net3679 _10696_ VGND VGND VPWR VPWR _10702_ sky130_fd_sc_hd__mux2_1
Xhold2074 datamem.data_ram\[15\]\[21\] VGND VGND VPWR VPWR net3224 sky130_fd_sc_hd__dlygate4sd3_1
X_20088_ datamem.data_ram\[52\]\[10\] _06805_ _07380_ _07381_ VGND VGND VPWR VPWR
+ _07382_ sky130_fd_sc_hd__o211a_1
Xhold1340 datamem.data_ram\[30\]\[17\] VGND VGND VPWR VPWR net2490 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2085 rvcpu.dp.rf.reg_file_arr\[13\]\[17\] VGND VGND VPWR VPWR net3235 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2096 datamem.data_ram\[3\]\[25\] VGND VGND VPWR VPWR net3246 sky130_fd_sc_hd__dlygate4sd3_1
X_26704_ _10816_ net2764 _11704_ VGND VGND VPWR VPWR _11707_ sky130_fd_sc_hd__mux2_1
Xhold1351 datamem.data_ram\[16\]\[14\] VGND VGND VPWR VPWR net2501 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1362 datamem.data_ram\[28\]\[25\] VGND VGND VPWR VPWR net2512 sky130_fd_sc_hd__dlygate4sd3_1
X_24896_ _10450_ net2884 _10659_ VGND VGND VPWR VPWR _10665_ sky130_fd_sc_hd__mux2_1
X_27684_ _06997_ VGND VGND VPWR VPWR _12279_ sky130_fd_sc_hd__buf_8
Xhold1373 rvcpu.dp.rf.reg_file_arr\[20\]\[28\] VGND VGND VPWR VPWR net2523 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1384 rvcpu.dp.rf.reg_file_arr\[22\]\[11\] VGND VGND VPWR VPWR net2534 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1395 datamem.data_ram\[22\]\[12\] VGND VGND VPWR VPWR net2545 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_502 _11603_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29423_ clknet_leaf_97_clk _01158_ VGND VGND VPWR VPWR datamem.data_ram\[5\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__10204_ clknet_0__10204_ VGND VGND VPWR VPWR clknet_1_1__leaf__10204_
+ sky130_fd_sc_hd__clkbuf_16
X_26635_ _11078_ _11663_ VGND VGND VPWR VPWR _11664_ sky130_fd_sc_hd__and2_1
XANTENNA_513 _13222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_524 _13257_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_170_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_535 rvcpu.dp.plmw.ReadDataW\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_185_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_546 _06780_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_212_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29354_ clknet_leaf_141_clk _01089_ VGND VGND VPWR VPWR datamem.data_ram\[61\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__10135_ clknet_0__10135_ VGND VGND VPWR VPWR clknet_1_1__leaf__10135_
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_557 _07859_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_184_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23778_ clknet_1_0__leaf__10203_ VGND VGND VPWR VPWR _10204_ sky130_fd_sc_hd__buf_1
X_26566_ _10826_ net2214 _11620_ VGND VGND VPWR VPWR _11628_ sky130_fd_sc_hd__mux2_1
XANTENNA_568 _06610_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_184_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28305_ _12452_ net4169 net72 VGND VGND VPWR VPWR _12626_ sky130_fd_sc_hd__mux2_1
X_25517_ _10067_ _11010_ VGND VGND VPWR VPWR _11015_ sky130_fd_sc_hd__and2_1
XFILLER_0_177_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23304__945 clknet_1_1__leaf__10133_ VGND VGND VPWR VPWR net1071 sky130_fd_sc_hd__inv_2
XFILLER_0_55_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22729_ _09391_ _09872_ VGND VGND VPWR VPWR _09873_ sky130_fd_sc_hd__or2_1
X_29285_ _09317_ net3285 _13159_ VGND VGND VPWR VPWR _13164_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_188_5006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23916__473 clknet_1_1__leaf__10225_ VGND VGND VPWR VPWR net599 sky130_fd_sc_hd__inv_2
X_16250_ _14485_ VGND VGND VPWR VPWR _01917_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_188_5017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25448_ _10780_ _10981_ VGND VGND VPWR VPWR _10982_ sky130_fd_sc_hd__nor2_2
X_28236_ _12587_ VGND VGND VPWR VPWR _03938_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_192_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15201_ _13740_ _13499_ _13742_ VGND VGND VPWR VPWR _13743_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_213_5596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_209_Right_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16181_ net2531 _14438_ _14422_ VGND VGND VPWR VPWR _14439_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25379_ _10938_ net1517 _10934_ _10941_ VGND VGND VPWR VPWR _02727_ sky130_fd_sc_hd__a31o_1
X_28167_ _12550_ VGND VGND VPWR VPWR _03906_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23615__234 clknet_1_0__leaf__10179_ VGND VGND VPWR VPWR net360 sky130_fd_sc_hd__inv_2
XFILLER_0_35_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15132_ _13372_ _13336_ _13510_ _13401_ VGND VGND VPWR VPWR _13677_ sky130_fd_sc_hd__o22a_1
X_27118_ _11829_ _11953_ VGND VGND VPWR VPWR _11958_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28098_ _12454_ net3801 net75 VGND VGND VPWR VPWR _12514_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_226_5913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_226_5924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15063_ _13335_ _13294_ VGND VGND VPWR VPWR _13610_ sky130_fd_sc_hd__nand2_1
X_27049_ _11829_ _11911_ VGND VGND VPWR VPWR _11915_ sky130_fd_sc_hd__and2_1
X_19940_ datamem.data_ram\[34\]\[18\] _06613_ _07229_ _07233_ VGND VGND VPWR VPWR
+ _07234_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_147_4013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_4024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_4035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30060_ net422 _01795_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[12\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_19871_ datamem.data_ram\[30\]\[1\] _07159_ _06949_ datamem.data_ram\[25\]\[1\] VGND
+ VGND VPWR VPWR _07166_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_243_clk clknet_5_17__leaf_clk VGND VGND VPWR VPWR clknet_leaf_243_clk
+ sky130_fd_sc_hd__clkbuf_8
X_18822_ _05504_ _05513_ _05616_ _05569_ VGND VGND VPWR VPWR _06168_ sky130_fd_sc_hd__o31a_1
XFILLER_0_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23350__987 clknet_1_1__leaf__10137_ VGND VGND VPWR VPWR net1113 sky130_fd_sc_hd__inv_2
XFILLER_0_208_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18753_ _06087_ _06088_ _06103_ VGND VGND VPWR VPWR rvcpu.ALUResultE\[13\] sky130_fd_sc_hd__a21o_1
XFILLER_0_218_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15965_ _14319_ VGND VGND VPWR VPWR _02044_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_106_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17704_ _05126_ VGND VGND VPWR VPWR _01188_ sky130_fd_sc_hd__clkbuf_1
X_14916_ _13412_ VGND VGND VPWR VPWR _13466_ sky130_fd_sc_hd__clkbuf_4
X_30962_ clknet_leaf_91_clk _02697_ VGND VGND VPWR VPWR datamem.data_ram\[3\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_18684_ _05419_ _06036_ _05239_ VGND VGND VPWR VPWR _06038_ sky130_fd_sc_hd__o21a_1
X_15896_ net3873 _13204_ _14275_ VGND VGND VPWR VPWR _14283_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_177_4732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32701_ clknet_leaf_237_clk _04123_ VGND VGND VPWR VPWR datamem.data_ram\[17\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_177_4743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17635_ net2012 _13203_ _05082_ VGND VGND VPWR VPWR _05090_ sky130_fd_sc_hd__mux2_1
X_14847_ rvcpu.dp.pcreg.q\[3\] rvcpu.dp.pcreg.q\[2\] VGND VGND VPWR VPWR _13400_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_177_4754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30893_ clknet_leaf_155_clk _02628_ VGND VGND VPWR VPWR datamem.data_ram\[41\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32632_ clknet_leaf_90_clk _04054_ VGND VGND VPWR VPWR datamem.data_ram\[1\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17566_ _05053_ VGND VGND VPWR VPWR _01253_ sky130_fd_sc_hd__clkbuf_1
X_14778_ rvcpu.dp.pcreg.q\[6\] VGND VGND VPWR VPWR _13331_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_19_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_175_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19305_ _06600_ VGND VGND VPWR VPWR _06601_ sky130_fd_sc_hd__buf_8
X_16517_ _04496_ VGND VGND VPWR VPWR _01785_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_191_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32563_ clknet_leaf_171_clk _03985_ VGND VGND VPWR VPWR datamem.data_ram\[22\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_17497_ _13201_ net3325 _05010_ VGND VGND VPWR VPWR _05017_ sky130_fd_sc_hd__mux2_1
X_23244__892 clknet_1_0__leaf__10126_ VGND VGND VPWR VPWR net1018 sky130_fd_sc_hd__inv_2
XFILLER_0_156_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31514_ clknet_leaf_51_clk net1226 VGND VGND VPWR VPWR rvcpu.dp.plem.PCPlus4M\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_190_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19236_ rvcpu.dp.plde.ImmExtE\[28\] rvcpu.dp.plde.PCE\[28\] VGND VGND VPWR VPWR _06541_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16448_ net2485 _14478_ _04451_ VGND VGND VPWR VPWR _04459_ sky130_fd_sc_hd__mux2_1
X_32494_ clknet_leaf_74_clk _03916_ VGND VGND VPWR VPWR datamem.data_ram\[25\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_3750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_136_3761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19167_ rvcpu.dp.plde.ImmExtE\[19\] rvcpu.dp.plde.PCE\[19\] VGND VGND VPWR VPWR _06481_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_144_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31445_ clknet_leaf_76_clk rvcpu.dp.SrcBFW_Mux.y\[3\] VGND VGND VPWR VPWR rvcpu.dp.plem.WriteDataM\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_82_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16379_ _14554_ VGND VGND VPWR VPWR _01849_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18118_ rvcpu.dp.plde.ImmExtE\[19\] rvcpu.dp.SrcBFW_Mux.y\[19\] _05278_ VGND VGND
+ VPWR VPWR _05485_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_132_3658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_3669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19098_ _06420_ VGND VGND VPWR VPWR rvcpu.dp.lAuiPCE\[10\] sky130_fd_sc_hd__clkbuf_1
X_31376_ clknet_leaf_22_clk _03079_ VGND VGND VPWR VPWR rvcpu.dp.plde.ImmExtE\[25\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f__10224_ clknet_0__10224_ VGND VGND VPWR VPWR clknet_1_0__leaf__10224_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_170_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18049_ _05416_ _05417_ VGND VGND VPWR VPWR _05418_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30327_ net673 _02062_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[4\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_197_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__10155_ clknet_0__10155_ VGND VGND VPWR VPWR clknet_1_0__leaf__10155_
+ sky130_fd_sc_hd__clkbuf_16
X_21060_ datamem.data_ram\[40\]\[31\] datamem.data_ram\[41\]\[31\] datamem.data_ram\[42\]\[31\]
+ datamem.data_ram\[43\]\[31\] _07824_ _07819_ VGND VGND VPWR VPWR _08349_ sky130_fd_sc_hd__mux4_1
XFILLER_0_1_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30258_ net612 _01993_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[6\]\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_35_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__10086_ clknet_0__10086_ VGND VGND VPWR VPWR clknet_1_0__leaf__10086_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_201_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20011_ datamem.data_ram\[48\]\[2\] _06937_ _06954_ datamem.data_ram\[52\]\[2\] VGND
+ VGND VPWR VPWR _07305_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_35_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_234_clk clknet_5_20__leaf_clk VGND VGND VPWR VPWR clknet_leaf_234_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_35_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30189_ net543 _01924_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[8\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_225_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24750_ _10584_ VGND VGND VPWR VPWR _02455_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21962_ _08623_ _09185_ _09189_ _09193_ VGND VGND VPWR VPWR _09194_ sky130_fd_sc_hd__and4_1
XFILLER_0_193_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20913_ datamem.data_ram\[22\]\[22\] _07028_ _07019_ datamem.data_ram\[21\]\[22\]
+ _08202_ VGND VGND VPWR VPWR _08203_ sky130_fd_sc_hd__o221a_1
X_23562__185 clknet_1_1__leaf__10175_ VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__inv_2
X_24681_ _10547_ VGND VGND VPWR VPWR _02423_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21893_ rvcpu.dp.rf.reg_file_arr\[20\]\[27\] rvcpu.dp.rf.reg_file_arr\[21\]\[27\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[27\] rvcpu.dp.rf.reg_file_arr\[23\]\[27\] _08516_
+ _08518_ VGND VGND VPWR VPWR _09128_ sky130_fd_sc_hd__mux4_1
XFILLER_0_222_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_178_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_221_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26420_ net2171 _11542_ _11557_ _11534_ VGND VGND VPWR VPWR _03152_ sky130_fd_sc_hd__o211a_1
X_23632_ _10142_ _09269_ _09361_ VGND VGND VPWR VPWR _10182_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_179_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20844_ datamem.data_ram\[16\]\[14\] datamem.data_ram\[17\]\[14\] datamem.data_ram\[18\]\[14\]
+ datamem.data_ram\[19\]\[14\] _07826_ _07821_ VGND VGND VPWR VPWR _08134_ sky130_fd_sc_hd__mux4_1
XFILLER_0_194_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26351_ _10073_ _11507_ _11508_ net1330 VGND VGND VPWR VPWR _03132_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23026__728 clknet_1_0__leaf__10088_ VGND VGND VPWR VPWR net854 sky130_fd_sc_hd__inv_2
X_20775_ datamem.data_ram\[58\]\[6\] _07136_ _07137_ datamem.data_ram\[59\]\[6\] VGND
+ VGND VPWR VPWR _08065_ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25302_ _10764_ net2234 _10887_ VGND VGND VPWR VPWR _10894_ sky130_fd_sc_hd__mux2_1
XFILLER_0_175_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22514_ _09476_ _09667_ _09669_ _09474_ VGND VGND VPWR VPWR _09670_ sky130_fd_sc_hd__o211a_1
XFILLER_0_107_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26282_ _11473_ VGND VGND VPWR VPWR _03098_ sky130_fd_sc_hd__clkbuf_1
X_29070_ _10777_ _10960_ _12977_ VGND VGND VPWR VPWR _13049_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_88_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25233_ _10766_ net2020 _10848_ VGND VGND VPWR VPWR _10856_ sky130_fd_sc_hd__mux2_1
X_28021_ _12472_ VGND VGND VPWR VPWR _03838_ sky130_fd_sc_hd__clkbuf_1
X_22445_ _09401_ VGND VGND VPWR VPWR _09604_ sky130_fd_sc_hd__buf_4
XFILLER_0_88_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25164_ _09309_ VGND VGND VPWR VPWR _10816_ sky130_fd_sc_hd__buf_2
X_22376_ _09538_ VGND VGND VPWR VPWR _01127_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21327_ rvcpu.dp.plfd.InstrD\[24\] VGND VGND VPWR VPWR _08589_ sky130_fd_sc_hd__inv_2
X_25095_ _10780_ _10779_ VGND VGND VPWR VPWR _10781_ sky130_fd_sc_hd__nor2_2
X_29972_ net342 _01707_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[15\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_24046_ clknet_1_1__leaf__10244_ VGND VGND VPWR VPWR _10246_ sky130_fd_sc_hd__buf_1
X_28923_ _12702_ net1987 _12959_ VGND VGND VPWR VPWR _12967_ sky130_fd_sc_hd__mux2_1
Xhold470 datamem.data_ram\[18\]\[2\] VGND VGND VPWR VPWR net1620 sky130_fd_sc_hd__dlygate4sd3_1
X_21258_ rvcpu.dp.rf.reg_file_arr\[16\]\[0\] rvcpu.dp.rf.reg_file_arr\[17\]\[0\] rvcpu.dp.rf.reg_file_arr\[18\]\[0\]
+ rvcpu.dp.rf.reg_file_arr\[19\]\[0\] _08517_ _08519_ VGND VGND VPWR VPWR _08520_
+ sky130_fd_sc_hd__mux4_1
Xhold481 datamem.data_ram\[49\]\[6\] VGND VGND VPWR VPWR net1631 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold492 datamem.data_ram\[8\]\[5\] VGND VGND VPWR VPWR net1642 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_221_5810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_225_clk clknet_5_21__leaf_clk VGND VGND VPWR VPWR clknet_leaf_225_clk
+ sky130_fd_sc_hd__clkbuf_8
X_20209_ datamem.data_ram\[51\]\[11\] _06738_ _07498_ _07501_ VGND VGND VPWR VPWR
+ _07502_ sky130_fd_sc_hd__o211a_1
X_28854_ _12930_ VGND VGND VPWR VPWR _04213_ sky130_fd_sc_hd__clkbuf_1
X_21189_ _08471_ _08474_ VGND VGND VPWR VPWR _08475_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27805_ _12344_ VGND VGND VPWR VPWR _03750_ sky130_fd_sc_hd__clkbuf_1
X_28785_ _12764_ net2740 _12887_ VGND VGND VPWR VPWR _12894_ sky130_fd_sc_hd__mux2_1
X_25997_ net12 _11317_ VGND VGND VPWR VPWR _11323_ sky130_fd_sc_hd__or2_1
XFILLER_0_176_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27736_ _10838_ _10908_ _12260_ VGND VGND VPWR VPWR _12307_ sky130_fd_sc_hd__a21oi_4
X_15750_ _14139_ net2758 _14199_ VGND VGND VPWR VPWR _14204_ sky130_fd_sc_hd__mux2_1
X_24948_ _10450_ net3107 _10687_ VGND VGND VPWR VPWR _10693_ sky130_fd_sc_hd__mux2_1
Xhold1170 datamem.data_ram\[49\]\[13\] VGND VGND VPWR VPWR net2320 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14701_ net2487 _13260_ _13245_ VGND VGND VPWR VPWR _13261_ sky130_fd_sc_hd__mux2_1
Xhold1181 rvcpu.dp.rf.reg_file_arr\[9\]\[22\] VGND VGND VPWR VPWR net2331 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1192 datamem.data_ram\[62\]\[24\] VGND VGND VPWR VPWR net2342 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_310 _14160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15681_ _13222_ VGND VGND VPWR VPWR _14158_ sky130_fd_sc_hd__buf_4
X_27667_ _10570_ _10898_ _12260_ VGND VGND VPWR VPWR _12270_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_219_5750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24879_ _10476_ net2661 net92 VGND VGND VPWR VPWR _10656_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_219_5761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_321 _14434_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17420_ _04976_ VGND VGND VPWR VPWR _01330_ sky130_fd_sc_hd__clkbuf_1
X_29406_ clknet_leaf_0_clk _01141_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD2E\[17\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_332 _14457_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_343 _14474_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14632_ _13208_ VGND VGND VPWR VPWR _03195_ sky130_fd_sc_hd__clkbuf_1
X_26618_ _10824_ net3228 _11650_ VGND VGND VPWR VPWR _11657_ sky130_fd_sc_hd__mux2_1
XANTENNA_354 rvcpu.dp.SrcBFW_Mux.y\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_365 rvcpu.dp.plde.ImmExtE\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27598_ _10741_ _12106_ _12168_ VGND VGND VPWR VPWR _12233_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_157_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_215_5647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_376 rvcpu.dp.plmw.ReadDataW\[24\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_215_5658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_387 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_630 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17351_ _14133_ net2953 _04938_ VGND VGND VPWR VPWR _04940_ sky130_fd_sc_hd__mux2_1
X_23459__108 clknet_1_0__leaf__10157_ VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__inv_2
X_29337_ clknet_leaf_181_clk _01072_ VGND VGND VPWR VPWR datamem.data_ram\[62\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_26549_ _11064_ _11610_ VGND VGND VPWR VPWR _11619_ sky130_fd_sc_hd__and2_1
XANTENNA_398 _06600_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_222_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16302_ net3484 _14468_ _14511_ VGND VGND VPWR VPWR _14514_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_745 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_600 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17282_ _04903_ VGND VGND VPWR VPWR _01403_ sky130_fd_sc_hd__clkbuf_1
X_29268_ _09281_ net4148 _13150_ VGND VGND VPWR VPWR _13155_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19021_ _06352_ _06353_ VGND VGND VPWR VPWR _06354_ sky130_fd_sc_hd__and2_1
XFILLER_0_83_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_183_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28219_ _12578_ VGND VGND VPWR VPWR _03930_ sky130_fd_sc_hd__clkbuf_1
X_16233_ _13259_ VGND VGND VPWR VPWR _14474_ sky130_fd_sc_hd__buf_4
XFILLER_0_153_655 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29199_ _13117_ VGND VGND VPWR VPWR _04371_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload307 clknet_1_1__leaf__10196_ VGND VGND VPWR VPWR clkload307/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_36_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload15 clknet_5_17__leaf_clk VGND VGND VPWR VPWR clkload15/X sky130_fd_sc_hd__clkbuf_8
Xclkload318 clknet_1_1__leaf__10161_ VGND VGND VPWR VPWR clkload318/Y sky130_fd_sc_hd__clkinvlp_4
X_31230_ clknet_leaf_43_clk _02933_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCD\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload26 clknet_5_31__leaf_clk VGND VGND VPWR VPWR clkload26/Y sky130_fd_sc_hd__clkinv_8
Xclkload329 clknet_1_1__leaf__10265_ VGND VGND VPWR VPWR clkload329/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_180_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload37 clknet_leaf_25_clk VGND VGND VPWR VPWR clkload37/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_152_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16164_ _14427_ VGND VGND VPWR VPWR _01945_ sky130_fd_sc_hd__clkbuf_1
Xclkload48 clknet_leaf_44_clk VGND VGND VPWR VPWR clkload48/Y sky130_fd_sc_hd__clkinv_4
Xclkload59 clknet_leaf_6_clk VGND VGND VPWR VPWR clkload59/Y sky130_fd_sc_hd__inv_8
XFILLER_0_2_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15115_ _13657_ _13659_ _13353_ VGND VGND VPWR VPWR _13660_ sky130_fd_sc_hd__o21a_1
X_31161_ clknet_leaf_8_clk rvcpu.ALUResultE\[20\] VGND VGND VPWR VPWR rvcpu.dp.plem.ALUResultM\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_16095_ _14389_ VGND VGND VPWR VPWR _01976_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_71_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_192_Right_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15046_ _13297_ _13592_ VGND VGND VPWR VPWR _13593_ sky130_fd_sc_hd__and2_1
X_19923_ datamem.data_ram\[59\]\[17\] _06636_ _07214_ _07217_ VGND VGND VPWR VPWR
+ _07218_ sky130_fd_sc_hd__o211a_1
X_30112_ net474 _01847_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[10\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_31092_ clknet_leaf_101_clk _02827_ VGND VGND VPWR VPWR datamem.data_ram\[21\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_166_4477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_4488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24025__556 clknet_1_1__leaf__10243_ VGND VGND VPWR VPWR net682 sky130_fd_sc_hd__inv_2
XFILLER_0_208_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_216_clk clknet_5_21__leaf_clk VGND VGND VPWR VPWR clknet_leaf_216_clk
+ sky130_fd_sc_hd__clkbuf_8
X_30043_ net405 _01778_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[13\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_19854_ datamem.data_ram\[59\]\[1\] _06961_ _06948_ datamem.data_ram\[57\]\[1\] _07031_
+ VGND VGND VPWR VPWR _07149_ sky130_fd_sc_hd__a221o_1
XFILLER_0_208_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18805_ _05504_ _06151_ VGND VGND VPWR VPWR _06152_ sky130_fd_sc_hd__xnor2_1
X_19785_ datamem.data_ram\[45\]\[9\] _06703_ _06779_ datamem.data_ram\[40\]\[9\] _07079_
+ VGND VGND VPWR VPWR _07080_ sky130_fd_sc_hd__o221a_1
X_16997_ net2392 _14480_ _04742_ VGND VGND VPWR VPWR _04751_ sky130_fd_sc_hd__mux2_1
XFILLER_0_223_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18736_ _06085_ _06086_ VGND VGND VPWR VPWR _06087_ sky130_fd_sc_hd__or2_1
X_15948_ _13179_ _14271_ VGND VGND VPWR VPWR _14310_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_69_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31994_ clknet_leaf_127_clk _03416_ VGND VGND VPWR VPWR datamem.data_ram\[31\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_190_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_3484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_3495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30945_ clknet_leaf_100_clk _02680_ VGND VGND VPWR VPWR datamem.data_ram\[3\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_18667_ _05866_ _05696_ VGND VGND VPWR VPWR _06022_ sky130_fd_sc_hd__nand2_1
X_15879_ _14272_ VGND VGND VPWR VPWR _14273_ sky130_fd_sc_hd__buf_4
XFILLER_0_203_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17618_ _05080_ VGND VGND VPWR VPWR _01228_ sky130_fd_sc_hd__clkbuf_1
X_30876_ clknet_leaf_62_clk _02611_ VGND VGND VPWR VPWR datamem.data_ram\[42\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_18598_ _05589_ _05593_ _05356_ VGND VGND VPWR VPWR _05956_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_138_3801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32615_ clknet_leaf_81_clk _04037_ VGND VGND VPWR VPWR datamem.data_ram\[20\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17549_ _13278_ net2454 _05009_ VGND VGND VPWR VPWR _05044_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20560_ _06940_ VGND VGND VPWR VPWR _07851_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_134_3709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32546_ clknet_leaf_273_clk _03968_ VGND VGND VPWR VPWR datamem.data_ram\[23\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload9 clknet_5_10__leaf_clk VGND VGND VPWR VPWR clkload9/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_132_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19219_ _06526_ VGND VGND VPWR VPWR rvcpu.dp.lAuiPCE\[25\] sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_99_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20491_ _06589_ _07692_ _07782_ VGND VGND VPWR VPWR _07783_ sky130_fd_sc_hd__and3b_1
XFILLER_0_116_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32477_ clknet_leaf_253_clk _03899_ VGND VGND VPWR VPWR datamem.data_ram\[26\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_694 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22230_ rvcpu.dp.rf.reg_file_arr\[24\]\[0\] rvcpu.dp.rf.reg_file_arr\[25\]\[0\] rvcpu.dp.rf.reg_file_arr\[26\]\[0\]
+ rvcpu.dp.rf.reg_file_arr\[27\]\[0\] _09393_ _09395_ VGND VGND VPWR VPWR _09396_
+ sky130_fd_sc_hd__mux4_1
X_31428_ clknet_leaf_59_clk _03131_ VGND VGND VPWR VPWR datamem.data_ram\[44\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22161_ _09350_ VGND VGND VPWR VPWR _09351_ sky130_fd_sc_hd__buf_8
X_31359_ clknet_leaf_35_clk _03062_ VGND VGND VPWR VPWR rvcpu.dp.plde.ImmExtE\[8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_42_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__10207_ clknet_0__10207_ VGND VGND VPWR VPWR clknet_1_0__leaf__10207_
+ sky130_fd_sc_hd__clkbuf_16
X_21112_ datamem.data_ram\[29\]\[7\] _06639_ VGND VGND VPWR VPWR _08401_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22092_ rvcpu.dp.plem.WriteDataM\[25\] _09304_ _09215_ VGND VGND VPWR VPWR _09305_
+ sky130_fd_sc_hd__mux2_8
XTAP_TAPCELL_ROW_58_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__10138_ clknet_0__10138_ VGND VGND VPWR VPWR clknet_1_0__leaf__10138_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_58_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_207_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_207_clk
+ sky130_fd_sc_hd__clkbuf_8
X_25920_ rvcpu.dp.plfd.PCD\[16\] _11279_ VGND VGND VPWR VPWR _11280_ sky130_fd_sc_hd__or2_1
X_21043_ datamem.data_ram\[6\]\[31\] datamem.data_ram\[7\]\[31\] _07874_ VGND VGND
+ VPWR VPWR _08332_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_54_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_227_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25851_ _11206_ _11207_ _11232_ VGND VGND VPWR VPWR _11233_ sky130_fd_sc_hd__and3_1
XFILLER_0_226_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24802_ _10614_ VGND VGND VPWR VPWR _02477_ sky130_fd_sc_hd__clkbuf_1
X_28570_ _12779_ VGND VGND VPWR VPWR _04080_ sky130_fd_sc_hd__clkbuf_1
X_25782_ rvcpu.dp.pcreg.q\[12\] rvcpu.dp.pcreg.q\[11\] _11171_ VGND VGND VPWR VPWR
+ _11178_ sky130_fd_sc_hd__and3_1
X_27521_ _12192_ VGND VGND VPWR VPWR _03618_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24733_ _10575_ VGND VGND VPWR VPWR _02447_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21945_ _09169_ _09173_ _09177_ _08624_ VGND VGND VPWR VPWR _01057_ sky130_fd_sc_hd__o31a_1
XFILLER_0_222_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24664_ _10412_ net1523 _10531_ _10537_ VGND VGND VPWR VPWR _02416_ sky130_fd_sc_hd__a31o_1
XFILLER_0_167_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27452_ _12153_ net1994 _12143_ VGND VGND VPWR VPWR _12154_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21876_ rvcpu.dp.rf.reg_file_arr\[28\]\[26\] rvcpu.dp.rf.reg_file_arr\[30\]\[26\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[26\] rvcpu.dp.rf.reg_file_arr\[31\]\[26\] _08629_
+ _08683_ VGND VGND VPWR VPWR _09112_ sky130_fd_sc_hd__mux4_1
XFILLER_0_96_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26403_ rvcpu.dp.plde.JalrE VGND VGND VPWR VPWR _11545_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_77_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20827_ datamem.data_ram\[14\]\[30\] _07085_ _06618_ datamem.data_ram\[12\]\[30\]
+ VGND VGND VPWR VPWR _08117_ sky130_fd_sc_hd__o22a_1
X_24595_ _10498_ VGND VGND VPWR VPWR _02386_ sky130_fd_sc_hd__clkbuf_1
X_27383_ _10731_ net2426 net86 VGND VGND VPWR VPWR _12111_ sky130_fd_sc_hd__mux2_1
XFILLER_0_194_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29122_ _09223_ net3595 _13076_ VGND VGND VPWR VPWR _13077_ sky130_fd_sc_hd__mux2_1
X_26334_ _11501_ net1689 _11496_ _11502_ VGND VGND VPWR VPWR _03121_ sky130_fd_sc_hd__a31o_1
X_20758_ _08046_ _08047_ _07840_ VGND VGND VPWR VPWR _08048_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_210_5533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_210_5544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26265_ _11464_ VGND VGND VPWR VPWR _03090_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29053_ _10777_ _11020_ _12977_ VGND VGND VPWR VPWR _13040_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_108_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23477_ clknet_1_0__leaf__10152_ VGND VGND VPWR VPWR _10159_ sky130_fd_sc_hd__buf_1
X_23987__522 clknet_1_0__leaf__10239_ VGND VGND VPWR VPWR net648 sky130_fd_sc_hd__inv_2
X_20689_ datamem.data_ram\[48\]\[5\] _07122_ _07978_ _07979_ VGND VGND VPWR VPWR _07980_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_150_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28004_ _12463_ VGND VGND VPWR VPWR _03830_ sky130_fd_sc_hd__clkbuf_1
X_25216_ _10826_ net2332 net56 VGND VGND VPWR VPWR _10847_ sky130_fd_sc_hd__mux2_1
X_22428_ _09528_ _09587_ _09426_ VGND VGND VPWR VPWR _09588_ sky130_fd_sc_hd__a21o_1
XFILLER_0_162_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26196_ _11435_ VGND VGND VPWR VPWR _03050_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25147_ _10758_ net3703 _10802_ VGND VGND VPWR VPWR _10806_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22359_ _09390_ _09521_ VGND VGND VPWR VPWR _09522_ sky130_fd_sc_hd__or2_1
XFILLER_0_209_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25078_ _10770_ VGND VGND VPWR VPWR _02597_ sky130_fd_sc_hd__clkbuf_1
X_29955_ net325 _01690_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[15\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_208_5484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_208_5495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16920_ _04710_ VGND VGND VPWR VPWR _01580_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28906_ _12749_ net2745 net68 VGND VGND VPWR VPWR _12958_ sky130_fd_sc_hd__mux2_1
X_29886_ net264 _01621_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[17\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28837_ _12921_ VGND VGND VPWR VPWR _04205_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_161_4352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16851_ net3046 _14470_ _04670_ VGND VGND VPWR VPWR _04674_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_161_4363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15802_ _14191_ net3848 _14221_ VGND VGND VPWR VPWR _14231_ sky130_fd_sc_hd__mux2_1
XFILLER_0_176_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19570_ datamem.data_ram\[5\]\[8\] _06865_ _06672_ datamem.data_ram\[7\]\[8\] VGND
+ VGND VPWR VPWR _06866_ sky130_fd_sc_hd__o22a_1
X_16782_ _04637_ VGND VGND VPWR VPWR _01653_ sky130_fd_sc_hd__clkbuf_1
X_28768_ _12884_ VGND VGND VPWR VPWR _04173_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_217_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18521_ _05879_ _05864_ _05880_ _05881_ VGND VGND VPWR VPWR _05882_ sky130_fd_sc_hd__a211o_1
X_15733_ _13274_ VGND VGND VPWR VPWR _14193_ sky130_fd_sc_hd__buf_4
X_27719_ _10838_ _10898_ _12260_ VGND VGND VPWR VPWR _12298_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_217_5709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28699_ _12747_ net2230 net42 VGND VGND VPWR VPWR _12848_ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18452_ _05810_ _05786_ _05813_ _05814_ VGND VGND VPWR VPWR _05815_ sky130_fd_sc_hd__a2bb2o_1
X_30730_ clknet_leaf_221_clk _02465_ VGND VGND VPWR VPWR datamem.data_ram\[48\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_64_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15664_ _14146_ VGND VGND VPWR VPWR _02180_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_140 _07833_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_151 _07874_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17403_ _14185_ net3155 _04960_ VGND VGND VPWR VPWR _04967_ sky130_fd_sc_hd__mux2_1
XANTENNA_162 _08568_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14615_ net2016 _13195_ _13181_ VGND VGND VPWR VPWR _13196_ sky130_fd_sc_hd__mux2_1
XANTENNA_173 _08744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18383_ _05743_ _05744_ _05746_ VGND VGND VPWR VPWR _05747_ sky130_fd_sc_hd__a21oi_1
X_30661_ clknet_leaf_149_clk _02396_ VGND VGND VPWR VPWR datamem.data_ram\[50\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_184 _09059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15595_ _14105_ VGND VGND VPWR VPWR _02208_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_195 _09321_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32400_ clknet_leaf_4_clk _03822_ VGND VGND VPWR VPWR datamem.data_ram\[29\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_17334_ _04930_ VGND VGND VPWR VPWR _01378_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30592_ clknet_leaf_117_clk _02327_ VGND VGND VPWR VPWR datamem.data_ram\[53\]\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_102_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32331_ clknet_leaf_249_clk _03753_ VGND VGND VPWR VPWR datamem.data_ram\[31\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_17265_ _04893_ VGND VGND VPWR VPWR _01410_ sky130_fd_sc_hd__clkbuf_1
Xclkload104 clknet_leaf_90_clk VGND VGND VPWR VPWR clkload104/Y sky130_fd_sc_hd__clkinvlp_2
X_19004_ _06335_ _06336_ _05240_ VGND VGND VPWR VPWR _06338_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_12_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16216_ _14462_ VGND VGND VPWR VPWR _01928_ sky130_fd_sc_hd__clkbuf_1
Xclkload115 clknet_leaf_94_clk VGND VGND VPWR VPWR clkload115/Y sky130_fd_sc_hd__inv_6
XFILLER_0_141_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32262_ clknet_leaf_272_clk _03684_ VGND VGND VPWR VPWR datamem.data_ram\[34\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_168_4517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17196_ _14183_ net3131 _04851_ VGND VGND VPWR VPWR _04857_ sky130_fd_sc_hd__mux2_1
Xclkload126 clknet_leaf_253_clk VGND VGND VPWR VPWR clkload126/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_168_4528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload137 clknet_leaf_242_clk VGND VGND VPWR VPWR clkload137/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_70_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_180_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_168_4539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload148 clknet_leaf_261_clk VGND VGND VPWR VPWR clkload148/Y sky130_fd_sc_hd__clkinvlp_4
X_31213_ clknet_leaf_32_clk _02916_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCD\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_94_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload159 clknet_leaf_174_clk VGND VGND VPWR VPWR clkload159/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_0_24_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16147_ _14416_ VGND VGND VPWR VPWR _01951_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32193_ clknet_leaf_226_clk _03615_ VGND VGND VPWR VPWR datamem.data_ram\[36\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_23356__993 clknet_1_0__leaf__10137_ VGND VGND VPWR VPWR net1119 sky130_fd_sc_hd__inv_2
XFILLER_0_84_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31144_ clknet_leaf_63_clk rvcpu.ALUResultE\[3\] VGND VGND VPWR VPWR rvcpu.dp.plem.ALUResultM\[3\]
+ sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_90_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16078_ net2229 _13269_ _14371_ VGND VGND VPWR VPWR _14380_ sky130_fd_sc_hd__mux2_1
XFILLER_0_220_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_227_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15029_ _13553_ _13575_ VGND VGND VPWR VPWR _13576_ sky130_fd_sc_hd__and2b_1
X_19906_ datamem.data_ram\[12\]\[17\] _07182_ _07197_ _07200_ VGND VGND VPWR VPWR
+ _07201_ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31075_ clknet_leaf_157_clk _02810_ VGND VGND VPWR VPWR datamem.data_ram\[9\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2607 rvcpu.dp.rf.reg_file_arr\[13\]\[25\] VGND VGND VPWR VPWR net3757 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2618 datamem.data_ram\[27\]\[22\] VGND VGND VPWR VPWR net3768 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_127_3535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2629 datamem.data_ram\[14\]\[28\] VGND VGND VPWR VPWR net3779 sky130_fd_sc_hd__dlygate4sd3_1
X_19837_ _06921_ VGND VGND VPWR VPWR _07132_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_127_3546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30026_ net388 _01761_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[13\]\[13\] sky130_fd_sc_hd__dfxtp_1
Xhold1906 datamem.data_ram\[27\]\[15\] VGND VGND VPWR VPWR net3056 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1917 datamem.data_ram\[19\]\[29\] VGND VGND VPWR VPWR net3067 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1928 datamem.data_ram\[25\]\[29\] VGND VGND VPWR VPWR net3078 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1939 datamem.data_ram\[1\]\[25\] VGND VGND VPWR VPWR net3089 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19768_ datamem.data_ram\[30\]\[25\] _06763_ _06691_ datamem.data_ram\[26\]\[25\]
+ VGND VGND VPWR VPWR _07063_ sky130_fd_sc_hd__o22a_1
X_18719_ _05776_ _05922_ _05926_ _05858_ VGND VGND VPWR VPWR _06071_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_88_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19699_ datamem.data_ram\[13\]\[0\] _06921_ _06993_ datamem.data_ram\[15\]\[0\] _06994_
+ VGND VGND VPWR VPWR _06995_ sky130_fd_sc_hd__a221o_1
X_31977_ clknet_leaf_150_clk _03399_ VGND VGND VPWR VPWR datamem.data_ram\[53\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23856__419 clknet_1_1__leaf__10219_ VGND VGND VPWR VPWR net545 sky130_fd_sc_hd__inv_2
X_21730_ rvcpu.dp.rf.reg_file_arr\[24\]\[18\] rvcpu.dp.rf.reg_file_arr\[25\]\[18\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[18\] rvcpu.dp.rf.reg_file_arr\[27\]\[18\] _08536_
+ _08693_ VGND VGND VPWR VPWR _08974_ sky130_fd_sc_hd__mux4_1
X_30928_ clknet_leaf_155_clk _02663_ VGND VGND VPWR VPWR datamem.data_ram\[40\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21661_ rvcpu.dp.rf.reg_file_arr\[4\]\[14\] rvcpu.dp.rf.reg_file_arr\[5\]\[14\] rvcpu.dp.rf.reg_file_arr\[6\]\[14\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[14\] _08687_ _08856_ VGND VGND VPWR VPWR _08909_
+ sky130_fd_sc_hd__mux4_1
X_30859_ clknet_leaf_156_clk _02594_ VGND VGND VPWR VPWR datamem.data_ram\[43\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23400_ _09330_ net2981 _10143_ VGND VGND VPWR VPWR _10151_ sky130_fd_sc_hd__mux2_1
X_20612_ _05347_ _06594_ VGND VGND VPWR VPWR _07903_ sky130_fd_sc_hd__nand2_8
XFILLER_0_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24380_ _09236_ net4359 _10367_ VGND VGND VPWR VPWR _10369_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21592_ _08842_ _08843_ VGND VGND VPWR VPWR _08844_ sky130_fd_sc_hd__or2_1
XFILLER_0_188_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20543_ datamem.data_ram\[5\]\[21\] _07833_ VGND VGND VPWR VPWR _07834_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32529_ clknet_leaf_245_clk _03951_ VGND VGND VPWR VPWR datamem.data_ram\[23\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_26050_ _11081_ _11351_ VGND VGND VPWR VPWR _11354_ sky130_fd_sc_hd__and2_1
XFILLER_0_7_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20474_ datamem.data_ram\[34\]\[20\] _06690_ _06633_ datamem.data_ram\[35\]\[20\]
+ _06678_ VGND VGND VPWR VPWR _07766_ sky130_fd_sc_hd__o221a_1
XFILLER_0_15_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25001_ _10721_ VGND VGND VPWR VPWR _02569_ sky130_fd_sc_hd__clkbuf_1
X_22213_ _09379_ VGND VGND VPWR VPWR _01123_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_160_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23193_ _10117_ VGND VGND VPWR VPWR _01365_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Left_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22144_ _09267_ net3441 net62 VGND VGND VPWR VPWR _09342_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29740_ net1086 _01475_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[21\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_26952_ _11829_ _11854_ VGND VGND VPWR VPWR _11858_ sky130_fd_sc_hd__and2_1
X_22075_ rvcpu.dp.plem.WriteDataM\[7\] _09264_ _09265_ rvcpu.dp.plem.WriteDataM\[15\]
+ VGND VGND VPWR VPWR _09290_ sky130_fd_sc_hd__a22o_4
XFILLER_0_227_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25903_ _13539_ _11268_ VGND VGND VPWR VPWR _11270_ sky130_fd_sc_hd__nand2_1
X_21026_ _06917_ _08314_ VGND VGND VPWR VPWR _08315_ sky130_fd_sc_hd__or2_1
X_29671_ net1017 _01406_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[23\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_26883_ _11681_ _11810_ VGND VGND VPWR VPWR _11814_ sky130_fd_sc_hd__and2_1
X_23568__191 clknet_1_0__leaf__10175_ VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_203_5370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28622_ _12807_ VGND VGND VPWR VPWR _04104_ sky130_fd_sc_hd__clkbuf_1
X_25834_ rvcpu.dp.plfd.PCPlus4D\[23\] _11218_ _11142_ VGND VGND VPWR VPWR _11219_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_199_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28553_ _12770_ VGND VGND VPWR VPWR _04072_ sky130_fd_sc_hd__clkbuf_1
X_25765_ _13514_ _13876_ VGND VGND VPWR VPWR _11165_ sky130_fd_sc_hd__nand2_1
X_22977_ clknet_1_0__leaf__10080_ VGND VGND VPWR VPWR _10083_ sky130_fd_sc_hd__buf_1
XFILLER_0_214_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_195_5171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_198_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_195_5182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_27_Left_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27504_ _12183_ VGND VGND VPWR VPWR _03610_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24716_ _10474_ net4220 net59 VGND VGND VPWR VPWR _10566_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28484_ _11968_ _12724_ VGND VGND VPWR VPWR _12726_ sky130_fd_sc_hd__and2_1
XFILLER_0_179_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21928_ rvcpu.dp.rf.reg_file_arr\[16\]\[29\] rvcpu.dp.rf.reg_file_arr\[17\]\[29\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[29\] rvcpu.dp.rf.reg_file_arr\[19\]\[29\] _08631_
+ _08632_ VGND VGND VPWR VPWR _09161_ sky130_fd_sc_hd__mux4_1
XFILLER_0_70_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25696_ _11091_ _11113_ VGND VGND VPWR VPWR _11120_ sky130_fd_sc_hd__and2_1
XFILLER_0_214_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_191_5068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_191_5079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27435_ _09266_ VGND VGND VPWR VPWR _12142_ sky130_fd_sc_hd__buf_2
XFILLER_0_155_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24647_ _10527_ VGND VGND VPWR VPWR _02409_ sky130_fd_sc_hd__clkbuf_1
X_21859_ _08515_ _09095_ VGND VGND VPWR VPWR _09096_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24054__582 clknet_1_0__leaf__10246_ VGND VGND VPWR VPWR net708 sky130_fd_sc_hd__inv_2
XFILLER_0_195_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15380_ _13432_ _13773_ _13441_ VGND VGND VPWR VPWR _13914_ sky130_fd_sc_hd__or3_1
XFILLER_0_37_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27366_ _12101_ VGND VGND VPWR VPWR _03554_ sky130_fd_sc_hd__clkbuf_1
X_24578_ _10489_ VGND VGND VPWR VPWR _02378_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_5_19__f_clk clknet_2_2_0_clk VGND VGND VPWR VPWR clknet_5_19__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_167_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29105_ _09266_ net3158 _13067_ VGND VGND VPWR VPWR _13068_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_203_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26317_ _11491_ VGND VGND VPWR VPWR _03115_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27297_ _11978_ _12054_ VGND VGND VPWR VPWR _12062_ sky130_fd_sc_hd__and2_1
XFILLER_0_151_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29036_ _10932_ _10778_ VGND VGND VPWR VPWR _13031_ sky130_fd_sc_hd__nor2_1
X_17050_ net4090 _14463_ _04779_ VGND VGND VPWR VPWR _04780_ sky130_fd_sc_hd__mux2_1
X_26248_ _11438_ _11458_ _11459_ net2479 VGND VGND VPWR VPWR _03078_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_150_4086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_4097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16001_ _14338_ VGND VGND VPWR VPWR _02027_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_36_Left_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26179_ _11426_ VGND VGND VPWR VPWR _03042_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_4403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_4414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17952_ _05320_ _05323_ VGND VGND VPWR VPWR _05324_ sky130_fd_sc_hd__nor2_1
X_29938_ net308 _01673_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[16\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_26515__3 clknet_1_1__leaf__10080_ VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__inv_2
X_16903_ _04701_ VGND VGND VPWR VPWR _01588_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_224_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17883_ rvcpu.dp.plde.Rs1E\[1\] rvcpu.dp.plmw.RdW\[1\] VGND VGND VPWR VPWR _05256_
+ sky130_fd_sc_hd__xor2_1
X_29869_ net247 _01604_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[17\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31900_ _04442_ net121 VGND VGND VPWR VPWR datamem.rd_data_mem\[5\] sky130_fd_sc_hd__dlxtn_1
X_19622_ _06605_ _06917_ VGND VGND VPWR VPWR _06918_ sky130_fd_sc_hd__nor2_1
X_16834_ net1876 _14453_ _04659_ VGND VGND VPWR VPWR _04665_ sky130_fd_sc_hd__mux2_1
X_32880_ clknet_leaf_57_clk _04302_ VGND VGND VPWR VPWR datamem.data_ram\[10\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_122_3421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_45_Left_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_221_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_178_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_3432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19553_ datamem.data_ram\[14\]\[24\] _06625_ _06689_ datamem.data_ram\[10\]\[24\]
+ VGND VGND VPWR VPWR _06849_ sky130_fd_sc_hd__o22a_1
X_31831_ clknet_leaf_235_clk _03285_ VGND VGND VPWR VPWR datamem.data_ram\[3\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_16765_ _04628_ VGND VGND VPWR VPWR _01661_ sky130_fd_sc_hd__clkbuf_1
X_18504_ _05590_ VGND VGND VPWR VPWR _05866_ sky130_fd_sc_hd__buf_2
X_15716_ _14181_ net2468 _14173_ VGND VGND VPWR VPWR _14182_ sky130_fd_sc_hd__mux2_1
X_31762_ clknet_leaf_107_clk _03216_ VGND VGND VPWR VPWR datamem.data_ram\[18\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_19484_ _06654_ VGND VGND VPWR VPWR _06780_ sky130_fd_sc_hd__buf_8
X_16696_ _14160_ net2911 _04587_ VGND VGND VPWR VPWR _04592_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18435_ _05797_ VGND VGND VPWR VPWR _05798_ sky130_fd_sc_hd__inv_2
X_30713_ clknet_leaf_147_clk _02448_ VGND VGND VPWR VPWR datamem.data_ram\[49\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_83_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15647_ _13186_ VGND VGND VPWR VPWR _14135_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_83_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31693_ clknet_leaf_39_clk _03151_ VGND VGND VPWR VPWR rvcpu.dp.pcreg.q\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30644_ clknet_leaf_139_clk _02379_ VGND VGND VPWR VPWR datamem.data_ram\[51\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_18366_ _05236_ rvcpu.dp.plde.ALUControlE\[0\] rvcpu.dp.plde.ALUControlE\[1\] VGND
+ VGND VPWR VPWR _05731_ sky130_fd_sc_hd__or3b_1
XFILLER_0_173_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15578_ _14096_ VGND VGND VPWR VPWR _02216_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17317_ _04921_ VGND VGND VPWR VPWR _01386_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_96_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18297_ _05576_ VGND VGND VPWR VPWR _05662_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_44_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30575_ clknet_leaf_182_clk _02310_ VGND VGND VPWR VPWR datamem.data_ram\[54\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_54_Left_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32314_ clknet_leaf_213_clk _03736_ VGND VGND VPWR VPWR datamem.data_ram\[31\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17248_ _04884_ VGND VGND VPWR VPWR _01418_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_189_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_181_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32245_ clknet_leaf_224_clk _03667_ VGND VGND VPWR VPWR datamem.data_ram\[34\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_17179_ _14166_ net4367 _04840_ VGND VGND VPWR VPWR _04848_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20190_ datamem.data_ram\[40\]\[11\] _06697_ _07024_ datamem.data_ram\[44\]\[11\]
+ VGND VGND VPWR VPWR _07483_ sky130_fd_sc_hd__o22a_1
X_32176_ clknet_leaf_200_clk _03598_ VGND VGND VPWR VPWR datamem.data_ram\[37\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3105 datamem.data_ram\[28\]\[24\] VGND VGND VPWR VPWR net4255 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3116 datamem.data_ram\[61\]\[17\] VGND VGND VPWR VPWR net4266 sky130_fd_sc_hd__dlygate4sd3_1
X_31127_ clknet_leaf_125_clk _02862_ VGND VGND VPWR VPWR datamem.data_ram\[25\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3127 rvcpu.dp.rf.reg_file_arr\[21\]\[17\] VGND VGND VPWR VPWR net4277 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3138 rvcpu.dp.rf.reg_file_arr\[22\]\[19\] VGND VGND VPWR VPWR net4288 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2404 datamem.data_ram\[57\]\[19\] VGND VGND VPWR VPWR net3554 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3149 rvcpu.dp.rf.reg_file_arr\[27\]\[23\] VGND VGND VPWR VPWR net4299 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2415 datamem.data_ram\[49\]\[9\] VGND VGND VPWR VPWR net3565 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2426 datamem.data_ram\[20\]\[11\] VGND VGND VPWR VPWR net3576 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31058_ clknet_leaf_93_clk _02793_ VGND VGND VPWR VPWR datamem.data_ram\[38\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2437 datamem.data_ram\[36\]\[8\] VGND VGND VPWR VPWR net3587 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1703 datamem.data_ram\[0\]\[18\] VGND VGND VPWR VPWR net2853 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2448 rvcpu.dp.rf.reg_file_arr\[25\]\[31\] VGND VGND VPWR VPWR net3598 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2459 datamem.data_ram\[47\]\[30\] VGND VGND VPWR VPWR net3609 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1714 datamem.data_ram\[47\]\[26\] VGND VGND VPWR VPWR net2864 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_3988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1725 rvcpu.dp.rf.reg_file_arr\[21\]\[30\] VGND VGND VPWR VPWR net2875 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_3999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_63_Left_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22900_ _09429_ _10032_ _10034_ VGND VGND VPWR VPWR _10035_ sky130_fd_sc_hd__a21o_1
X_30009_ clknet_leaf_181_clk _01744_ VGND VGND VPWR VPWR datamem.data_ram\[59\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1736 rvcpu.dp.rf.reg_file_arr\[22\]\[26\] VGND VGND VPWR VPWR net2886 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1747 datamem.data_ram\[19\]\[11\] VGND VGND VPWR VPWR net2897 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1758 rvcpu.dp.rf.reg_file_arr\[31\]\[23\] VGND VGND VPWR VPWR net2908 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1769 rvcpu.dp.rf.reg_file_arr\[15\]\[15\] VGND VGND VPWR VPWR net2919 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22831_ _09969_ VGND VGND VPWR VPWR _01151_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_194_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25550_ _11033_ VGND VGND VPWR VPWR _02806_ sky130_fd_sc_hd__clkbuf_1
X_22762_ rvcpu.dp.rf.reg_file_arr\[28\]\[24\] rvcpu.dp.rf.reg_file_arr\[30\]\[24\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[24\] rvcpu.dp.rf.reg_file_arr\[31\]\[24\] _09446_
+ _09402_ VGND VGND VPWR VPWR _09904_ sky130_fd_sc_hd__mux4_1
XFILLER_0_154_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24501_ _09235_ VGND VGND VPWR VPWR _10442_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_49_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26495__48 clknet_1_1__leaf__11601_ VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__inv_2
X_21713_ _08686_ _08957_ _08748_ VGND VGND VPWR VPWR _08958_ sky130_fd_sc_hd__o21ai_1
X_25481_ _10061_ net35 _10996_ net1334 VGND VGND VPWR VPWR _02774_ sky130_fd_sc_hd__a22o_1
XFILLER_0_177_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_566 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22693_ _09516_ _09836_ _09838_ _09523_ VGND VGND VPWR VPWR _09839_ sky130_fd_sc_hd__o211a_1
XFILLER_0_13_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27220_ _12005_ net1578 _12018_ _12021_ VGND VGND VPWR VPWR _03488_ sky130_fd_sc_hd__a31o_1
XFILLER_0_176_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24432_ _10399_ VGND VGND VPWR VPWR _02322_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21644_ _08813_ _08892_ _08689_ VGND VGND VPWR VPWR _08893_ sky130_fd_sc_hd__a21o_1
XFILLER_0_192_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_536 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27151_ _11974_ net1694 _11964_ _11979_ VGND VGND VPWR VPWR _03461_ sky130_fd_sc_hd__a31o_1
XFILLER_0_164_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24363_ _10359_ VGND VGND VPWR VPWR _02293_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_40 _06677_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21575_ _08824_ _08826_ _08743_ VGND VGND VPWR VPWR _08827_ sky130_fd_sc_hd__mux2_2
XFILLER_0_62_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_51 _06686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26102_ _11371_ VGND VGND VPWR VPWR _11386_ sky130_fd_sc_hd__buf_2
XFILLER_0_117_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23314_ clknet_1_0__leaf__10130_ VGND VGND VPWR VPWR _10134_ sky130_fd_sc_hd__buf_1
XANTENNA_62 _06742_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_73 _06776_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27082_ _11526_ _11934_ VGND VGND VPWR VPWR _11935_ sky130_fd_sc_hd__or2_1
XFILLER_0_191_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20526_ datamem.data_ram\[21\]\[21\] _07019_ _07815_ _07816_ VGND VGND VPWR VPWR
+ _07817_ sky130_fd_sc_hd__o211a_1
XANTENNA_84 _06784_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24294_ _10320_ VGND VGND VPWR VPWR _02263_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_95 _06810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26033_ _11121_ net1739 _11339_ _11343_ VGND VGND VPWR VPWR _02979_ sky130_fd_sc_hd__a31o_1
XFILLER_0_31_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20457_ datamem.data_ram\[24\]\[20\] _06821_ _06781_ datamem.data_ram\[25\]\[20\]
+ VGND VGND VPWR VPWR _07749_ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20388_ datamem.data_ram\[22\]\[28\] _06744_ _07243_ datamem.data_ram\[17\]\[28\]
+ VGND VGND VPWR VPWR _07680_ sky130_fd_sc_hd__o22a_1
XFILLER_0_24_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_205_5410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_205_5421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22127_ _09224_ net4043 _09332_ VGND VGND VPWR VPWR _09333_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_330 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27984_ _09272_ VGND VGND VPWR VPWR _12450_ sky130_fd_sc_hd__clkbuf_2
X_29723_ net1069 _01458_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[22\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26935_ _11831_ net1549 _11841_ _11847_ VGND VGND VPWR VPWR _03377_ sky130_fd_sc_hd__a31o_1
X_22058_ _09277_ VGND VGND VPWR VPWR _01070_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_201_5318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_201_5329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23724__316 clknet_1_0__leaf__10198_ VGND VGND VPWR VPWR net442 sky130_fd_sc_hd__inv_2
XFILLER_0_215_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_197_5222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_197_5233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21009_ _07872_ _08254_ _08269_ _08297_ VGND VGND VPWR VPWR _08298_ sky130_fd_sc_hd__o211a_2
Xhold2960 rvcpu.dp.rf.reg_file_arr\[10\]\[26\] VGND VGND VPWR VPWR net4110 sky130_fd_sc_hd__dlygate4sd3_1
X_29654_ net1000 _01389_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[24\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_14880_ rvcpu.dp.pcreg.q\[3\] _13280_ VGND VGND VPWR VPWR _13432_ sky130_fd_sc_hd__nor2b_4
XFILLER_0_214_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26866_ _10066_ VGND VGND VPWR VPWR _11803_ sky130_fd_sc_hd__clkbuf_4
Xhold2971 datamem.data_ram\[25\]\[21\] VGND VGND VPWR VPWR net4121 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2982 rvcpu.dp.rf.reg_file_arr\[11\]\[12\] VGND VGND VPWR VPWR net4132 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2993 datamem.data_ram\[51\]\[21\] VGND VGND VPWR VPWR net4143 sky130_fd_sc_hd__dlygate4sd3_1
X_28605_ _12798_ VGND VGND VPWR VPWR _04096_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_193_5119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25817_ _11203_ _11204_ _11157_ VGND VGND VPWR VPWR _11205_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_3_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29585_ net939 _01320_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[26\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_26797_ _10297_ _08066_ _11609_ VGND VGND VPWR VPWR _11762_ sky130_fd_sc_hd__and3_2
XFILLER_0_173_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28536_ _12759_ VGND VGND VPWR VPWR _04066_ sky130_fd_sc_hd__clkbuf_1
X_16550_ _04502_ VGND VGND VPWR VPWR _04514_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_74_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25748_ _11151_ VGND VGND VPWR VPWR _11152_ sky130_fd_sc_hd__buf_2
Xmax_cap64 _13094_ VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__buf_4
Xmax_cap75 _12510_ VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__buf_4
XFILLER_0_98_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15501_ _13398_ _13488_ _13402_ _14009_ VGND VGND VPWR VPWR _14029_ sky130_fd_sc_hd__o31a_1
Xmax_cap86 _12107_ VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__buf_4
Xmax_cap97 _12464_ VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__buf_4
XFILLER_0_167_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_4240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28467_ _12452_ net2747 _12713_ VGND VGND VPWR VPWR _12716_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16481_ _04477_ VGND VGND VPWR VPWR _01802_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25679_ _08125_ VGND VGND VPWR VPWR _11109_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_156_4251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18220_ _05582_ _05583_ _05584_ VGND VGND VPWR VPWR _05585_ sky130_fd_sc_hd__o21ai_1
X_15432_ _13506_ _13398_ _13703_ VGND VGND VPWR VPWR _13963_ sky130_fd_sc_hd__or3b_1
XFILLER_0_167_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27418_ _12130_ net2538 _12126_ VGND VGND VPWR VPWR _12131_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_171 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28398_ _12675_ VGND VGND VPWR VPWR _04012_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_152_4137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_4148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18151_ _05503_ _05515_ VGND VGND VPWR VPWR _05516_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15363_ _13528_ _13512_ _13514_ VGND VGND VPWR VPWR _13898_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_26_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27349_ _09321_ VGND VGND VPWR VPWR _12091_ sky130_fd_sc_hd__buf_2
XFILLER_0_93_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23770__358 clknet_1_0__leaf__10202_ VGND VGND VPWR VPWR net484 sky130_fd_sc_hd__inv_2
X_17102_ _04807_ VGND VGND VPWR VPWR _01487_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18082_ _05447_ _05448_ _05449_ VGND VGND VPWR VPWR _05450_ sky130_fd_sc_hd__o21ai_1
X_30360_ net706 _02095_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[3\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_15294_ _13298_ _13488_ _13447_ VGND VGND VPWR VPWR _13832_ sky130_fd_sc_hd__or3_1
XFILLER_0_41_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17033_ net2227 _14447_ _04768_ VGND VGND VPWR VPWR _04771_ sky130_fd_sc_hd__mux2_1
X_29019_ _13021_ VGND VGND VPWR VPWR _04287_ sky130_fd_sc_hd__clkbuf_1
X_30291_ net637 _02026_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[5\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23885__445 clknet_1_1__leaf__10222_ VGND VGND VPWR VPWR net571 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_229_5988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32030_ clknet_leaf_128_clk _03452_ VGND VGND VPWR VPWR datamem.data_ram\[26\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_111_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_229_5999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_186_4970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_111_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_221_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24104__612 clknet_1_0__leaf__10258_ VGND VGND VPWR VPWR net738 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_182_4856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18984_ _05886_ _06307_ _06309_ _06319_ VGND VGND VPWR VPWR rvcpu.ALUResultE\[28\]
+ sky130_fd_sc_hd__o211ai_4
XTAP_TAPCELL_ROW_182_4867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17935_ _13234_ rvcpu.dp.plde.RD2E\[14\] _05194_ VGND VGND VPWR VPWR _05308_ sky130_fd_sc_hd__mux2_1
XFILLER_0_225_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23664__263 clknet_1_0__leaf__10191_ VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__inv_2
XFILLER_0_79_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32932_ clknet_leaf_153_clk _04354_ VGND VGND VPWR VPWR datamem.data_ram\[7\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_17866_ _05238_ VGND VGND VPWR VPWR _05239_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_1_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19605_ datamem.data_ram\[22\]\[8\] _06682_ _06790_ datamem.data_ram\[17\]\[8\] _06900_
+ VGND VGND VPWR VPWR _06901_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_1_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16817_ net2244 _14436_ _04648_ VGND VGND VPWR VPWR _04656_ sky130_fd_sc_hd__mux2_1
X_32863_ clknet_leaf_55_clk _04285_ VGND VGND VPWR VPWR datamem.data_ram\[11\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_85_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17797_ _05179_ _05180_ rvcpu.dp.plde.RD2E\[4\] VGND VGND VPWR VPWR _05191_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_85_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_141_3874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31814_ clknet_leaf_106_clk _03268_ VGND VGND VPWR VPWR datamem.data_ram\[17\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_141_3885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19536_ datamem.data_ram\[32\]\[24\] _06811_ _06655_ datamem.data_ram\[33\]\[24\]
+ _06831_ VGND VGND VPWR VPWR _06832_ sky130_fd_sc_hd__o221a_1
XFILLER_0_152_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16748_ _04619_ VGND VGND VPWR VPWR _01669_ sky130_fd_sc_hd__clkbuf_1
X_32794_ clknet_leaf_212_clk _04216_ VGND VGND VPWR VPWR datamem.data_ram\[13\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19467_ _06744_ VGND VGND VPWR VPWR _06763_ sky130_fd_sc_hd__buf_6
X_31745_ net130 _03203_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[9\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16679_ _14143_ net2729 _04576_ VGND VGND VPWR VPWR _04583_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18418_ _05749_ _05781_ VGND VGND VPWR VPWR _05782_ sky130_fd_sc_hd__nand2_2
XFILLER_0_115_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24150__654 clknet_1_1__leaf__10262_ VGND VGND VPWR VPWR net780 sky130_fd_sc_hd__inv_2
XFILLER_0_173_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31676_ clknet_leaf_8_clk net1272 VGND VGND VPWR VPWR rvcpu.dp.plmw.ALUResultW\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_19398_ datamem.data_ram\[6\]\[16\] _06683_ _06688_ datamem.data_ram\[4\]\[16\] _06693_
+ VGND VGND VPWR VPWR _06694_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_44_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18349_ _05527_ _05533_ _05665_ VGND VGND VPWR VPWR _05714_ sky130_fd_sc_hd__mux2_1
X_30627_ clknet_leaf_177_clk _02362_ VGND VGND VPWR VPWR datamem.data_ram\[52\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_100_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21360_ _08598_ _08620_ _08621_ VGND VGND VPWR VPWR _08622_ sky130_fd_sc_hd__and3_4
XFILLER_0_127_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30558_ clknet_leaf_218_clk _02293_ VGND VGND VPWR VPWR datamem.data_ram\[54\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_20311_ datamem.data_ram\[0\]\[4\] _07138_ _07601_ _07602_ _07081_ VGND VGND VPWR
+ VPWR _07603_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_140_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold800 rvcpu.dp.rf.reg_file_arr\[7\]\[21\] VGND VGND VPWR VPWR net1950 sky130_fd_sc_hd__dlygate4sd3_1
X_21291_ _08552_ VGND VGND VPWR VPWR _08553_ sky130_fd_sc_hd__buf_4
Xhold811 rvcpu.dp.rf.reg_file_arr\[20\]\[3\] VGND VGND VPWR VPWR net1961 sky130_fd_sc_hd__dlygate4sd3_1
X_30489_ clknet_leaf_204_clk _02224_ VGND VGND VPWR VPWR datamem.data_ram\[57\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold822 rvcpu.dp.rf.reg_file_arr\[2\]\[10\] VGND VGND VPWR VPWR net1972 sky130_fd_sc_hd__dlygate4sd3_1
X_20242_ datamem.data_ram\[62\]\[3\] _07127_ _06976_ datamem.data_ram\[60\]\[3\] VGND
+ VGND VPWR VPWR _07535_ sky130_fd_sc_hd__a22o_1
X_32228_ clknet_leaf_169_clk _03650_ VGND VGND VPWR VPWR datamem.data_ram\[35\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold833 rvcpu.dp.rf.reg_file_arr\[11\]\[6\] VGND VGND VPWR VPWR net1983 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold844 datamem.data_ram\[38\]\[13\] VGND VGND VPWR VPWR net1994 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold855 rvcpu.dp.rf.reg_file_arr\[3\]\[28\] VGND VGND VPWR VPWR net2005 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold866 rvcpu.dp.rf.reg_file_arr\[9\]\[27\] VGND VGND VPWR VPWR net2016 sky130_fd_sc_hd__dlygate4sd3_1
Xhold877 rvcpu.dp.rf.reg_file_arr\[6\]\[4\] VGND VGND VPWR VPWR net2027 sky130_fd_sc_hd__dlygate4sd3_1
X_32159_ clknet_leaf_89_clk _03581_ VGND VGND VPWR VPWR datamem.data_ram\[38\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold888 datamem.data_ram\[14\]\[23\] VGND VGND VPWR VPWR net2038 sky130_fd_sc_hd__dlygate4sd3_1
X_20173_ datamem.data_ram\[19\]\[11\] _06731_ _06656_ datamem.data_ram\[17\]\[11\]
+ VGND VGND VPWR VPWR _07466_ sky130_fd_sc_hd__o22a_1
XFILLER_0_228_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold899 datamem.data_ram\[54\]\[1\] VGND VGND VPWR VPWR net2049 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2201 rvcpu.dp.rf.reg_file_arr\[13\]\[2\] VGND VGND VPWR VPWR net3351 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_71_Left_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2212 datamem.data_ram\[56\]\[20\] VGND VGND VPWR VPWR net3362 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2223 datamem.data_ram\[34\]\[9\] VGND VGND VPWR VPWR net3373 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24981_ _10474_ net3933 net101 VGND VGND VPWR VPWR _10711_ sky130_fd_sc_hd__mux2_1
Xhold2234 datamem.data_ram\[29\]\[17\] VGND VGND VPWR VPWR net3384 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1500 rvcpu.dp.rf.reg_file_arr\[15\]\[3\] VGND VGND VPWR VPWR net2650 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2245 rvcpu.dp.rf.reg_file_arr\[11\]\[26\] VGND VGND VPWR VPWR net3395 sky130_fd_sc_hd__dlygate4sd3_1
X_26720_ _10754_ net2616 _11714_ VGND VGND VPWR VPWR _11716_ sky130_fd_sc_hd__mux2_1
Xhold2256 datamem.data_ram\[29\]\[26\] VGND VGND VPWR VPWR net3406 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1511 datamem.data_ram\[46\]\[29\] VGND VGND VPWR VPWR net2661 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2267 rvcpu.dp.rf.reg_file_arr\[15\]\[10\] VGND VGND VPWR VPWR net3417 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1522 rvcpu.dp.rf.reg_file_arr\[22\]\[9\] VGND VGND VPWR VPWR net2672 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1533 rvcpu.dp.rf.reg_file_arr\[2\]\[27\] VGND VGND VPWR VPWR net2683 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2278 datamem.data_ram\[56\]\[12\] VGND VGND VPWR VPWR net3428 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1544 rvcpu.dp.rf.reg_file_arr\[19\]\[27\] VGND VGND VPWR VPWR net2694 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2289 datamem.data_ram\[4\]\[22\] VGND VGND VPWR VPWR net3439 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f__10220_ clknet_0__10220_ VGND VGND VPWR VPWR clknet_1_1__leaf__10220_
+ sky130_fd_sc_hd__clkbuf_16
Xhold1555 rvcpu.dp.rf.reg_file_arr\[28\]\[25\] VGND VGND VPWR VPWR net2705 sky130_fd_sc_hd__dlygate4sd3_1
X_26651_ _11672_ _11663_ VGND VGND VPWR VPWR _11673_ sky130_fd_sc_hd__and2_1
Xhold1566 datamem.data_ram\[9\]\[20\] VGND VGND VPWR VPWR net2716 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1577 datamem.data_ram\[8\]\[30\] VGND VGND VPWR VPWR net2727 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_165_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1588 datamem.data_ram\[25\]\[25\] VGND VGND VPWR VPWR net2738 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1599 rvcpu.dp.rf.reg_file_arr\[28\]\[19\] VGND VGND VPWR VPWR net2749 sky130_fd_sc_hd__dlygate4sd3_1
X_25602_ _11064_ _11055_ VGND VGND VPWR VPWR _11065_ sky130_fd_sc_hd__and2_1
X_22814_ rvcpu.dp.rf.reg_file_arr\[24\]\[27\] rvcpu.dp.rf.reg_file_arr\[25\]\[27\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[27\] rvcpu.dp.rf.reg_file_arr\[27\]\[27\] _09406_
+ _09395_ VGND VGND VPWR VPWR _09953_ sky130_fd_sc_hd__mux4_2
X_29370_ clknet_leaf_206_clk _01105_ VGND VGND VPWR VPWR datamem.data_ram\[60\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_26582_ _11636_ VGND VGND VPWR VPWR _03235_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_196_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28321_ _12634_ VGND VGND VPWR VPWR _03976_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_211_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25533_ _11024_ VGND VGND VPWR VPWR _02798_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1__f__10082_ clknet_0__10082_ VGND VGND VPWR VPWR clknet_1_1__leaf__10082_
+ sky130_fd_sc_hd__clkbuf_16
X_22745_ rvcpu.dp.rf.reg_file_arr\[28\]\[23\] rvcpu.dp.rf.reg_file_arr\[30\]\[23\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[23\] rvcpu.dp.rf.reg_file_arr\[31\]\[23\] _09381_
+ _09423_ VGND VGND VPWR VPWR _09888_ sky130_fd_sc_hd__mux4_1
XFILLER_0_183_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_80_Left_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28252_ _12454_ net4055 net44 VGND VGND VPWR VPWR _12596_ sky130_fd_sc_hd__mux2_1
X_25464_ _10410_ _10985_ VGND VGND VPWR VPWR _10988_ sky130_fd_sc_hd__and2_1
XFILLER_0_165_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22676_ rvcpu.dp.rf.reg_file_arr\[0\]\[19\] rvcpu.dp.rf.reg_file_arr\[1\]\[19\] rvcpu.dp.rf.reg_file_arr\[2\]\[19\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[19\] _09714_ _09585_ VGND VGND VPWR VPWR _09823_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_176_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27203_ _12005_ net1413 _12007_ _12011_ VGND VGND VPWR VPWR _03481_ sky130_fd_sc_hd__a31o_1
XFILLER_0_137_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24415_ _09272_ VGND VGND VPWR VPWR _10388_ sky130_fd_sc_hd__buf_2
X_21627_ rvcpu.dp.rf.reg_file_arr\[0\]\[12\] rvcpu.dp.rf.reg_file_arr\[1\]\[12\] rvcpu.dp.rf.reg_file_arr\[2\]\[12\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[12\] _08683_ _08684_ VGND VGND VPWR VPWR _08877_
+ sky130_fd_sc_hd__mux4_1
X_28183_ _12437_ net2675 _12555_ VGND VGND VPWR VPWR _12559_ sky130_fd_sc_hd__mux2_1
X_25395_ _10408_ _10950_ VGND VGND VPWR VPWR _10952_ sky130_fd_sc_hd__and2_1
XFILLER_0_164_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27134_ _10057_ VGND VGND VPWR VPWR _11968_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_168_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_180_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24346_ _10350_ VGND VGND VPWR VPWR _02285_ sky130_fd_sc_hd__clkbuf_1
X_21558_ _08560_ VGND VGND VPWR VPWR _08811_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_145_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20509_ datamem.data_ram\[50\]\[21\] _06613_ _07077_ datamem.data_ram\[51\]\[21\]
+ _07799_ VGND VGND VPWR VPWR _07800_ sky130_fd_sc_hd__o221a_1
XFILLER_0_133_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27065_ _11919_ net1725 _11923_ _11925_ VGND VGND VPWR VPWR _03429_ sky130_fd_sc_hd__a31o_1
X_24277_ _10311_ VGND VGND VPWR VPWR _02255_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21489_ rvcpu.dp.rf.reg_file_arr\[28\]\[6\] rvcpu.dp.rf.reg_file_arr\[30\]\[6\] rvcpu.dp.rf.reg_file_arr\[29\]\[6\]
+ rvcpu.dp.rf.reg_file_arr\[31\]\[6\] _08635_ _08637_ VGND VGND VPWR VPWR _08745_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_133_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26016_ net1306 _11329_ _11325_ _11333_ VGND VGND VPWR VPWR _02972_ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_200_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_224_5863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_224_5874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27967_ _12438_ VGND VGND VPWR VPWR _03818_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_8_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15981_ net2015 _13229_ _14322_ VGND VGND VPWR VPWR _14328_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29706_ net1052 _01441_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[22\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_17720_ _13229_ net2097 _05129_ VGND VGND VPWR VPWR _05135_ sky130_fd_sc_hd__mux2_1
X_14932_ _13328_ _13425_ VGND VGND VPWR VPWR _13481_ sky130_fd_sc_hd__nand2_1
X_26918_ _11831_ net1385 _11821_ _11836_ VGND VGND VPWR VPWR _03371_ sky130_fd_sc_hd__a31o_1
X_27898_ _11976_ _12394_ VGND VGND VPWR VPWR _12400_ sky130_fd_sc_hd__and2_1
XFILLER_0_216_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29637_ net983 _01372_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[24\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_17651_ _05098_ VGND VGND VPWR VPWR _01213_ sky130_fd_sc_hd__clkbuf_1
Xhold2790 datamem.data_ram\[21\]\[13\] VGND VGND VPWR VPWR net3940 sky130_fd_sc_hd__dlygate4sd3_1
X_14863_ _13380_ _13414_ VGND VGND VPWR VPWR _13415_ sky130_fd_sc_hd__nand2_2
XFILLER_0_215_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26849_ _11781_ net1809 _11785_ _11792_ VGND VGND VPWR VPWR _03346_ sky130_fd_sc_hd__a31o_1
XFILLER_0_188_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_203_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16602_ _04542_ VGND VGND VPWR VPWR _01738_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_19_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29568_ net922 _01303_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[26\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_17582_ _13226_ net2516 _05057_ VGND VGND VPWR VPWR _05062_ sky130_fd_sc_hd__mux2_1
X_14794_ _13286_ _13280_ VGND VGND VPWR VPWR _13347_ sky130_fd_sc_hd__or2b_1
XFILLER_0_187_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19321_ _06616_ VGND VGND VPWR VPWR _06617_ sky130_fd_sc_hd__buf_6
X_16533_ _04505_ VGND VGND VPWR VPWR _01778_ sky130_fd_sc_hd__clkbuf_1
X_28519_ _12747_ net4417 _12735_ VGND VGND VPWR VPWR _12748_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29499_ net861 _01234_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[28\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31530_ clknet_leaf_27_clk net1213 VGND VGND VPWR VPWR rvcpu.dp.plem.PCPlus4M\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19252_ _06553_ _06554_ VGND VGND VPWR VPWR _06555_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_175_4693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16464_ net2438 _14424_ _04467_ VGND VGND VPWR VPWR _04469_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_183_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18203_ _05504_ _05567_ VGND VGND VPWR VPWR _05568_ sky130_fd_sc_hd__or2_1
X_23694__289 clknet_1_1__leaf__10195_ VGND VGND VPWR VPWR net415 sky130_fd_sc_hd__inv_2
X_15415_ _13431_ _13628_ _13423_ _13945_ _13946_ VGND VGND VPWR VPWR _13947_ sky130_fd_sc_hd__o311a_1
XFILLER_0_171_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19183_ rvcpu.dp.plde.ImmExtE\[21\] rvcpu.dp.plde.PCE\[21\] VGND VGND VPWR VPWR _06495_
+ sky130_fd_sc_hd__nor2_1
X_31461_ clknet_leaf_75_clk rvcpu.dp.SrcBFW_Mux.y\[19\] VGND VGND VPWR VPWR rvcpu.dp.plem.WriteDataM\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16395_ _14563_ VGND VGND VPWR VPWR _01842_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18134_ rvcpu.dp.plde.RD1E\[17\] _05292_ _05499_ VGND VGND VPWR VPWR _05500_ sky130_fd_sc_hd__o21a_2
X_30412_ net750 _02147_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[31\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_15346_ _13428_ _13880_ _13881_ VGND VGND VPWR VPWR _13882_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_113_3206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31392_ clknet_leaf_40_clk _03095_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCE\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_3217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_887 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__10240_ clknet_0__10240_ VGND VGND VPWR VPWR clknet_1_0__leaf__10240_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_108_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18065_ _05432_ VGND VGND VPWR VPWR _05433_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_78_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30343_ net689 _02078_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[4\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_15277_ _13630_ _13776_ _13798_ _13441_ VGND VGND VPWR VPWR _13816_ sky130_fd_sc_hd__a31o_1
XFILLER_0_151_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_184_4907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold107 rvcpu.dp.plem.ALUResultM\[9\] VGND VGND VPWR VPWR net1257 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__10171_ clknet_0__10171_ VGND VGND VPWR VPWR clknet_1_0__leaf__10171_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_184_4918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold118 rvcpu.dp.plem.RegWriteM VGND VGND VPWR VPWR net1268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 rvcpu.dp.plem.ALUResultM\[22\] VGND VGND VPWR VPWR net1279 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_145_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17016_ net4401 _14430_ _04757_ VGND VGND VPWR VPWR _04762_ sky130_fd_sc_hd__mux2_1
XFILLER_0_229_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30274_ net628 _02009_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[6\]\[29\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_74_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32013_ clknet_leaf_128_clk _03435_ VGND VGND VPWR VPWR datamem.data_ram\[27\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23134__810 clknet_1_1__leaf__10106_ VGND VGND VPWR VPWR net936 sky130_fd_sc_hd__inv_2
XFILLER_0_95_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18967_ _05554_ _05730_ _06301_ _06303_ VGND VGND VPWR VPWR _06304_ sky130_fd_sc_hd__a211o_1
XFILLER_0_219_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_225_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_3925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17918_ _05252_ _05263_ VGND VGND VPWR VPWR _05291_ sky130_fd_sc_hd__nand2_4
XFILLER_0_193_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18898_ _05461_ _06238_ VGND VGND VPWR VPWR _06239_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_217_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32915_ clknet_leaf_164_clk _04337_ VGND VGND VPWR VPWR datamem.data_ram\[0\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_17849_ _05226_ _05227_ VGND VGND VPWR VPWR rvcpu.dp.SrcBFW_Mux.y\[13\] sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_33_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32846_ clknet_leaf_86_clk _04268_ VGND VGND VPWR VPWR datamem.data_ram\[7\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20860_ datamem.data_ram\[8\]\[14\] _06648_ _06658_ datamem.data_ram\[9\]\[14\] VGND
+ VGND VPWR VPWR _08150_ sky130_fd_sc_hd__o22a_1
XFILLER_0_117_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19519_ _06661_ VGND VGND VPWR VPWR _06815_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_102_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32777_ clknet_leaf_159_clk _04199_ VGND VGND VPWR VPWR datamem.data_ram\[14\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_20791_ _08078_ _08079_ _08080_ _06712_ VGND VGND VPWR VPWR _08081_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_102_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22530_ rvcpu.dp.rf.reg_file_arr\[8\]\[11\] rvcpu.dp.rf.reg_file_arr\[10\]\[11\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[11\] rvcpu.dp.rf.reg_file_arr\[11\]\[11\] _09424_
+ _09485_ VGND VGND VPWR VPWR _09685_ sky130_fd_sc_hd__mux4_1
X_31728_ net177 _03186_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[9\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22461_ rvcpu.dp.rf.reg_file_arr\[20\]\[8\] rvcpu.dp.rf.reg_file_arr\[21\]\[8\] rvcpu.dp.rf.reg_file_arr\[22\]\[8\]
+ rvcpu.dp.rf.reg_file_arr\[23\]\[8\] _09512_ _09408_ VGND VGND VPWR VPWR _09619_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_88_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31659_ clknet_leaf_64_clk net1986 VGND VGND VPWR VPWR rvcpu.dp.plmw.ALUResultW\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_24200_ _10268_ _09301_ _10269_ VGND VGND VPWR VPWR _10270_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_8_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21412_ _08662_ _08667_ _08671_ _08625_ VGND VGND VPWR VPWR _01030_ sky130_fd_sc_hd__o31a_1
XFILLER_0_127_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23221__871 clknet_1_0__leaf__10124_ VGND VGND VPWR VPWR net997 sky130_fd_sc_hd__inv_2
X_25180_ _10826_ net1873 net58 VGND VGND VPWR VPWR _10827_ sky130_fd_sc_hd__mux2_1
XFILLER_0_228_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22392_ _09534_ _09553_ VGND VGND VPWR VPWR _09554_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21343_ rvcpu.ALUResultE\[14\] rvcpu.ALUResultE\[17\] _08603_ _08604_ VGND VGND VPWR
+ VPWR _08605_ sky130_fd_sc_hd__or4_1
XFILLER_0_161_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_559 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold630 datamem.data_ram\[11\]\[1\] VGND VGND VPWR VPWR net1780 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21274_ _08535_ VGND VGND VPWR VPWR _08536_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold641 datamem.data_ram\[2\]\[2\] VGND VGND VPWR VPWR net1791 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold652 rvcpu.dp.plfd.PCD\[24\] VGND VGND VPWR VPWR net1802 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold663 datamem.data_ram\[19\]\[6\] VGND VGND VPWR VPWR net1813 sky130_fd_sc_hd__dlygate4sd3_1
X_20225_ datamem.data_ram\[10\]\[3\] _06932_ _06955_ datamem.data_ram\[12\]\[3\] VGND
+ VGND VPWR VPWR _07518_ sky130_fd_sc_hd__a22o_1
XFILLER_0_198_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold674 _02944_ VGND VGND VPWR VPWR net1824 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28870_ _12700_ net3099 _12932_ VGND VGND VPWR VPWR _12939_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold685 datamem.data_ram\[53\]\[5\] VGND VGND VPWR VPWR net1835 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_204_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold696 datamem.data_ram\[25\]\[7\] VGND VGND VPWR VPWR net1846 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_228_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27821_ _12353_ VGND VGND VPWR VPWR _03757_ sky130_fd_sc_hd__clkbuf_1
X_20156_ datamem.data_ram\[25\]\[27\] _06657_ VGND VGND VPWR VPWR _07449_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_5_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2020 datamem.data_ram\[53\]\[21\] VGND VGND VPWR VPWR net3170 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2031 rvcpu.dp.rf.reg_file_arr\[16\]\[27\] VGND VGND VPWR VPWR net3181 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2042 datamem.data_ram\[21\]\[10\] VGND VGND VPWR VPWR net3192 sky130_fd_sc_hd__dlygate4sd3_1
X_27752_ _12315_ VGND VGND VPWR VPWR _03726_ sky130_fd_sc_hd__clkbuf_1
Xhold2053 datamem.data_ram\[35\]\[28\] VGND VGND VPWR VPWR net3203 sky130_fd_sc_hd__dlygate4sd3_1
X_24964_ _10701_ VGND VGND VPWR VPWR _02552_ sky130_fd_sc_hd__clkbuf_1
X_20087_ datamem.data_ram\[50\]\[10\] _06802_ _06780_ datamem.data_ram\[49\]\[10\]
+ _06732_ VGND VGND VPWR VPWR _07381_ sky130_fd_sc_hd__o221a_1
Xhold2064 datamem.data_ram\[47\]\[21\] VGND VGND VPWR VPWR net3214 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2075 rvcpu.dp.rf.reg_file_arr\[23\]\[17\] VGND VGND VPWR VPWR net3225 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1330 rvcpu.dp.rf.reg_file_arr\[17\]\[1\] VGND VGND VPWR VPWR net2480 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2086 rvcpu.dp.rf.reg_file_arr\[26\]\[31\] VGND VGND VPWR VPWR net3236 sky130_fd_sc_hd__dlygate4sd3_1
X_26703_ _11706_ VGND VGND VPWR VPWR _03286_ sky130_fd_sc_hd__clkbuf_1
Xhold1341 rvcpu.dp.rf.reg_file_arr\[1\]\[18\] VGND VGND VPWR VPWR net2491 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2097 datamem.data_ram\[62\]\[21\] VGND VGND VPWR VPWR net3247 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1352 datamem.data_ram\[31\]\[20\] VGND VGND VPWR VPWR net2502 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1363 datamem.data_ram\[5\]\[28\] VGND VGND VPWR VPWR net2513 sky130_fd_sc_hd__dlygate4sd3_1
X_27683_ _12278_ VGND VGND VPWR VPWR _03694_ sky130_fd_sc_hd__clkbuf_1
X_24895_ _10664_ VGND VGND VPWR VPWR _02520_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1374 datamem.data_ram\[25\]\[23\] VGND VGND VPWR VPWR net2524 sky130_fd_sc_hd__dlygate4sd3_1
X_29422_ clknet_leaf_97_clk _01157_ VGND VGND VPWR VPWR datamem.data_ram\[5\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1385 rvcpu.dp.rf.reg_file_arr\[14\]\[29\] VGND VGND VPWR VPWR net2535 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f__10203_ clknet_0__10203_ VGND VGND VPWR VPWR clknet_1_1__leaf__10203_
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_503 _11679_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26634_ _10268_ _11054_ _11609_ VGND VGND VPWR VPWR _11663_ sky130_fd_sc_hd__and3_1
Xhold1396 rvcpu.dp.rf.reg_file_arr\[22\]\[3\] VGND VGND VPWR VPWR net2546 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_514 _13223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_525 _13260_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_536 rvcpu.dp.plmw.ReadDataW\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29353_ clknet_leaf_145_clk _01088_ VGND VGND VPWR VPWR datamem.data_ram\[61\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__10134_ clknet_0__10134_ VGND VGND VPWR VPWR clknet_1_1__leaf__10134_
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_547 _06780_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26565_ _11627_ VGND VGND VPWR VPWR _03227_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_558 _07912_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20989_ datamem.data_ram\[0\]\[15\] datamem.data_ram\[1\]\[15\] _06650_ VGND VGND
+ VPWR VPWR _08278_ sky130_fd_sc_hd__mux2_1
X_23777_ clknet_1_0__leaf__10078_ VGND VGND VPWR VPWR _10203_ sky130_fd_sc_hd__buf_1
XFILLER_0_178_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_569 _06744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_28304_ _12625_ VGND VGND VPWR VPWR _03968_ sky130_fd_sc_hd__clkbuf_1
X_25516_ _10991_ net1398 _11009_ _11014_ VGND VGND VPWR VPWR _02791_ sky130_fd_sc_hd__a31o_1
XFILLER_0_137_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29284_ _13163_ VGND VGND VPWR VPWR _04410_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22728_ rvcpu.dp.rf.reg_file_arr\[24\]\[22\] rvcpu.dp.rf.reg_file_arr\[25\]\[22\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[22\] rvcpu.dp.rf.reg_file_arr\[27\]\[22\] _09393_
+ _09465_ VGND VGND VPWR VPWR _09872_ sky130_fd_sc_hd__mux4_1
XFILLER_0_211_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28235_ _12437_ net3653 _12583_ VGND VGND VPWR VPWR _12587_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_188_5007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25447_ _10600_ _10980_ VGND VGND VPWR VPWR _10981_ sky130_fd_sc_hd__nor2_4
XFILLER_0_137_366 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_188_5018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22659_ rvcpu.dp.rf.reg_file_arr\[4\]\[18\] rvcpu.dp.rf.reg_file_arr\[5\]\[18\] rvcpu.dp.rf.reg_file_arr\[6\]\[18\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[18\] _09604_ _09716_ VGND VGND VPWR VPWR _09807_
+ sky130_fd_sc_hd__mux4_1
X_15200_ _13385_ _13672_ _13741_ _13598_ VGND VGND VPWR VPWR _13742_ sky130_fd_sc_hd__or4b_1
XPHY_EDGE_ROW_173_Right_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_213_5597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28166_ _12363_ net2281 _12546_ VGND VGND VPWR VPWR _12550_ sky130_fd_sc_hd__mux2_1
X_16180_ _13206_ VGND VGND VPWR VPWR _14438_ sky130_fd_sc_hd__buf_4
X_25378_ _10413_ _10936_ VGND VGND VPWR VPWR _10941_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_211_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27117_ _11956_ net1704 _11952_ _11957_ VGND VGND VPWR VPWR _03449_ sky130_fd_sc_hd__a31o_1
X_15131_ _13330_ _13603_ _13673_ _13675_ _13475_ VGND VGND VPWR VPWR _13676_ sky130_fd_sc_hd__a41o_1
XFILLER_0_180_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24329_ _09240_ net4306 _10338_ VGND VGND VPWR VPWR _10341_ sky130_fd_sc_hd__mux2_1
X_28097_ _12513_ VGND VGND VPWR VPWR _03873_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_226_5914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_226_5925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15062_ _13607_ _13473_ _13608_ VGND VGND VPWR VPWR _13609_ sky130_fd_sc_hd__o21a_1
X_27048_ _11904_ datamem.data_ram\[52\]\[2\] _11910_ _11914_ VGND VGND VPWR VPWR _03423_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_160_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_4014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_147_4025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19870_ _06604_ _07156_ _07158_ _07164_ VGND VGND VPWR VPWR _07165_ sky130_fd_sc_hd__o31a_1
XFILLER_0_102_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18821_ _05516_ _06165_ _05497_ VGND VGND VPWR VPWR _06167_ sky130_fd_sc_hd__o21ai_1
X_28999_ _10142_ _10935_ _10921_ VGND VGND VPWR VPWR _13010_ sky130_fd_sc_hd__and3_2
XFILLER_0_156_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18752_ _06090_ _06091_ _06092_ _06102_ VGND VGND VPWR VPWR _06103_ sky130_fd_sc_hd__a31o_1
X_15964_ net2609 _13204_ _14311_ VGND VGND VPWR VPWR _14319_ sky130_fd_sc_hd__mux2_1
XFILLER_0_223_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_216_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_222_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17703_ _13204_ net2937 _05118_ VGND VGND VPWR VPWR _05126_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_106_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14915_ _13425_ _13434_ VGND VGND VPWR VPWR _13465_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_106_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18683_ _05419_ _06036_ VGND VGND VPWR VPWR _06037_ sky130_fd_sc_hd__nand2_1
X_30961_ clknet_leaf_153_clk _02696_ VGND VGND VPWR VPWR datamem.data_ram\[3\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15895_ _14282_ VGND VGND VPWR VPWR _02077_ sky130_fd_sc_hd__clkbuf_1
X_32700_ clknet_leaf_233_clk _04122_ VGND VGND VPWR VPWR datamem.data_ram\[17\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_17634_ _05089_ VGND VGND VPWR VPWR _01221_ sky130_fd_sc_hd__clkbuf_1
X_14846_ rvcpu.dp.pcreg.q\[3\] _13280_ VGND VGND VPWR VPWR _13399_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_177_4733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_177_4744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30892_ clknet_leaf_194_clk _02627_ VGND VGND VPWR VPWR datamem.data_ram\[42\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_177_4755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32631_ clknet_leaf_90_clk _04053_ VGND VGND VPWR VPWR datamem.data_ram\[1\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_67_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23164__836 clknet_1_1__leaf__10110_ VGND VGND VPWR VPWR net962 sky130_fd_sc_hd__inv_2
X_17565_ _13201_ net2705 _05046_ VGND VGND VPWR VPWR _05053_ sky130_fd_sc_hd__mux2_1
X_14777_ _13283_ _13329_ VGND VGND VPWR VPWR _13330_ sky130_fd_sc_hd__or2_2
XFILLER_0_86_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_187_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23702__296 clknet_1_0__leaf__10196_ VGND VGND VPWR VPWR net422 sky130_fd_sc_hd__inv_2
X_19304_ _06599_ VGND VGND VPWR VPWR _06600_ sky130_fd_sc_hd__clkbuf_16
X_23776__364 clknet_1_0__leaf__10202_ VGND VGND VPWR VPWR net490 sky130_fd_sc_hd__inv_2
X_16516_ net2099 _14476_ _04489_ VGND VGND VPWR VPWR _04496_ sky130_fd_sc_hd__mux2_1
X_32562_ clknet_leaf_87_clk _03984_ VGND VGND VPWR VPWR datamem.data_ram\[22\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17496_ _05016_ VGND VGND VPWR VPWR _01294_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31513_ clknet_leaf_52_clk net1188 VGND VGND VPWR VPWR rvcpu.dp.plem.PCPlus4M\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_19235_ rvcpu.dp.plde.ImmExtE\[28\] rvcpu.dp.plde.PCE\[28\] VGND VGND VPWR VPWR _06540_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_156_664 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16447_ _04458_ VGND VGND VPWR VPWR _01817_ sky130_fd_sc_hd__clkbuf_1
X_32493_ clknet_leaf_78_clk _03915_ VGND VGND VPWR VPWR datamem.data_ram\[25\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_136_3751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_140_Right_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_3762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19166_ rvcpu.dp.plde.ImmExtE\[19\] rvcpu.dp.plde.PCE\[19\] VGND VGND VPWR VPWR _06480_
+ sky130_fd_sc_hd__nor2_1
X_31444_ clknet_leaf_7_clk rvcpu.dp.SrcBFW_Mux.y\[2\] VGND VGND VPWR VPWR rvcpu.dp.plem.WriteDataM\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_27_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16378_ net2174 _14476_ _14547_ VGND VGND VPWR VPWR _14554_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_76_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1271 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18117_ rvcpu.dp.plde.RD1E\[19\] _05292_ _05483_ VGND VGND VPWR VPWR _05484_ sky130_fd_sc_hd__o21a_2
XFILLER_0_42_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15329_ _13449_ _13694_ _13865_ _13455_ _13357_ VGND VGND VPWR VPWR _13866_ sky130_fd_sc_hd__o32a_1
X_19097_ _06418_ rvcpu.dp.plde.ImmExtE\[10\] _06419_ VGND VGND VPWR VPWR _06420_ sky130_fd_sc_hd__mux2_1
XFILLER_0_182_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31375_ clknet_leaf_18_clk _03078_ VGND VGND VPWR VPWR rvcpu.dp.plde.ImmExtE\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_3659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__10223_ clknet_0__10223_ VGND VGND VPWR VPWR clknet_1_0__leaf__10223_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_223_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18048_ _05412_ _05415_ VGND VGND VPWR VPWR _05417_ sky130_fd_sc_hd__nor2_1
X_30326_ net672 _02061_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[4\]\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_39_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__10154_ clknet_0__10154_ VGND VGND VPWR VPWR clknet_1_0__leaf__10154_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_223_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30257_ net611 _01992_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[6\]\[12\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f__10085_ clknet_0__10085_ VGND VGND VPWR VPWR clknet_1_0__leaf__10085_
+ sky130_fd_sc_hd__clkbuf_16
X_20010_ datamem.data_ram\[57\]\[2\] _06948_ _07301_ _07303_ VGND VGND VPWR VPWR _07304_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_1_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30188_ net542 _01923_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[8\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_19999_ datamem.data_ram\[30\]\[2\] _06950_ _06947_ datamem.data_ram\[25\]\[2\] VGND
+ VGND VPWR VPWR _07293_ sky130_fd_sc_hd__a22o_1
XFILLER_0_226_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24002__535 clknet_1_0__leaf__10241_ VGND VGND VPWR VPWR net661 sky130_fd_sc_hd__inv_2
XFILLER_0_20_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23482__129 clknet_1_1__leaf__10159_ VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__inv_2
XFILLER_0_225_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21961_ _08532_ _09190_ _09192_ _08699_ VGND VGND VPWR VPWR _09193_ sky130_fd_sc_hd__a211o_1
XFILLER_0_222_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_206_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23700_ clknet_1_0__leaf__10192_ VGND VGND VPWR VPWR _10196_ sky130_fd_sc_hd__buf_1
X_20912_ _08199_ _08200_ _08201_ _07822_ _07868_ VGND VGND VPWR VPWR _08202_ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24680_ _10392_ net3507 _10543_ VGND VGND VPWR VPWR _10547_ sky130_fd_sc_hd__mux2_1
X_21892_ _08514_ _09126_ VGND VGND VPWR VPWR _09127_ sky130_fd_sc_hd__or2_1
XFILLER_0_221_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20843_ _08132_ VGND VGND VPWR VPWR _08133_ sky130_fd_sc_hd__buf_6
X_32829_ clknet_leaf_153_clk _04251_ VGND VGND VPWR VPWR datamem.data_ram\[12\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26350_ _10070_ _11507_ _11508_ net1340 VGND VGND VPWR VPWR _03131_ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_620 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20774_ datamem.data_ram\[56\]\[6\] _07122_ _07133_ datamem.data_ram\[57\]\[6\] VGND
+ VGND VPWR VPWR _08064_ sky130_fd_sc_hd__a22o_1
XFILLER_0_159_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25301_ _10893_ VGND VGND VPWR VPWR _02697_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22513_ _09482_ _09668_ VGND VGND VPWR VPWR _09669_ sky130_fd_sc_hd__or2_1
X_26281_ net1838 _11467_ VGND VGND VPWR VPWR _11473_ sky130_fd_sc_hd__and2_1
XFILLER_0_92_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_170_clk clknet_5_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_170_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_134_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28020_ _12371_ net2001 _12464_ VGND VGND VPWR VPWR _12472_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25232_ _10855_ VGND VGND VPWR VPWR _02666_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_146_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22444_ rvcpu.dp.rf.reg_file_arr\[0\]\[7\] rvcpu.dp.rf.reg_file_arr\[1\]\[7\] rvcpu.dp.rf.reg_file_arr\[2\]\[7\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[7\] _09417_ _09585_ VGND VGND VPWR VPWR _09603_ sky130_fd_sc_hd__mux4_1
XFILLER_0_73_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25163_ _10815_ VGND VGND VPWR VPWR _02637_ sky130_fd_sc_hd__clkbuf_1
X_22375_ _09389_ _09526_ _09531_ _09537_ VGND VGND VPWR VPWR _09538_ sky130_fd_sc_hd__and4_1
XFILLER_0_32_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21326_ _08584_ _08585_ _08587_ VGND VGND VPWR VPWR _08588_ sky130_fd_sc_hd__and3b_2
X_25094_ _09231_ VGND VGND VPWR VPWR _10780_ sky130_fd_sc_hd__buf_4
X_29971_ net341 _01706_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[15\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23417__70 clknet_1_0__leaf__10153_ VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__inv_2
X_28922_ _12966_ VGND VGND VPWR VPWR _04245_ sky130_fd_sc_hd__clkbuf_1
Xhold460 datamem.data_ram\[11\]\[4\] VGND VGND VPWR VPWR net1610 sky130_fd_sc_hd__dlygate4sd3_1
X_21257_ _08518_ VGND VGND VPWR VPWR _08519_ sky130_fd_sc_hd__buf_4
XFILLER_0_64_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold471 rvcpu.dp.plfd.PCPlus4D\[31\] VGND VGND VPWR VPWR net1621 sky130_fd_sc_hd__dlygate4sd3_1
Xhold482 datamem.data_ram\[27\]\[3\] VGND VGND VPWR VPWR net1632 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_221_5800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold493 datamem.data_ram\[50\]\[5\] VGND VGND VPWR VPWR net1643 sky130_fd_sc_hd__dlygate4sd3_1
X_20208_ datamem.data_ram\[52\]\[11\] _06766_ _07500_ _06769_ VGND VGND VPWR VPWR
+ _07501_ sky130_fd_sc_hd__o211a_1
XFILLER_0_229_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_221_5811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28853_ _12747_ net4385 _12923_ VGND VGND VPWR VPWR _12930_ sky130_fd_sc_hd__mux2_1
X_21188_ _07277_ _07119_ _07070_ _06915_ VGND VGND VPWR VPWR _08474_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_102_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23432__84 clknet_1_0__leaf__10154_ VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__inv_2
X_27804_ _12140_ net3198 _12336_ VGND VGND VPWR VPWR _12344_ sky130_fd_sc_hd__mux2_1
X_20139_ datamem.data_ram\[46\]\[27\] _06627_ _06821_ datamem.data_ram\[40\]\[27\]
+ VGND VGND VPWR VPWR _07432_ sky130_fd_sc_hd__o22a_1
X_28784_ _12893_ VGND VGND VPWR VPWR _04180_ sky130_fd_sc_hd__clkbuf_1
X_25996_ _08513_ _11315_ _11312_ _11322_ VGND VGND VPWR VPWR _02963_ sky130_fd_sc_hd__o211a_1
XFILLER_0_204_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27735_ _12306_ VGND VGND VPWR VPWR _03718_ sky130_fd_sc_hd__clkbuf_1
X_24947_ _10692_ VGND VGND VPWR VPWR _02544_ sky130_fd_sc_hd__clkbuf_1
Xhold1160 rvcpu.dp.rf.reg_file_arr\[7\]\[29\] VGND VGND VPWR VPWR net2310 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1171 rvcpu.dp.pcreg.q\[29\] VGND VGND VPWR VPWR net2321 sky130_fd_sc_hd__dlygate4sd3_1
X_14700_ _13259_ VGND VGND VPWR VPWR _13260_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_73_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1182 datamem.data_ram\[40\]\[31\] VGND VGND VPWR VPWR net2332 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15680_ _14157_ VGND VGND VPWR VPWR _02175_ sky130_fd_sc_hd__clkbuf_1
X_27666_ _12269_ VGND VGND VPWR VPWR _03686_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_219_5740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_300 _13921_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1193 rvcpu.dp.rf.reg_file_arr\[10\]\[7\] VGND VGND VPWR VPWR net2343 sky130_fd_sc_hd__dlygate4sd3_1
X_24878_ _10655_ VGND VGND VPWR VPWR _02512_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_311 _14170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_219_5751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29405_ clknet_leaf_0_clk _01140_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD2E\[16\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_322 _14445_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_219_5762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_333 _14459_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14631_ net2391 _13207_ _13181_ VGND VGND VPWR VPWR _13208_ sky130_fd_sc_hd__mux2_1
X_26617_ _11656_ VGND VGND VPWR VPWR _03250_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23829_ _09298_ net3407 _10210_ VGND VGND VPWR VPWR _10211_ sky130_fd_sc_hd__mux2_1
X_27597_ _12232_ VGND VGND VPWR VPWR _03654_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_344 _14478_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23228__877 clknet_1_0__leaf__10125_ VGND VGND VPWR VPWR net1003 sky130_fd_sc_hd__inv_2
XFILLER_0_185_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_355 rvcpu.dp.SrcBFW_Mux.y\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_366 rvcpu.dp.plde.ImmExtE\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_377 rvcpu.dp.plmw.ReadDataW\[29\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17350_ _04939_ VGND VGND VPWR VPWR _01363_ sky130_fd_sc_hd__clkbuf_1
X_29336_ clknet_leaf_271_clk _01071_ VGND VGND VPWR VPWR datamem.data_ram\[62\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26548_ _11104_ VGND VGND VPWR VPWR _11618_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_215_5648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_388 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_215_5659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_4630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_399 _06610_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16301_ _14513_ VGND VGND VPWR VPWR _01886_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17281_ net4312 _13172_ _04902_ VGND VGND VPWR VPWR _04903_ sky130_fd_sc_hd__mux2_1
X_29267_ _13154_ VGND VGND VPWR VPWR _04402_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_222_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26479_ rvcpu.dp.plde.JalrE VGND VGND VPWR VPWR _11598_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_161_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_161_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_83_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19020_ rvcpu.dp.plde.ImmExtE\[0\] rvcpu.dp.plde.PCE\[0\] VGND VGND VPWR VPWR _06353_
+ sky130_fd_sc_hd__or2_1
X_28218_ _12363_ net3558 net45 VGND VGND VPWR VPWR _12578_ sky130_fd_sc_hd__mux2_1
X_16232_ _14473_ VGND VGND VPWR VPWR _01923_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__10079_ _10079_ VGND VGND VPWR VPWR clknet_0__10079_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_222_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29198_ _09317_ net3025 _13112_ VGND VGND VPWR VPWR _13117_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload308 clknet_1_0__leaf__10195_ VGND VGND VPWR VPWR clkload308/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload319 clknet_1_1__leaf__10159_ VGND VGND VPWR VPWR clkload319/Y sky130_fd_sc_hd__clkinvlp_4
X_28149_ _12454_ net3709 net73 VGND VGND VPWR VPWR _12541_ sky130_fd_sc_hd__mux2_1
X_16163_ net2258 _14426_ _14422_ VGND VGND VPWR VPWR _14427_ sky130_fd_sc_hd__mux2_1
Xclkload16 clknet_5_19__leaf_clk VGND VGND VPWR VPWR clkload16/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload27 clknet_leaf_15_clk VGND VGND VPWR VPWR clkload27/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_3_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload38 clknet_leaf_9_clk VGND VGND VPWR VPWR clkload38/Y sky130_fd_sc_hd__clkinv_4
Xclkload49 clknet_leaf_45_clk VGND VGND VPWR VPWR clkload49/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_2_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15114_ _13658_ _13484_ VGND VGND VPWR VPWR _13659_ sky130_fd_sc_hd__nor2_2
X_31160_ clknet_leaf_68_clk rvcpu.ALUResultE\[19\] VGND VGND VPWR VPWR rvcpu.dp.plem.ALUResultM\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16094_ net2688 _13190_ _14385_ VGND VGND VPWR VPWR _14389_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30111_ net473 _01846_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[10\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_15045_ _13282_ _13415_ VGND VGND VPWR VPWR _13592_ sky130_fd_sc_hd__nand2_1
X_19922_ datamem.data_ram\[58\]\[17\] _06612_ _07215_ _07216_ VGND VGND VPWR VPWR
+ _07217_ sky130_fd_sc_hd__o211a_1
X_31091_ clknet_leaf_95_clk _02826_ VGND VGND VPWR VPWR datamem.data_ram\[21\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_4478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_4489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30042_ net404 _01777_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[13\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_19853_ datamem.data_ram\[58\]\[1\] _06932_ _06973_ datamem.data_ram\[56\]\[1\] VGND
+ VGND VPWR VPWR _07148_ sky130_fd_sc_hd__a22o_1
XFILLER_0_208_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18804_ _05454_ _05513_ _05510_ VGND VGND VPWR VPWR _06151_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_207_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19784_ datamem.data_ram\[46\]\[9\] _06763_ _06611_ datamem.data_ram\[42\]\[9\] VGND
+ VGND VPWR VPWR _07079_ sky130_fd_sc_hd__o22a_1
X_16996_ _04750_ VGND VGND VPWR VPWR _01544_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_30_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18735_ _05436_ _06082_ _05331_ VGND VGND VPWR VPWR _06086_ sky130_fd_sc_hd__a21oi_1
X_15947_ _14309_ VGND VGND VPWR VPWR _02052_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_69_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31993_ clknet_leaf_127_clk _03415_ VGND VGND VPWR VPWR datamem.data_ram\[31\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_69_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_3485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_3496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30944_ clknet_leaf_95_clk _02679_ VGND VGND VPWR VPWR datamem.data_ram\[3\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_18666_ _05809_ _06019_ _06020_ VGND VGND VPWR VPWR _06021_ sky130_fd_sc_hd__and3_1
X_15878_ rvcpu.dp.plmw.RdW\[0\] rvcpu.dp.plmw.RdW\[1\] rvcpu.dp.plmw.RegWriteW VGND
+ VGND VPWR VPWR _14272_ sky130_fd_sc_hd__or3b_1
XFILLER_0_204_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14829_ _13379_ _13381_ _13331_ VGND VGND VPWR VPWR _13382_ sky130_fd_sc_hd__o21a_1
X_17617_ _13278_ net3570 _05045_ VGND VGND VPWR VPWR _05080_ sky130_fd_sc_hd__mux2_1
X_30875_ clknet_leaf_61_clk _02610_ VGND VGND VPWR VPWR datamem.data_ram\[42\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_18597_ _05356_ _05361_ _05404_ _05886_ _05954_ VGND VGND VPWR VPWR _05955_ sky130_fd_sc_hd__a311oi_1
XFILLER_0_148_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_175_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_3813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_188_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32614_ clknet_leaf_82_clk _04036_ VGND VGND VPWR VPWR datamem.data_ram\[20\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17548_ _05043_ VGND VGND VPWR VPWR _01269_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32545_ clknet_leaf_252_clk _03967_ VGND VGND VPWR VPWR datamem.data_ram\[23\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_152_clk clknet_5_28__leaf_clk VGND VGND VPWR VPWR clknet_leaf_152_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_132_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17479_ _14193_ net3699 _04973_ VGND VGND VPWR VPWR _05007_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19218_ _06525_ rvcpu.dp.plde.ImmExtE\[25\] _06493_ VGND VGND VPWR VPWR _06526_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20490_ rvcpu.dp.plem.ALUResultM\[1\] _07737_ _07781_ rvcpu.dp.plem.ALUResultM\[0\]
+ VGND VGND VPWR VPWR _07782_ sky130_fd_sc_hd__o22a_1
XFILLER_0_132_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32476_ clknet_leaf_253_clk _03898_ VGND VGND VPWR VPWR datamem.data_ram\[26\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22960__669 clknet_1_1__leaf__10081_ VGND VGND VPWR VPWR net795 sky130_fd_sc_hd__inv_2
X_31427_ clknet_leaf_99_clk _03130_ VGND VGND VPWR VPWR datamem.data_ram\[44\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_19149_ _06463_ _06464_ VGND VGND VPWR VPWR _06465_ sky130_fd_sc_hd__or2b_1
XFILLER_0_171_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22160_ _07123_ VGND VGND VPWR VPWR _09350_ sky130_fd_sc_hd__buf_12
X_31358_ clknet_leaf_22_clk _03061_ VGND VGND VPWR VPWR rvcpu.dp.plde.ImmExtE\[7\]
+ sky130_fd_sc_hd__dfxtp_2
Xclkbuf_1_0__f__10206_ clknet_0__10206_ VGND VGND VPWR VPWR clknet_1_0__leaf__10206_
+ sky130_fd_sc_hd__clkbuf_16
X_21111_ datamem.data_ram\[23\]\[7\] _06924_ _06953_ datamem.data_ram\[20\]\[7\] _08399_
+ VGND VGND VPWR VPWR _08400_ sky130_fd_sc_hd__a221o_1
XFILLER_0_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30309_ net655 _02044_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[5\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_22091_ rvcpu.dp.plem.WriteDataM\[1\] _08488_ _09293_ _09295_ rvcpu.dp.plem.WriteDataM\[9\]
+ VGND VGND VPWR VPWR _09304_ sky130_fd_sc_hd__a32o_1
X_31289_ clknet_leaf_108_clk _02992_ VGND VGND VPWR VPWR datamem.data_ram\[34\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_58_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__10137_ clknet_0__10137_ VGND VGND VPWR VPWR clknet_1_0__leaf__10137_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_58_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23333__972 clknet_1_1__leaf__10135_ VGND VGND VPWR VPWR net1098 sky130_fd_sc_hd__inv_2
X_21042_ datamem.data_ram\[9\]\[31\] _06655_ _08330_ _06599_ VGND VGND VPWR VPWR _08331_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_160_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_226_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25850_ rvcpu.dp.plfd.PCPlus4D\[26\] _11231_ _11142_ VGND VGND VPWR VPWR _11232_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24801_ _10442_ net4155 _10612_ VGND VGND VPWR VPWR _10614_ sky130_fd_sc_hd__mux2_1
X_25781_ _11146_ VGND VGND VPWR VPWR _11177_ sky130_fd_sc_hd__clkbuf_4
X_27520_ _12087_ net4081 net99 VGND VGND VPWR VPWR _12192_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24732_ _10446_ net3098 _10571_ VGND VGND VPWR VPWR _10575_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23112__790 clknet_1_1__leaf__10104_ VGND VGND VPWR VPWR net916 sky130_fd_sc_hd__inv_2
X_21944_ _08547_ _09174_ _09176_ _08652_ VGND VGND VPWR VPWR _09177_ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27451_ _09284_ VGND VGND VPWR VPWR _12153_ sky130_fd_sc_hd__buf_2
XFILLER_0_194_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24663_ _10067_ _10532_ VGND VGND VPWR VPWR _10537_ sky130_fd_sc_hd__and2_1
XFILLER_0_222_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21875_ _09109_ _09110_ _08673_ VGND VGND VPWR VPWR _09111_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26402_ _13706_ _11542_ _11544_ _11534_ VGND VGND VPWR VPWR _03147_ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27382_ _12110_ VGND VGND VPWR VPWR _03561_ sky130_fd_sc_hd__clkbuf_1
X_20826_ datamem.data_ram\[13\]\[30\] _06663_ _08115_ _07851_ VGND VGND VPWR VPWR
+ _08116_ sky130_fd_sc_hd__o22a_1
X_24594_ _10398_ net3448 _10491_ VGND VGND VPWR VPWR _10498_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29121_ _10979_ _10114_ _12977_ VGND VGND VPWR VPWR _13076_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_37_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26333_ _11086_ _11497_ VGND VGND VPWR VPWR _11502_ sky130_fd_sc_hd__and2_1
XFILLER_0_135_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20757_ datamem.data_ram\[4\]\[6\] datamem.data_ram\[5\]\[6\] _07828_ VGND VGND VPWR
+ VPWR _08047_ sky130_fd_sc_hd__mux2_1
XFILLER_0_175_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_143_clk clknet_5_29__leaf_clk VGND VGND VPWR VPWR clknet_leaf_143_clk
+ sky130_fd_sc_hd__clkbuf_8
X_29052_ _13018_ net1767 _13030_ _13039_ VGND VGND VPWR VPWR _04302_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_210_5534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26264_ net1801 _11432_ VGND VGND VPWR VPWR _11464_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_210_5545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20688_ datamem.data_ram\[54\]\[5\] _06978_ _07000_ datamem.data_ram\[50\]\[5\] VGND
+ VGND VPWR VPWR _07979_ sky130_fd_sc_hd__a22o_1
XFILLER_0_163_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_208_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28003_ _12462_ net3778 _12448_ VGND VGND VPWR VPWR _12463_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25215_ _10846_ VGND VGND VPWR VPWR _02658_ sky130_fd_sc_hd__clkbuf_1
X_22427_ rvcpu.dp.rf.reg_file_arr\[4\]\[6\] rvcpu.dp.rf.reg_file_arr\[5\]\[6\] rvcpu.dp.rf.reg_file_arr\[6\]\[6\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[6\] _09423_ _09424_ VGND VGND VPWR VPWR _09587_ sky130_fd_sc_hd__mux4_1
X_26195_ rvcpu.ALUControl\[3\] _11432_ VGND VGND VPWR VPWR _11435_ sky130_fd_sc_hd__and2_1
XFILLER_0_162_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25146_ _10805_ VGND VGND VPWR VPWR _02630_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22358_ rvcpu.dp.rf.reg_file_arr\[24\]\[3\] rvcpu.dp.rf.reg_file_arr\[25\]\[3\] rvcpu.dp.rf.reg_file_arr\[26\]\[3\]
+ rvcpu.dp.rf.reg_file_arr\[27\]\[3\] _09392_ _09394_ VGND VGND VPWR VPWR _09521_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_27_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21309_ rvcpu.dp.rf.reg_file_arr\[4\]\[0\] rvcpu.dp.rf.reg_file_arr\[5\]\[0\] rvcpu.dp.rf.reg_file_arr\[6\]\[0\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[0\] _08567_ _08570_ VGND VGND VPWR VPWR _08571_ sky130_fd_sc_hd__mux4_1
X_25077_ _10727_ net4036 _10768_ VGND VGND VPWR VPWR _10770_ sky130_fd_sc_hd__mux2_1
X_29954_ net324 _01689_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[15\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_22289_ rvcpu.dp.rf.reg_file_arr\[28\]\[1\] rvcpu.dp.rf.reg_file_arr\[30\]\[1\] rvcpu.dp.rf.reg_file_arr\[29\]\[1\]
+ rvcpu.dp.rf.reg_file_arr\[31\]\[1\] _09443_ _09453_ VGND VGND VPWR VPWR _09454_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_208_5485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28905_ _12957_ VGND VGND VPWR VPWR _04237_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_208_5496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold290 datamem.data_ram\[56\]\[6\] VGND VGND VPWR VPWR net1440 sky130_fd_sc_hd__dlygate4sd3_1
X_29885_ net263 _01620_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[17\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16850_ _04673_ VGND VGND VPWR VPWR _01613_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28836_ _12764_ net4060 _12914_ VGND VGND VPWR VPWR _12921_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_161_4353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_4364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15801_ _14230_ VGND VGND VPWR VPWR _02127_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_217_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16781_ net3033 _14468_ _04634_ VGND VGND VPWR VPWR _04637_ sky130_fd_sc_hd__mux2_1
X_28767_ _12700_ net2925 _12877_ VGND VGND VPWR VPWR _12884_ sky130_fd_sc_hd__mux2_1
XFILLER_0_204_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25979_ _13932_ _11268_ VGND VGND VPWR VPWR _11313_ sky130_fd_sc_hd__nand2_1
X_18520_ _05374_ _05732_ VGND VGND VPWR VPWR _05881_ sky130_fd_sc_hd__nor2_1
XFILLER_0_204_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23545__170 clknet_1_0__leaf__10173_ VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__inv_2
X_15732_ _14192_ VGND VGND VPWR VPWR _02158_ sky130_fd_sc_hd__clkbuf_1
X_27718_ _12297_ VGND VGND VPWR VPWR _03710_ sky130_fd_sc_hd__clkbuf_1
X_28698_ _12847_ VGND VGND VPWR VPWR _04140_ sky130_fd_sc_hd__clkbuf_1
X_18451_ _05810_ _05791_ VGND VGND VPWR VPWR _05814_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_64_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27649_ _10500_ VGND VGND VPWR VPWR _12260_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_64_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15663_ _14145_ net4382 _14131_ VGND VGND VPWR VPWR _14146_ sky130_fd_sc_hd__mux2_1
XANTENNA_130 _07808_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_198_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_141 _07836_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_152 _07874_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17402_ _04966_ VGND VGND VPWR VPWR _01338_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_120_3371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14614_ _13194_ VGND VGND VPWR VPWR _13195_ sky130_fd_sc_hd__buf_4
X_18382_ _05652_ rvcpu.dp.plde.ALUControlE\[1\] _05722_ _05745_ VGND VGND VPWR VPWR
+ _05746_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_120_3382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_163 _08634_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_30660_ clknet_leaf_198_clk _02395_ VGND VGND VPWR VPWR datamem.data_ram\[50\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15594_ net2242 _13217_ _14103_ VGND VGND VPWR VPWR _14105_ sky130_fd_sc_hd__mux2_1
XANTENNA_174 _08780_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_185 _09094_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_196 _09351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29319_ clknet_leaf_11_clk _01054_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD1E\[26\] sky130_fd_sc_hd__dfxtp_1
X_17333_ net4440 _13259_ _04924_ VGND VGND VPWR VPWR _04930_ sky130_fd_sc_hd__mux2_1
X_30591_ clknet_leaf_92_clk _02326_ VGND VGND VPWR VPWR datamem.data_ram\[53\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_134_clk clknet_5_27__leaf_clk VGND VGND VPWR VPWR clknet_leaf_134_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_138_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32330_ clknet_leaf_259_clk _03752_ VGND VGND VPWR VPWR datamem.data_ram\[31\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17264_ _14183_ net3894 _04887_ VGND VGND VPWR VPWR _04893_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19003_ _06335_ _06336_ VGND VGND VPWR VPWR _06337_ sky130_fd_sc_hd__and2_1
XFILLER_0_181_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16215_ net3320 _14461_ _14443_ VGND VGND VPWR VPWR _14462_ sky130_fd_sc_hd__mux2_1
Xclkload105 clknet_leaf_158_clk VGND VGND VPWR VPWR clkload105/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_24_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32261_ clknet_leaf_241_clk _03683_ VGND VGND VPWR VPWR datamem.data_ram\[34\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload116 clknet_leaf_95_clk VGND VGND VPWR VPWR clkload116/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_12_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17195_ _04856_ VGND VGND VPWR VPWR _01443_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_168_4518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload127 clknet_leaf_255_clk VGND VGND VPWR VPWR clkload127/Y sky130_fd_sc_hd__clkinv_1
X_23814__397 clknet_1_0__leaf__10207_ VGND VGND VPWR VPWR net523 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_168_4529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31212_ clknet_leaf_40_clk net1365 VGND VGND VPWR VPWR rvcpu.dp.plfd.PCD\[1\] sky130_fd_sc_hd__dfxtp_1
Xclkload138 clknet_leaf_243_clk VGND VGND VPWR VPWR clkload138/Y sky130_fd_sc_hd__inv_6
Xclkload149 clknet_leaf_271_clk VGND VGND VPWR VPWR clkload149/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_94_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16146_ net2070 _13269_ _14407_ VGND VGND VPWR VPWR _14416_ sky130_fd_sc_hd__mux2_1
XFILLER_0_178_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32192_ clknet_leaf_276_clk _03614_ VGND VGND VPWR VPWR datamem.data_ram\[37\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_94_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31143_ clknet_leaf_66_clk rvcpu.ALUResultE\[2\] VGND VGND VPWR VPWR rvcpu.dp.plem.ALUResultM\[2\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16077_ _14379_ VGND VGND VPWR VPWR _01984_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_90_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_911 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15028_ _13574_ _13546_ VGND VGND VPWR VPWR _13575_ sky130_fd_sc_hd__or2_1
X_19905_ datamem.data_ram\[9\]\[17\] _06659_ _07198_ _07199_ VGND VGND VPWR VPWR _07200_
+ sky130_fd_sc_hd__o211a_1
X_31074_ clknet_leaf_91_clk _02809_ VGND VGND VPWR VPWR datamem.data_ram\[9\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2608 datamem.data_ram\[58\]\[31\] VGND VGND VPWR VPWR net3758 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2619 datamem.data_ram\[7\]\[22\] VGND VGND VPWR VPWR net3769 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_127_3536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30025_ net387 _01760_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[13\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19836_ _06777_ VGND VGND VPWR VPWR _07131_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_127_3547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23628__245 clknet_1_0__leaf__10181_ VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__inv_2
XFILLER_0_120_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1907 rvcpu.dp.rf.reg_file_arr\[13\]\[13\] VGND VGND VPWR VPWR net3057 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1918 datamem.data_ram\[18\]\[13\] VGND VGND VPWR VPWR net3068 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1929 datamem.data_ram\[14\]\[26\] VGND VGND VPWR VPWR net3079 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19767_ datamem.data_ram\[22\]\[25\] _06683_ _06739_ datamem.data_ram\[19\]\[25\]
+ _07061_ VGND VGND VPWR VPWR _07062_ sky130_fd_sc_hd__o221a_1
XFILLER_0_224_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16979_ _04741_ VGND VGND VPWR VPWR _01552_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_194_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18718_ _05436_ _06069_ VGND VGND VPWR VPWR _06070_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_88_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19698_ datamem.data_ram\[14\]\[0\] _06952_ _06961_ datamem.data_ram\[11\]\[0\] VGND
+ VGND VPWR VPWR _06994_ sky130_fd_sc_hd__a22o_1
X_31976_ clknet_leaf_138_clk _03398_ VGND VGND VPWR VPWR datamem.data_ram\[53\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_188_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_204_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18649_ _05604_ _05596_ _05664_ VGND VGND VPWR VPWR _06005_ sky130_fd_sc_hd__mux2_1
X_30927_ clknet_leaf_151_clk _02662_ VGND VGND VPWR VPWR datamem.data_ram\[40\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_189_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30858_ clknet_leaf_137_clk _02593_ VGND VGND VPWR VPWR datamem.data_ram\[43\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_21660_ rvcpu.dp.rf.reg_file_arr\[0\]\[14\] rvcpu.dp.rf.reg_file_arr\[1\]\[14\] rvcpu.dp.rf.reg_file_arr\[2\]\[14\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[14\] _08810_ _08811_ VGND VGND VPWR VPWR _08908_
+ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20611_ datamem.data_ram\[46\]\[13\] _06682_ _06806_ datamem.data_ram\[44\]\[13\]
+ VGND VGND VPWR VPWR _07902_ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_125_clk clknet_5_30__leaf_clk VGND VGND VPWR VPWR clknet_leaf_125_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_188_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21591_ rvcpu.dp.rf.reg_file_arr\[8\]\[10\] rvcpu.dp.rf.reg_file_arr\[10\]\[10\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[10\] rvcpu.dp.rf.reg_file_arr\[11\]\[10\] _08649_
+ _08537_ VGND VGND VPWR VPWR _08843_ sky130_fd_sc_hd__mux4_1
X_30789_ clknet_leaf_264_clk _02524_ VGND VGND VPWR VPWR datamem.data_ram\[46\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20542_ _07832_ VGND VGND VPWR VPWR _07833_ sky130_fd_sc_hd__buf_6
X_32528_ clknet_leaf_275_clk _03950_ VGND VGND VPWR VPWR datamem.data_ram\[24\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20473_ datamem.data_ram\[37\]\[20\] _06662_ _06781_ datamem.data_ram\[33\]\[20\]
+ VGND VGND VPWR VPWR _07765_ sky130_fd_sc_hd__o22a_1
XFILLER_0_104_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32459_ clknet_leaf_241_clk _03881_ VGND VGND VPWR VPWR datamem.data_ram\[26\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25000_ _10450_ net2522 _10715_ VGND VGND VPWR VPWR _10721_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22212_ _09291_ net2306 _09371_ VGND VGND VPWR VPWR _09379_ sky130_fd_sc_hd__mux2_1
X_23192_ _09236_ datamem.data_ram\[5\]\[17\] _10115_ VGND VGND VPWR VPWR _10117_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22143_ _09299_ _09269_ _09231_ VGND VGND VPWR VPWR _09341_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_30_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24008__541 clknet_1_1__leaf__10241_ VGND VGND VPWR VPWR net667 sky130_fd_sc_hd__inv_2
XFILLER_0_2_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_679 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26951_ _11849_ net1547 _11853_ _11857_ VGND VGND VPWR VPWR _03383_ sky130_fd_sc_hd__a31o_1
XFILLER_0_100_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22074_ _09289_ VGND VGND VPWR VPWR _01074_ sky130_fd_sc_hd__clkbuf_1
X_25902_ net1593 _11181_ _11258_ _11269_ VGND VGND VPWR VPWR _02922_ sky130_fd_sc_hd__o211a_1
X_21025_ datamem.data_ram\[28\]\[31\] datamem.data_ram\[29\]\[31\] _07911_ VGND VGND
+ VPWR VPWR _08314_ sky130_fd_sc_hd__mux2_1
X_29670_ net1016 _01405_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[23\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_26882_ _11752_ VGND VGND VPWR VPWR _11813_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_226_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_203_5360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28621_ _12754_ net4175 _12805_ VGND VGND VPWR VPWR _12807_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_203_5371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25833_ rvcpu.dp.pcreg.q\[23\] _11213_ VGND VGND VPWR VPWR _11218_ sky130_fd_sc_hd__xor2_1
XFILLER_0_173_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28552_ _12690_ net3377 _12768_ VGND VGND VPWR VPWR _12770_ sky130_fd_sc_hd__mux2_1
X_25764_ net1571 _11144_ _11147_ _11164_ VGND VGND VPWR VPWR _02889_ sky130_fd_sc_hd__o211a_1
XFILLER_0_173_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_195_5172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27503_ _12149_ net2294 _12179_ VGND VGND VPWR VPWR _12183_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_195_5183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24715_ _10565_ VGND VGND VPWR VPWR _02439_ sky130_fd_sc_hd__clkbuf_1
X_28483_ _12391_ net1685 _12723_ _12725_ VGND VGND VPWR VPWR _04047_ sky130_fd_sc_hd__a31o_1
XFILLER_0_179_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21927_ _09160_ VGND VGND VPWR VPWR _01056_ sky130_fd_sc_hd__clkbuf_1
X_25695_ _11105_ net1687 _11111_ _11119_ VGND VGND VPWR VPWR _02865_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27434_ _12141_ VGND VGND VPWR VPWR _03582_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_191_5069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24646_ _10396_ net3722 _10521_ VGND VGND VPWR VPWR _10527_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21858_ rvcpu.dp.rf.reg_file_arr\[24\]\[25\] rvcpu.dp.rf.reg_file_arr\[25\]\[25\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[25\] rvcpu.dp.rf.reg_file_arr\[27\]\[25\] _08525_
+ _08528_ VGND VGND VPWR VPWR _09095_ sky130_fd_sc_hd__mux4_1
XFILLER_0_167_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20809_ _08097_ _08098_ _07820_ VGND VGND VPWR VPWR _08099_ sky130_fd_sc_hd__mux2_1
X_27365_ _12087_ net4265 _12097_ VGND VGND VPWR VPWR _12101_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_116_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_116_clk
+ sky130_fd_sc_hd__clkbuf_8
X_24577_ _10452_ net3550 _10482_ VGND VGND VPWR VPWR _10489_ sky130_fd_sc_hd__mux2_1
X_21789_ _08510_ _09029_ VGND VGND VPWR VPWR _09030_ sky130_fd_sc_hd__nor2_1
XFILLER_0_203_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29104_ _12601_ _10092_ _12977_ VGND VGND VPWR VPWR _13067_ sky130_fd_sc_hd__a21oi_4
X_26316_ net1651 _11436_ VGND VGND VPWR VPWR _11491_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_4190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27296_ _11918_ VGND VGND VPWR VPWR _12061_ sky130_fd_sc_hd__buf_2
XFILLER_0_80_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29035_ _13029_ VGND VGND VPWR VPWR _13030_ sky130_fd_sc_hd__clkbuf_2
X_26247_ _11438_ _11458_ _11459_ _09457_ VGND VGND VPWR VPWR _03077_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_123_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_150_4087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16000_ net4282 _13257_ _14333_ VGND VGND VPWR VPWR _14338_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_4098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26178_ _08567_ _11413_ VGND VGND VPWR VPWR _11426_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25129_ _10796_ VGND VGND VPWR VPWR _02622_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_221_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_4404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_4415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17951_ _05321_ _05226_ _05227_ _05322_ VGND VGND VPWR VPWR _05323_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_20_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29937_ net307 _01672_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[16\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_23119__796 clknet_1_1__leaf__10105_ VGND VGND VPWR VPWR net922 sky130_fd_sc_hd__inv_2
XFILLER_0_228_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16902_ net2366 _14453_ _04695_ VGND VGND VPWR VPWR _04701_ sky130_fd_sc_hd__mux2_1
X_17882_ rvcpu.dp.plmw.RdW\[4\] rvcpu.dp.plde.Rs1E\[4\] VGND VGND VPWR VPWR _05255_
+ sky130_fd_sc_hd__and2b_1
X_29868_ net246 _01603_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[18\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19621_ _05371_ _06641_ VGND VGND VPWR VPWR _06917_ sky130_fd_sc_hd__nand2_8
XFILLER_0_219_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16833_ _04664_ VGND VGND VPWR VPWR _01621_ sky130_fd_sc_hd__clkbuf_1
X_28819_ _12700_ net3539 _12905_ VGND VGND VPWR VPWR _12912_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29799_ clknet_leaf_198_clk _01534_ VGND VGND VPWR VPWR datamem.data_ram\[59\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_122_3422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31830_ clknet_leaf_105_clk _03284_ VGND VGND VPWR VPWR datamem.data_ram\[16\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_122_3433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16764_ net2696 _14451_ _04623_ VGND VGND VPWR VPWR _04628_ sky130_fd_sc_hd__mux2_1
X_19552_ datamem.data_ram\[13\]\[24\] _06823_ _06789_ datamem.data_ram\[9\]\[24\]
+ VGND VGND VPWR VPWR _06848_ sky130_fd_sc_hd__o22a_1
XFILLER_0_219_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_100_Left_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18503_ _05275_ _05709_ _05864_ VGND VGND VPWR VPWR _05865_ sky130_fd_sc_hd__and3_1
X_15715_ _13256_ VGND VGND VPWR VPWR _14181_ sky130_fd_sc_hd__buf_4
X_31761_ clknet_leaf_107_clk _03215_ VGND VGND VPWR VPWR datamem.data_ram\[18\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_19483_ _06778_ VGND VGND VPWR VPWR _06779_ sky130_fd_sc_hd__buf_6
X_16695_ _04591_ VGND VGND VPWR VPWR _01694_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_201_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30712_ clknet_leaf_138_clk _02447_ VGND VGND VPWR VPWR datamem.data_ram\[49\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18434_ _05674_ _05796_ VGND VGND VPWR VPWR _05797_ sky130_fd_sc_hd__or2_1
X_15646_ _14134_ VGND VGND VPWR VPWR _02186_ sky130_fd_sc_hd__clkbuf_1
X_31692_ clknet_leaf_39_clk _03150_ VGND VGND VPWR VPWR rvcpu.dp.pcreg.q\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_556 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30643_ clknet_leaf_139_clk _02378_ VGND VGND VPWR VPWR datamem.data_ram\[51\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18365_ _05729_ VGND VGND VPWR VPWR _05730_ sky130_fd_sc_hd__buf_2
XFILLER_0_150_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_107_clk clknet_5_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_107_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_200_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15577_ net2511 _13190_ _14092_ VGND VGND VPWR VPWR _14096_ sky130_fd_sc_hd__mux2_1
XFILLER_0_200_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17316_ net4402 _13234_ _04913_ VGND VGND VPWR VPWR _04921_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18296_ _05658_ _05660_ VGND VGND VPWR VPWR _05661_ sky130_fd_sc_hd__nor2_2
X_30574_ clknet_leaf_190_clk _02309_ VGND VGND VPWR VPWR datamem.data_ram\[54\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32313_ clknet_leaf_230_clk _03735_ VGND VGND VPWR VPWR datamem.data_ram\[31\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_17247_ _14166_ net3209 _04876_ VGND VGND VPWR VPWR _04884_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_92_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32244_ clknet_leaf_225_clk _03666_ VGND VGND VPWR VPWR datamem.data_ram\[34\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17178_ _04847_ VGND VGND VPWR VPWR _01451_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16129_ _14384_ VGND VGND VPWR VPWR _14407_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32175_ clknet_leaf_194_clk _03597_ VGND VGND VPWR VPWR datamem.data_ram\[37\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3106 datamem.data_ram\[54\]\[13\] VGND VGND VPWR VPWR net4256 sky130_fd_sc_hd__dlygate4sd3_1
X_31126_ clknet_leaf_125_clk _02861_ VGND VGND VPWR VPWR datamem.data_ram\[25\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3117 rvcpu.dp.rf.reg_file_arr\[1\]\[10\] VGND VGND VPWR VPWR net4267 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_161_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold3128 datamem.data_ram\[13\]\[9\] VGND VGND VPWR VPWR net4278 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3139 rvcpu.dp.rf.reg_file_arr\[15\]\[23\] VGND VGND VPWR VPWR net4289 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2405 datamem.data_ram\[58\]\[26\] VGND VGND VPWR VPWR net3555 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2416 datamem.data_ram\[7\]\[21\] VGND VGND VPWR VPWR net3566 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31057_ clknet_leaf_114_clk _02792_ VGND VGND VPWR VPWR datamem.data_ram\[38\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_51_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2427 datamem.data_ram\[57\]\[10\] VGND VGND VPWR VPWR net3577 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2438 rvcpu.dp.rf.reg_file_arr\[29\]\[19\] VGND VGND VPWR VPWR net3588 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1704 datamem.data_ram\[16\]\[30\] VGND VGND VPWR VPWR net2854 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2449 datamem.data_ram\[17\]\[13\] VGND VGND VPWR VPWR net3599 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_3989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30008_ clknet_leaf_266_clk _01743_ VGND VGND VPWR VPWR datamem.data_ram\[59\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1715 datamem.data_ram\[45\]\[26\] VGND VGND VPWR VPWR net2865 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1726 datamem.data_ram\[24\]\[18\] VGND VGND VPWR VPWR net2876 sky130_fd_sc_hd__dlygate4sd3_1
X_19819_ datamem.data_ram\[26\]\[9\] _06611_ _06634_ datamem.data_ram\[27\]\[9\] _06601_
+ VGND VGND VPWR VPWR _07114_ sky130_fd_sc_hd__o221a_1
Xhold1737 rvcpu.dp.rf.reg_file_arr\[3\]\[9\] VGND VGND VPWR VPWR net2887 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1748 datamem.data_ram\[0\]\[26\] VGND VGND VPWR VPWR net2898 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_5_25__f_clk clknet_2_3_0_clk VGND VGND VPWR VPWR clknet_5_25__leaf_clk sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_81_Right_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1759 datamem.data_ram\[22\]\[30\] VGND VGND VPWR VPWR net2909 sky130_fd_sc_hd__dlygate4sd3_1
X_22830_ _09705_ _09960_ _09964_ _09968_ VGND VGND VPWR VPWR _09969_ sky130_fd_sc_hd__and4_1
XFILLER_0_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_205_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22761_ _09511_ _09902_ VGND VGND VPWR VPWR _09903_ sky130_fd_sc_hd__or2_1
X_31959_ clknet_leaf_120_clk _03381_ VGND VGND VPWR VPWR datamem.data_ram\[28\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24038__567 clknet_1_0__leaf__10245_ VGND VGND VPWR VPWR net693 sky130_fd_sc_hd__inv_2
X_24500_ _10441_ VGND VGND VPWR VPWR _02348_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_49_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_220_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_188_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21712_ rvcpu.dp.rf.reg_file_arr\[24\]\[17\] rvcpu.dp.rf.reg_file_arr\[25\]\[17\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[17\] rvcpu.dp.rf.reg_file_arr\[27\]\[17\] _08536_
+ _08693_ VGND VGND VPWR VPWR _08957_ sky130_fd_sc_hd__mux4_1
X_25480_ _10058_ net35 _10996_ net1311 VGND VGND VPWR VPWR _02773_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22692_ _09390_ _09837_ VGND VGND VPWR VPWR _09838_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_192_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24431_ _10398_ net4418 _10386_ VGND VGND VPWR VPWR _10399_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21643_ rvcpu.dp.rf.reg_file_arr\[4\]\[13\] rvcpu.dp.rf.reg_file_arr\[5\]\[13\] rvcpu.dp.rf.reg_file_arr\[6\]\[13\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[13\] _08687_ _08856_ VGND VGND VPWR VPWR _08892_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_164_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27150_ _11978_ _11966_ VGND VGND VPWR VPWR _11979_ sky130_fd_sc_hd__and2_1
XFILLER_0_90_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24362_ _09306_ net3456 net61 VGND VGND VPWR VPWR _10359_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21574_ rvcpu.dp.rf.reg_file_arr\[20\]\[10\] rvcpu.dp.rf.reg_file_arr\[21\]\[10\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[10\] rvcpu.dp.rf.reg_file_arr\[23\]\[10\] _08778_
+ _08825_ VGND VGND VPWR VPWR _08826_ sky130_fd_sc_hd__mux4_1
XANTENNA_30 _06634_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_41 _06677_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26101_ _11385_ VGND VGND VPWR VPWR _03004_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_52 _06688_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_90_Right_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_63 _06751_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27081_ rvcpu.ALUResultE\[0\] _06354_ _11598_ VGND VGND VPWR VPWR _11934_ sky130_fd_sc_hd__mux2_1
X_20525_ datamem.data_ram\[16\]\[21\] _06649_ _06636_ datamem.data_ram\[19\]\[21\]
+ _06777_ VGND VGND VPWR VPWR _07816_ sky130_fd_sc_hd__o221a_1
XFILLER_0_90_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_74 _06776_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24293_ _09279_ net3404 _10316_ VGND VGND VPWR VPWR _10320_ sky130_fd_sc_hd__mux2_1
XANTENNA_85 _06784_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_96 _06810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26032_ _11083_ _11340_ VGND VGND VPWR VPWR _11343_ sky130_fd_sc_hd__and2_1
X_20456_ datamem.data_ram\[30\]\[20\] _06628_ _07230_ datamem.data_ram\[28\]\[20\]
+ VGND VGND VPWR VPWR _07748_ sky130_fd_sc_hd__o22a_1
XFILLER_0_160_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20387_ _06751_ _07673_ _07678_ VGND VGND VPWR VPWR _07679_ sky130_fd_sc_hd__or3_1
XFILLER_0_219_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_205_5411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_205_5422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22126_ _09299_ _09229_ _09231_ VGND VGND VPWR VPWR _09332_ sky130_fd_sc_hd__a21oi_4
X_27983_ _12449_ VGND VGND VPWR VPWR _03823_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26934_ _11803_ _11842_ VGND VGND VPWR VPWR _11847_ sky130_fd_sc_hd__and2_1
X_29722_ net1068 _01457_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[22\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_201_5308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22057_ _09276_ net3409 _09270_ VGND VGND VPWR VPWR _09277_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_201_5319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_197_5212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_197_5223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21008_ _07176_ _08284_ _08296_ _06592_ VGND VGND VPWR VPWR _08297_ sky130_fd_sc_hd__a22o_1
Xhold2950 datamem.data_ram\[26\]\[29\] VGND VGND VPWR VPWR net4100 sky130_fd_sc_hd__dlygate4sd3_1
X_26865_ _11795_ net1469 _11797_ _11802_ VGND VGND VPWR VPWR _03352_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_197_5234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2961 datamem.data_ram\[33\]\[9\] VGND VGND VPWR VPWR net4111 sky130_fd_sc_hd__dlygate4sd3_1
X_29653_ net999 _01388_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[24\]\[16\] sky130_fd_sc_hd__dfxtp_1
Xhold2972 datamem.data_ram\[20\]\[25\] VGND VGND VPWR VPWR net4122 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2983 rvcpu.dp.rf.reg_file_arr\[22\]\[20\] VGND VGND VPWR VPWR net4133 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25816_ rvcpu.dp.pcreg.q\[20\] _11200_ VGND VGND VPWR VPWR _11204_ sky130_fd_sc_hd__or2_1
XFILLER_0_173_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28604_ _12690_ net3300 _12796_ VGND VGND VPWR VPWR _12798_ sky130_fd_sc_hd__mux2_1
Xhold2994 datamem.data_ram\[11\]\[31\] VGND VGND VPWR VPWR net4144 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29584_ net938 _01319_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[26\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_26796_ _11760_ VGND VGND VPWR VPWR _11761_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_3_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28535_ _12758_ net3305 _12752_ VGND VGND VPWR VPWR _12759_ sky130_fd_sc_hd__mux2_1
XFILLER_0_186_106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25747_ _08588_ _08597_ rvcpu.dp.hu.ResultSrcE0 VGND VGND VPWR VPWR _11151_ sky130_fd_sc_hd__o21a_1
Xmax_cap43 _12735_ VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__buf_4
Xmax_cap54 _11021_ VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__buf_4
XFILLER_0_134_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap65 _13040_ VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__buf_4
X_15500_ _13475_ _14025_ _14026_ _14027_ VGND VGND VPWR VPWR _14028_ sky130_fd_sc_hd__o211a_1
XFILLER_0_186_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap76 _12448_ VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_4
XFILLER_0_57_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap87 _10793_ VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_156_4230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16480_ net3095 _14440_ _04467_ VGND VGND VPWR VPWR _04477_ sky130_fd_sc_hd__mux2_1
X_28466_ _12715_ VGND VGND VPWR VPWR _04040_ sky130_fd_sc_hd__clkbuf_1
X_25678_ _11105_ net4342 _11097_ _11108_ VGND VGND VPWR VPWR _02859_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_156_4241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap98 _12206_ VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__buf_4
X_15431_ _13431_ _13432_ _13613_ _13333_ VGND VGND VPWR VPWR _13962_ sky130_fd_sc_hd__a211o_1
X_27417_ _09239_ VGND VGND VPWR VPWR _12130_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_194_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_182_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24629_ _10517_ VGND VGND VPWR VPWR _02401_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_14_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28397_ _12441_ net4021 _12669_ VGND VGND VPWR VPWR _12675_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_183_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_152_4138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18150_ _05502_ _05510_ VGND VGND VPWR VPWR _05515_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_152_4149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15362_ _13466_ _13841_ VGND VGND VPWR VPWR _13897_ sky130_fd_sc_hd__or2_1
XFILLER_0_183_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27348_ _12090_ VGND VGND VPWR VPWR _03547_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17101_ _14156_ net3113 _04804_ VGND VGND VPWR VPWR _04807_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18081_ _05446_ _05409_ VGND VGND VPWR VPWR _05449_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15293_ _13415_ _13510_ VGND VGND VPWR VPWR _13831_ sky130_fd_sc_hd__or2_1
X_27279_ _10826_ net4225 _12043_ VGND VGND VPWR VPWR _12051_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17032_ _04770_ VGND VGND VPWR VPWR _01520_ sky130_fd_sc_hd__clkbuf_1
X_29018_ _12734_ net2607 net66 VGND VGND VPWR VPWR _13021_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23273__918 clknet_1_0__leaf__10129_ VGND VGND VPWR VPWR net1044 sky130_fd_sc_hd__inv_2
X_30290_ net636 _02025_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[5\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_229_5989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_186_4960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_186_4971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_221_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18983_ _05703_ _06312_ _06318_ VGND VGND VPWR VPWR _06319_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_182_4857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_4868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17934_ rvcpu.dp.plem.ALUResultM\[14\] _05272_ _05270_ _13234_ _05306_ VGND VGND
+ VPWR VPWR _05307_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_178_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32931_ clknet_leaf_147_clk _04353_ VGND VGND VPWR VPWR datamem.data_ram\[7\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17865_ rvcpu.dp.plde.ALUControlE\[0\] _00003_ VGND VGND VPWR VPWR _05238_ sky130_fd_sc_hd__nor2_1
X_24185__25 clknet_1_0__leaf__10266_ VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__inv_2
XFILLER_0_84_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_206_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_205_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_191_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19604_ datamem.data_ram\[21\]\[8\] _06723_ _06726_ datamem.data_ram\[23\]\[8\] VGND
+ VGND VPWR VPWR _06900_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_1_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16816_ _04655_ VGND VGND VPWR VPWR _01629_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_85_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32862_ clknet_leaf_55_clk _04284_ VGND VGND VPWR VPWR datamem.data_ram\[11\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_85_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17796_ _05190_ VGND VGND VPWR VPWR rvcpu.dp.SrcBFW_Mux.y\[3\] sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_85_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_141_3875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31813_ clknet_leaf_109_clk _03267_ VGND VGND VPWR VPWR datamem.data_ram\[17\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_19535_ datamem.data_ram\[34\]\[24\] _06689_ _06668_ datamem.data_ram\[39\]\[24\]
+ VGND VGND VPWR VPWR _06831_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_187_Right_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_141_3886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16747_ net4229 _14434_ _04612_ VGND VGND VPWR VPWR _04619_ sky130_fd_sc_hd__mux2_1
XFILLER_0_191_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32793_ clknet_leaf_234_clk _04215_ VGND VGND VPWR VPWR datamem.data_ram\[13\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_19466_ datamem.data_ram\[48\]\[16\] _06697_ _06761_ datamem.data_ram\[55\]\[16\]
+ VGND VGND VPWR VPWR _06762_ sky130_fd_sc_hd__o22a_1
X_16678_ _04582_ VGND VGND VPWR VPWR _01702_ sky130_fd_sc_hd__clkbuf_1
X_31744_ net129 _03202_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[9\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_174_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18417_ _05590_ _05375_ VGND VGND VPWR VPWR _05781_ sky130_fd_sc_hd__nor2_2
XFILLER_0_57_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15629_ net2380 _13269_ _14114_ VGND VGND VPWR VPWR _14123_ sky130_fd_sc_hd__mux2_1
X_31675_ clknet_leaf_8_clk net1282 VGND VGND VPWR VPWR rvcpu.dp.plmw.ALUResultW\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_19397_ datamem.data_ram\[2\]\[16\] _06692_ _06635_ datamem.data_ram\[3\]\[16\] VGND
+ VGND VPWR VPWR _06693_ sky130_fd_sc_hd__o22a_1
XFILLER_0_146_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18348_ _05539_ _05545_ _05666_ VGND VGND VPWR VPWR _05713_ sky130_fd_sc_hd__mux2_1
X_30626_ clknet_leaf_191_clk _02361_ VGND VGND VPWR VPWR datamem.data_ram\[52\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_228_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18279_ _05643_ _05301_ VGND VGND VPWR VPWR _05644_ sky130_fd_sc_hd__or2_1
X_30557_ clknet_leaf_217_clk _02292_ VGND VGND VPWR VPWR datamem.data_ram\[54\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23671__268 clknet_1_0__leaf__10193_ VGND VGND VPWR VPWR net394 sky130_fd_sc_hd__inv_2
XFILLER_0_44_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20310_ datamem.data_ram\[6\]\[4\] _06978_ _06943_ datamem.data_ram\[3\]\[4\] VGND
+ VGND VPWR VPWR _07602_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21290_ rvcpu.dp.plfd.InstrD\[16\] VGND VGND VPWR VPWR _08552_ sky130_fd_sc_hd__buf_4
XFILLER_0_13_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30488_ clknet_leaf_204_clk _02223_ VGND VGND VPWR VPWR datamem.data_ram\[57\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold801 datamem.data_ram\[46\]\[31\] VGND VGND VPWR VPWR net1951 sky130_fd_sc_hd__dlygate4sd3_1
Xhold812 rvcpu.dp.plfd.PCPlus4D\[30\] VGND VGND VPWR VPWR net1962 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_226_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20241_ datamem.data_ram\[50\]\[3\] _07136_ _07530_ _07533_ VGND VGND VPWR VPWR _07534_
+ sky130_fd_sc_hd__a211o_1
Xhold823 rvcpu.dp.rf.reg_file_arr\[6\]\[22\] VGND VGND VPWR VPWR net1973 sky130_fd_sc_hd__dlygate4sd3_1
X_32227_ clknet_leaf_170_clk _03649_ VGND VGND VPWR VPWR datamem.data_ram\[35\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold834 rvcpu.dp.rf.reg_file_arr\[11\]\[22\] VGND VGND VPWR VPWR net1984 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold845 datamem.data_ram\[2\]\[14\] VGND VGND VPWR VPWR net1995 sky130_fd_sc_hd__dlygate4sd3_1
Xhold856 rvcpu.dp.rf.reg_file_arr\[9\]\[4\] VGND VGND VPWR VPWR net2006 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold867 datamem.data_ram\[0\]\[21\] VGND VGND VPWR VPWR net2017 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32158_ clknet_leaf_88_clk _03580_ VGND VGND VPWR VPWR datamem.data_ram\[38\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20172_ datamem.data_ram\[29\]\[11\] _06865_ _06863_ datamem.data_ram\[27\]\[11\]
+ _07464_ VGND VGND VPWR VPWR _07465_ sky130_fd_sc_hd__o221a_1
Xhold878 rvcpu.dp.rf.reg_file_arr\[3\]\[21\] VGND VGND VPWR VPWR net2028 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold889 rvcpu.dp.rf.reg_file_arr\[3\]\[29\] VGND VGND VPWR VPWR net2039 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31109_ clknet_leaf_60_clk _02844_ VGND VGND VPWR VPWR datamem.data_ram\[43\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2202 datamem.data_ram\[30\]\[12\] VGND VGND VPWR VPWR net3352 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2213 rvcpu.dp.rf.reg_file_arr\[13\]\[12\] VGND VGND VPWR VPWR net3363 sky130_fd_sc_hd__dlygate4sd3_1
X_32089_ clknet_leaf_234_clk _03511_ VGND VGND VPWR VPWR datamem.data_ram\[8\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_24980_ _10710_ VGND VGND VPWR VPWR _02559_ sky130_fd_sc_hd__clkbuf_1
Xhold2224 datamem.data_ram\[55\]\[26\] VGND VGND VPWR VPWR net3374 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2235 datamem.data_ram\[32\]\[17\] VGND VGND VPWR VPWR net3385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1501 datamem.data_ram\[20\]\[8\] VGND VGND VPWR VPWR net2651 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2246 rvcpu.dp.rf.reg_file_arr\[1\]\[20\] VGND VGND VPWR VPWR net3396 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1512 rvcpu.dp.rf.reg_file_arr\[28\]\[18\] VGND VGND VPWR VPWR net2662 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2257 datamem.data_ram\[58\]\[24\] VGND VGND VPWR VPWR net3407 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1523 rvcpu.dp.rf.reg_file_arr\[29\]\[18\] VGND VGND VPWR VPWR net2673 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2268 rvcpu.dp.rf.reg_file_arr\[0\]\[7\] VGND VGND VPWR VPWR net3418 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1534 datamem.data_ram\[16\]\[29\] VGND VGND VPWR VPWR net2684 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2279 datamem.data_ram\[8\]\[27\] VGND VGND VPWR VPWR net3429 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1545 datamem.data_ram\[1\]\[22\] VGND VGND VPWR VPWR net2695 sky130_fd_sc_hd__dlygate4sd3_1
X_26650_ _10075_ VGND VGND VPWR VPWR _11672_ sky130_fd_sc_hd__buf_2
Xhold1556 datamem.data_ram\[5\]\[22\] VGND VGND VPWR VPWR net2706 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1567 rvcpu.dp.rf.reg_file_arr\[16\]\[14\] VGND VGND VPWR VPWR net2717 sky130_fd_sc_hd__dlygate4sd3_1
X_23862_ clknet_1_1__leaf__10203_ VGND VGND VPWR VPWR _10220_ sky130_fd_sc_hd__buf_1
Xhold1578 rvcpu.dp.rf.reg_file_arr\[18\]\[28\] VGND VGND VPWR VPWR net2728 sky130_fd_sc_hd__dlygate4sd3_1
X_25601_ _10075_ VGND VGND VPWR VPWR _11064_ sky130_fd_sc_hd__clkbuf_4
Xhold1589 rvcpu.dp.rf.reg_file_arr\[12\]\[6\] VGND VGND VPWR VPWR net2739 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22813_ _09944_ _09948_ _09952_ _09389_ VGND VGND VPWR VPWR _01150_ sky130_fd_sc_hd__o31a_1
X_26581_ _10737_ net2629 _11629_ VGND VGND VPWR VPWR _11636_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_154_Right_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28320_ _12359_ net3800 _12632_ VGND VGND VPWR VPWR _12634_ sky130_fd_sc_hd__mux2_1
Xclkbuf_0__10181_ _10181_ VGND VGND VPWR VPWR clknet_0__10181_ sky130_fd_sc_hd__clkbuf_16
X_25532_ _10729_ net3436 net54 VGND VGND VPWR VPWR _11024_ sky130_fd_sc_hd__mux2_1
X_22744_ _09398_ _09886_ VGND VGND VPWR VPWR _09887_ sky130_fd_sc_hd__or2_1
Xclkbuf_1_1__f__10081_ clknet_0__10081_ VGND VGND VPWR VPWR clknet_1_1__leaf__10081_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_211_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28251_ _12595_ VGND VGND VPWR VPWR _03945_ sky130_fd_sc_hd__clkbuf_1
X_25463_ _10954_ net1536 _10984_ _10987_ VGND VGND VPWR VPWR _02765_ sky130_fd_sc_hd__a31o_1
XFILLER_0_192_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_211_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22675_ _09412_ _09817_ _09819_ _09821_ _09525_ VGND VGND VPWR VPWR _09822_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_192_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27202_ _11970_ _12008_ VGND VGND VPWR VPWR _12011_ sky130_fd_sc_hd__and2_1
X_24414_ _10387_ VGND VGND VPWR VPWR _02316_ sky130_fd_sc_hd__clkbuf_1
X_28182_ _12558_ VGND VGND VPWR VPWR _03913_ sky130_fd_sc_hd__clkbuf_1
X_21626_ _08532_ _08873_ _08875_ _08699_ VGND VGND VPWR VPWR _08876_ sky130_fd_sc_hd__a211o_1
X_25394_ _10938_ net1533 _10949_ _10951_ VGND VGND VPWR VPWR _02732_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_205_Left_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_180_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27133_ _11956_ net1451 _11964_ _11967_ VGND VGND VPWR VPWR _03455_ sky130_fd_sc_hd__a31o_1
XFILLER_0_191_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24345_ _09273_ net3916 _10348_ VGND VGND VPWR VPWR _10350_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21557_ _08628_ VGND VGND VPWR VPWR _08810_ sky130_fd_sc_hd__buf_4
XFILLER_0_168_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27064_ _11822_ _11924_ VGND VGND VPWR VPWR _11925_ sky130_fd_sc_hd__and2_1
X_20508_ datamem.data_ram\[54\]\[21\] _06630_ _06665_ datamem.data_ram\[53\]\[21\]
+ VGND VGND VPWR VPWR _07799_ sky130_fd_sc_hd__o22a_1
XFILLER_0_90_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24276_ _09244_ net4298 _10307_ VGND VGND VPWR VPWR _10311_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_1275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21488_ _08740_ _08741_ _08743_ VGND VGND VPWR VPWR _08744_ sky130_fd_sc_hd__mux2_2
XFILLER_0_43_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26015_ net21 _11152_ VGND VGND VPWR VPWR _11333_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20439_ datamem.data_ram\[29\]\[12\] _06721_ _06654_ datamem.data_ram\[25\]\[12\]
+ VGND VGND VPWR VPWR _07731_ sky130_fd_sc_hd__o22a_1
XFILLER_0_120_437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_224_5864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22109_ _09318_ net2860 _09302_ VGND VGND VPWR VPWR _09319_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_224_5875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15980_ _14327_ VGND VGND VPWR VPWR _02037_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_214_Left_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27966_ _12437_ net3589 _12431_ VGND VGND VPWR VPWR _12438_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14931_ _13329_ _13422_ VGND VGND VPWR VPWR _13480_ sky130_fd_sc_hd__or2_1
X_29705_ net1051 _01440_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[22\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_209_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26917_ _11835_ _11823_ VGND VGND VPWR VPWR _11836_ sky130_fd_sc_hd__and2_1
X_27897_ _12391_ net1677 _12393_ _12399_ VGND VGND VPWR VPWR _03787_ sky130_fd_sc_hd__a31o_1
XFILLER_0_76_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2780 datamem.data_ram\[46\]\[18\] VGND VGND VPWR VPWR net3930 sky130_fd_sc_hd__dlygate4sd3_1
X_14862_ rvcpu.dp.pcreg.q\[4\] rvcpu.dp.pcreg.q\[3\] VGND VGND VPWR VPWR _13414_ sky130_fd_sc_hd__nand2_8
Xhold2791 datamem.data_ram\[26\]\[16\] VGND VGND VPWR VPWR net3941 sky130_fd_sc_hd__dlygate4sd3_1
X_29636_ clknet_leaf_146_clk _01371_ VGND VGND VPWR VPWR datamem.data_ram\[5\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_17650_ net1953 _13225_ _05093_ VGND VGND VPWR VPWR _05098_ sky130_fd_sc_hd__mux2_1
X_26848_ _11687_ _11786_ VGND VGND VPWR VPWR _11792_ sky130_fd_sc_hd__and2_1
XFILLER_0_215_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16601_ _14133_ net4071 _04540_ VGND VGND VPWR VPWR _04542_ sky130_fd_sc_hd__mux2_1
X_17581_ _05061_ VGND VGND VPWR VPWR _01246_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26779_ _11679_ _11749_ VGND VGND VPWR VPWR _11751_ sky130_fd_sc_hd__and2_1
X_14793_ _13345_ VGND VGND VPWR VPWR _13346_ sky130_fd_sc_hd__clkbuf_4
X_29567_ net921 _01302_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[26\]\[2\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_121_Right_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19320_ _06605_ _06615_ VGND VGND VPWR VPWR _06616_ sky130_fd_sc_hd__nand2_4
X_16532_ _14133_ net3687 _04503_ VGND VGND VPWR VPWR _04505_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24134__639 clknet_1_1__leaf__10261_ VGND VGND VPWR VPWR net765 sky130_fd_sc_hd__inv_2
XFILLER_0_168_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28518_ _09287_ VGND VGND VPWR VPWR _12747_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_80_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29498_ net860 _01233_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[28\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19251_ rvcpu.dp.plde.ImmExtE\[30\] rvcpu.dp.plde.PCE\[30\] VGND VGND VPWR VPWR _06554_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16463_ _04468_ VGND VGND VPWR VPWR _01811_ sky130_fd_sc_hd__clkbuf_1
X_28449_ _12706_ VGND VGND VPWR VPWR _04032_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_223_Left_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_175_4694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15414_ _13309_ _13809_ _13428_ VGND VGND VPWR VPWR _13946_ sky130_fd_sc_hd__o21ai_1
X_18202_ _05566_ _05509_ VGND VGND VPWR VPWR _05567_ sky130_fd_sc_hd__or2_1
XFILLER_0_155_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19182_ _06494_ VGND VGND VPWR VPWR rvcpu.dp.lAuiPCE\[20\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31460_ clknet_leaf_76_clk rvcpu.dp.SrcBFW_Mux.y\[18\] VGND VGND VPWR VPWR rvcpu.dp.plem.WriteDataM\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_117_3310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16394_ net2950 _14424_ _14561_ VGND VGND VPWR VPWR _14563_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18133_ rvcpu.dp.plem.ALUResultM\[17\] _05339_ _05340_ _13225_ VGND VGND VPWR VPWR
+ _05499_ sky130_fd_sc_hd__o22a_1
X_23590__211 clknet_1_1__leaf__10177_ VGND VGND VPWR VPWR net337 sky130_fd_sc_hd__inv_2
X_30411_ net749 _02146_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[31\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_15345_ _13332_ _13307_ _13350_ _13314_ VGND VGND VPWR VPWR _13881_ sky130_fd_sc_hd__a211o_1
XFILLER_0_155_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31391_ clknet_leaf_40_clk _03094_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCE\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_3218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18064_ _05410_ _05419_ _05427_ _05431_ VGND VGND VPWR VPWR _05432_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_78_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30342_ net688 _02077_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[4\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_15276_ _13806_ _13808_ _13810_ _13814_ VGND VGND VPWR VPWR _13815_ sky130_fd_sc_hd__o31a_1
XFILLER_0_112_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold108 rvcpu.dp.plem.ALUResultM\[10\] VGND VGND VPWR VPWR net1258 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_184_4908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17015_ _04761_ VGND VGND VPWR VPWR _01528_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_184_4919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold119 rvcpu.dp.plde.funct3E\[0\] VGND VGND VPWR VPWR net1269 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30273_ net627 _02008_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[6\]\[28\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_74_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32012_ clknet_leaf_128_clk _03434_ VGND VGND VPWR VPWR datamem.data_ram\[27\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18966_ _05661_ _06059_ _06302_ _05733_ VGND VGND VPWR VPWR _06303_ sky130_fd_sc_hd__a22o_1
X_23707__301 clknet_1_0__leaf__10196_ VGND VGND VPWR VPWR net427 sky130_fd_sc_hd__inv_2
XFILLER_0_225_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17917_ _05288_ _05289_ VGND VGND VPWR VPWR _05290_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_143_3926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_225_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18897_ _05467_ _06225_ _05466_ VGND VGND VPWR VPWR _06238_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_143_3937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32914_ clknet_leaf_156_clk _04336_ VGND VGND VPWR VPWR datamem.data_ram\[0\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_33_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17848_ rvcpu.dp.plem.ALUResultM\[13\] _05177_ VGND VGND VPWR VPWR _05227_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_33_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32845_ clknet_leaf_96_clk _04267_ VGND VGND VPWR VPWR datamem.data_ram\[7\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_17779_ _05176_ VGND VGND VPWR VPWR _05177_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19518_ datamem.data_ram\[63\]\[24\] _06670_ _06781_ datamem.data_ram\[57\]\[24\]
+ _06813_ VGND VGND VPWR VPWR _06814_ sky130_fd_sc_hd__o221a_1
XFILLER_0_159_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20790_ datamem.data_ram\[22\]\[30\] _06629_ _06703_ datamem.data_ram\[21\]\[30\]
+ VGND VGND VPWR VPWR _08080_ sky130_fd_sc_hd__o22a_1
X_32776_ clknet_leaf_185_clk _04198_ VGND VGND VPWR VPWR datamem.data_ram\[14\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_102_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_102_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19449_ datamem.data_ram\[46\]\[16\] _06744_ _06695_ datamem.data_ram\[40\]\[16\]
+ VGND VGND VPWR VPWR _06745_ sky130_fd_sc_hd__o22a_1
X_31727_ net176 _03185_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[9\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22460_ rvcpu.dp.rf.reg_file_arr\[16\]\[8\] rvcpu.dp.rf.reg_file_arr\[17\]\[8\] rvcpu.dp.rf.reg_file_arr\[18\]\[8\]
+ rvcpu.dp.rf.reg_file_arr\[19\]\[8\] _09406_ _09408_ VGND VGND VPWR VPWR _09618_
+ sky130_fd_sc_hd__mux4_1
X_31658_ clknet_leaf_64_clk net1887 VGND VGND VPWR VPWR rvcpu.dp.plmw.ALUResultW\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_23753__343 clknet_1_0__leaf__10200_ VGND VGND VPWR VPWR net469 sky130_fd_sc_hd__inv_2
XFILLER_0_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_518 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21411_ _08565_ _08668_ _08670_ _08576_ VGND VGND VPWR VPWR _08671_ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30609_ clknet_leaf_218_clk _02344_ VGND VGND VPWR VPWR datamem.data_ram\[52\]\[28\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22391_ rvcpu.dp.rf.reg_file_arr\[12\]\[4\] rvcpu.dp.rf.reg_file_arr\[13\]\[4\] rvcpu.dp.rf.reg_file_arr\[14\]\[4\]
+ rvcpu.dp.rf.reg_file_arr\[15\]\[4\] _09552_ _09382_ VGND VGND VPWR VPWR _09553_
+ sky130_fd_sc_hd__mux4_1
X_31589_ clknet_leaf_57_clk net1247 VGND VGND VPWR VPWR rvcpu.dp.plmw.PCPlus4W\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21342_ rvcpu.ALUResultE\[11\] rvcpu.ALUResultE\[13\] VGND VGND VPWR VPWR _08604_
+ sky130_fd_sc_hd__or2_1
X_23868__430 clknet_1_1__leaf__10220_ VGND VGND VPWR VPWR net556 sky130_fd_sc_hd__inv_2
XFILLER_0_60_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold620 rvcpu.dp.plfd.PCPlus4D\[28\] VGND VGND VPWR VPWR net1770 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21273_ rvcpu.dp.plfd.InstrD\[15\] VGND VGND VPWR VPWR _08535_ sky130_fd_sc_hd__buf_4
Xhold631 datamem.data_ram\[19\]\[5\] VGND VGND VPWR VPWR net1781 sky130_fd_sc_hd__dlygate4sd3_1
Xhold642 datamem.data_ram\[58\]\[5\] VGND VGND VPWR VPWR net1792 sky130_fd_sc_hd__dlygate4sd3_1
Xhold653 rvcpu.dp.plfd.PCD\[15\] VGND VGND VPWR VPWR net1803 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20224_ datamem.data_ram\[21\]\[3\] _07132_ _07513_ _07516_ VGND VGND VPWR VPWR _07517_
+ sky130_fd_sc_hd__a211o_1
Xhold664 datamem.data_ram\[35\]\[2\] VGND VGND VPWR VPWR net1814 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold675 datamem.data_ram\[5\]\[0\] VGND VGND VPWR VPWR net1825 sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 datamem.data_ram\[52\]\[4\] VGND VGND VPWR VPWR net1836 sky130_fd_sc_hd__dlygate4sd3_1
Xhold697 rvcpu.dp.plfd.PCD\[25\] VGND VGND VPWR VPWR net1847 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_223_Right_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20155_ _06751_ _07442_ _07447_ VGND VGND VPWR VPWR _07448_ sky130_fd_sc_hd__or3_1
X_27820_ _12155_ net3893 net78 VGND VGND VPWR VPWR _12353_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2010 datamem.data_ram\[49\]\[14\] VGND VGND VPWR VPWR net3160 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2021 datamem.data_ram\[31\]\[12\] VGND VGND VPWR VPWR net3171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2032 datamem.data_ram\[11\]\[26\] VGND VGND VPWR VPWR net3182 sky130_fd_sc_hd__dlygate4sd3_1
X_27751_ _12140_ net1936 _12307_ VGND VGND VPWR VPWR _12315_ sky130_fd_sc_hd__mux2_1
Xhold2043 datamem.data_ram\[20\]\[12\] VGND VGND VPWR VPWR net3193 sky130_fd_sc_hd__dlygate4sd3_1
X_24963_ _10394_ net3966 _10696_ VGND VGND VPWR VPWR _10701_ sky130_fd_sc_hd__mux2_1
X_20086_ datamem.data_ram\[54\]\[10\] _06626_ _06811_ datamem.data_ram\[48\]\[10\]
+ VGND VGND VPWR VPWR _07380_ sky130_fd_sc_hd__o22a_1
Xhold2054 rvcpu.dp.rf.reg_file_arr\[22\]\[0\] VGND VGND VPWR VPWR net3204 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_96_clk clknet_5_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_96_clk sky130_fd_sc_hd__clkbuf_8
Xhold2065 rvcpu.dp.rf.reg_file_arr\[4\]\[29\] VGND VGND VPWR VPWR net3215 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1320 datamem.data_ram\[42\]\[30\] VGND VGND VPWR VPWR net2470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1331 datamem.data_ram\[35\]\[30\] VGND VGND VPWR VPWR net2481 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2076 datamem.data_ram\[23\]\[24\] VGND VGND VPWR VPWR net3226 sky130_fd_sc_hd__dlygate4sd3_1
X_26702_ _10814_ net3246 _11704_ VGND VGND VPWR VPWR _11706_ sky130_fd_sc_hd__mux2_1
XFILLER_0_225_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2087 datamem.data_ram\[15\]\[24\] VGND VGND VPWR VPWR net3237 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1342 datamem.data_ram\[32\]\[8\] VGND VGND VPWR VPWR net2492 sky130_fd_sc_hd__dlygate4sd3_1
X_27682_ _12095_ net2139 net51 VGND VGND VPWR VPWR _12278_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24894_ _10448_ net3749 _10659_ VGND VGND VPWR VPWR _10664_ sky130_fd_sc_hd__mux2_1
Xhold2098 datamem.data_ram\[46\]\[25\] VGND VGND VPWR VPWR net3248 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1353 datamem.data_ram\[2\]\[28\] VGND VGND VPWR VPWR net2503 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1364 rvcpu.dp.rf.reg_file_arr\[18\]\[25\] VGND VGND VPWR VPWR net2514 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1375 rvcpu.dp.rf.reg_file_arr\[30\]\[8\] VGND VGND VPWR VPWR net2525 sky130_fd_sc_hd__dlygate4sd3_1
X_26633_ _11661_ VGND VGND VPWR VPWR _11662_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_196_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29421_ clknet_leaf_98_clk _01156_ VGND VGND VPWR VPWR datamem.data_ram\[5\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1386 rvcpu.dp.rf.reg_file_arr\[13\]\[18\] VGND VGND VPWR VPWR net2536 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f__10202_ clknet_0__10202_ VGND VGND VPWR VPWR clknet_1_1__leaf__10202_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_212_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_504 _11681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1397 rvcpu.dp.rf.reg_file_arr\[6\]\[24\] VGND VGND VPWR VPWR net2547 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_515 _13223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_526 _13272_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_197_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_196_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_537 rvcpu.dp.plmw.ReadDataW\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29352_ clknet_leaf_144_clk _01087_ VGND VGND VPWR VPWR datamem.data_ram\[61\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__10133_ clknet_0__10133_ VGND VGND VPWR VPWR clknet_1_1__leaf__10133_
+ sky130_fd_sc_hd__clkbuf_16
X_26564_ _10824_ net3060 _11620_ VGND VGND VPWR VPWR _11627_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_548 _06780_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_170_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20988_ datamem.data_ram\[4\]\[15\] datamem.data_ram\[5\]\[15\] _06652_ VGND VGND
+ VPWR VPWR _08277_ sky130_fd_sc_hd__mux2_1
XANTENNA_559 _08986_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_211_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25515_ _10413_ _11010_ VGND VGND VPWR VPWR _11014_ sky130_fd_sc_hd__and2_1
X_28303_ _12450_ net3581 net72 VGND VGND VPWR VPWR _12625_ sky130_fd_sc_hd__mux2_1
X_29283_ _09313_ net2341 _13159_ VGND VGND VPWR VPWR _13163_ sky130_fd_sc_hd__mux2_1
X_22727_ rvcpu.dp.rf.reg_file_arr\[28\]\[22\] rvcpu.dp.rf.reg_file_arr\[30\]\[22\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[22\] rvcpu.dp.rf.reg_file_arr\[31\]\[22\] _09443_
+ _09453_ VGND VGND VPWR VPWR _09871_ sky130_fd_sc_hd__mux4_1
XFILLER_0_149_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28234_ _12586_ VGND VGND VPWR VPWR _03937_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25446_ _10979_ _10051_ VGND VGND VPWR VPWR _10980_ sky130_fd_sc_hd__nand2_4
X_23081__762 clknet_1_1__leaf__10091_ VGND VGND VPWR VPWR net888 sky130_fd_sc_hd__inv_2
XFILLER_0_48_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_188_5008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22658_ rvcpu.dp.rf.reg_file_arr\[0\]\[18\] rvcpu.dp.rf.reg_file_arr\[1\]\[18\] rvcpu.dp.rf.reg_file_arr\[2\]\[18\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[18\] _09714_ _09585_ VGND VGND VPWR VPWR _09806_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_188_5019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_213_5598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28165_ _12549_ VGND VGND VPWR VPWR _03905_ sky130_fd_sc_hd__clkbuf_1
X_21609_ rvcpu.dp.rf.reg_file_arr\[8\]\[11\] rvcpu.dp.rf.reg_file_arr\[10\]\[11\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[11\] rvcpu.dp.rf.reg_file_arr\[11\]\[11\] _08693_
+ _08818_ VGND VGND VPWR VPWR _08860_ sky130_fd_sc_hd__mux4_1
X_23003__708 clknet_1_1__leaf__10085_ VGND VGND VPWR VPWR net834 sky130_fd_sc_hd__inv_2
XFILLER_0_91_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25377_ _10938_ net1573 _10934_ _10940_ VGND VGND VPWR VPWR _02726_ sky130_fd_sc_hd__a31o_1
XFILLER_0_192_495 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_4580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22589_ _09482_ _09740_ VGND VGND VPWR VPWR _09741_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_20_clk clknet_5_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_20_clk sky130_fd_sc_hd__clkbuf_8
X_27116_ _11827_ _11953_ VGND VGND VPWR VPWR _11957_ sky130_fd_sc_hd__and2_1
X_15130_ _13674_ VGND VGND VPWR VPWR _13675_ sky130_fd_sc_hd__inv_2
X_24328_ _10340_ VGND VGND VPWR VPWR _02277_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28096_ _12452_ net3807 net75 VGND VGND VPWR VPWR _12513_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_226_5915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15061_ rvcpu.dp.pcreg.q\[8\] _13513_ VGND VGND VPWR VPWR _13608_ sky130_fd_sc_hd__nor2_2
X_27047_ _11827_ _11911_ VGND VGND VPWR VPWR _11914_ sky130_fd_sc_hd__and2_1
X_24259_ _09314_ net3963 _10298_ VGND VGND VPWR VPWR _10302_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_226_5926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_147_4015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_147_4026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18820_ _05497_ _05516_ _06165_ VGND VGND VPWR VPWR _06166_ sky130_fd_sc_hd__or3_1
XFILLER_0_207_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28998_ _13008_ VGND VGND VPWR VPWR _13009_ sky130_fd_sc_hd__clkbuf_2
X_18751_ _06077_ _06096_ _06101_ VGND VGND VPWR VPWR _06102_ sky130_fd_sc_hd__o21ai_1
X_27949_ _12367_ net4200 _12421_ VGND VGND VPWR VPWR _12427_ sky130_fd_sc_hd__mux2_1
X_15963_ _14318_ VGND VGND VPWR VPWR _02045_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_87_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_87_clk sky130_fd_sc_hd__clkbuf_8
X_23923__479 clknet_1_1__leaf__10226_ VGND VGND VPWR VPWR net605 sky130_fd_sc_hd__inv_2
X_17702_ _05125_ VGND VGND VPWR VPWR _01189_ sky130_fd_sc_hd__clkbuf_1
X_14914_ _13379_ _13462_ _13463_ VGND VGND VPWR VPWR _13464_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_106_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18682_ _05427_ _05406_ _05431_ _05445_ VGND VGND VPWR VPWR _06036_ sky130_fd_sc_hd__a31o_1
X_30960_ clknet_leaf_163_clk _02695_ VGND VGND VPWR VPWR datamem.data_ram\[3\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_15894_ net2735 _13201_ _14275_ VGND VGND VPWR VPWR _14282_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_106_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17633_ net2207 _13200_ _05082_ VGND VGND VPWR VPWR _05089_ sky130_fd_sc_hd__mux2_1
X_29619_ net973 _01354_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[25\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_14845_ _13331_ _13397_ VGND VGND VPWR VPWR _13398_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_177_4734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_177_4745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1138 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30891_ clknet_leaf_193_clk _02626_ VGND VGND VPWR VPWR datamem.data_ram\[42\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32630_ clknet_leaf_93_clk _04052_ VGND VGND VPWR VPWR datamem.data_ram\[1\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_14776_ _13296_ _13300_ VGND VGND VPWR VPWR _13329_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17564_ _05052_ VGND VGND VPWR VPWR _01254_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_67_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19303_ _06598_ VGND VGND VPWR VPWR _06599_ sky130_fd_sc_hd__buf_6
XFILLER_0_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16515_ _04495_ VGND VGND VPWR VPWR _01786_ sky130_fd_sc_hd__clkbuf_1
X_32561_ clknet_leaf_79_clk _03983_ VGND VGND VPWR VPWR datamem.data_ram\[22\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_17495_ _13198_ net4048 _05010_ VGND VGND VPWR VPWR _05016_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31512_ clknet_leaf_57_clk net1250 VGND VGND VPWR VPWR rvcpu.dp.plem.PCPlus4M\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_19234_ _06539_ VGND VGND VPWR VPWR rvcpu.dp.lAuiPCE\[27\] sky130_fd_sc_hd__clkbuf_1
X_16446_ net2088 _14476_ _04451_ VGND VGND VPWR VPWR _04458_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32492_ clknet_leaf_169_clk _03914_ VGND VGND VPWR VPWR datamem.data_ram\[25\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_23279__924 clknet_1_1__leaf__10129_ VGND VGND VPWR VPWR net1050 sky130_fd_sc_hd__inv_2
XFILLER_0_2_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_3752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_3763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19165_ _06479_ VGND VGND VPWR VPWR rvcpu.dp.lAuiPCE\[18\] sky130_fd_sc_hd__clkbuf_1
X_31443_ clknet_leaf_6_clk rvcpu.dp.SrcBFW_Mux.y\[1\] VGND VGND VPWR VPWR rvcpu.dp.plem.WriteDataM\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_6_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16377_ _14553_ VGND VGND VPWR VPWR _01850_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_11_clk clknet_5_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15328_ _13615_ _13472_ VGND VGND VPWR VPWR _13865_ sky130_fd_sc_hd__nand2_1
XFILLER_0_205_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18116_ rvcpu.dp.plem.ALUResultM\[19\] _05339_ _05340_ _13219_ VGND VGND VPWR VPWR
+ _05483_ sky130_fd_sc_hd__o22a_1
XFILLER_0_121_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31374_ clknet_leaf_18_clk _03077_ VGND VGND VPWR VPWR rvcpu.dp.plde.ImmExtE\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19096_ rvcpu.dp.plde.luiE VGND VGND VPWR VPWR _06419_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_0__f__10222_ clknet_0__10222_ VGND VGND VPWR VPWR clknet_1_0__leaf__10222_
+ sky130_fd_sc_hd__clkbuf_16
X_30325_ net671 _02060_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[4\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_15259_ _13675_ _13776_ _13798_ _13441_ VGND VGND VPWR VPWR _13799_ sky130_fd_sc_hd__a31o_1
X_18047_ _05412_ _05415_ VGND VGND VPWR VPWR _05416_ sky130_fd_sc_hd__and2_1
XFILLER_0_151_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__10153_ clknet_0__10153_ VGND VGND VPWR VPWR clknet_1_0__leaf__10153_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_112_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30256_ net610 _01991_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[6\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__10084_ clknet_0__10084_ VGND VGND VPWR VPWR clknet_1_0__leaf__10084_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30187_ net541 _01922_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[8\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_19998_ datamem.data_ram\[19\]\[2\] _06942_ _07288_ _07291_ VGND VGND VPWR VPWR _07292_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_201_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23783__369 clknet_1_0__leaf__10204_ VGND VGND VPWR VPWR net495 sky130_fd_sc_hd__inv_2
XFILLER_0_226_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18949_ _05549_ _05727_ _06108_ _05547_ _06286_ VGND VGND VPWR VPWR _06287_ sky130_fd_sc_hd__a221o_1
X_23251__898 clknet_1_1__leaf__10127_ VGND VGND VPWR VPWR net1024 sky130_fd_sc_hd__inv_2
XFILLER_0_226_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_78_clk clknet_5_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_78_clk sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_129_Left_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21960_ _08541_ _09191_ VGND VGND VPWR VPWR _09192_ sky130_fd_sc_hd__and2_1
XFILLER_0_207_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20911_ datamem.data_ram\[18\]\[22\] datamem.data_ram\[19\]\[22\] _07836_ VGND VGND
+ VPWR VPWR _08201_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21891_ rvcpu.dp.rf.reg_file_arr\[16\]\[27\] rvcpu.dp.rf.reg_file_arr\[17\]\[27\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[27\] rvcpu.dp.rf.reg_file_arr\[19\]\[27\] _08799_
+ _08800_ VGND VGND VPWR VPWR _09126_ sky130_fd_sc_hd__mux4_1
XFILLER_0_90_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20842_ _08124_ _07177_ VGND VGND VPWR VPWR _08132_ sky130_fd_sc_hd__or2_1
X_32828_ clknet_leaf_162_clk _04250_ VGND VGND VPWR VPWR datamem.data_ram\[12\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_23597__217 clknet_1_0__leaf__10178_ VGND VGND VPWR VPWR net343 sky130_fd_sc_hd__inv_2
XFILLER_0_89_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_221_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23561_ clknet_1_1__leaf__10172_ VGND VGND VPWR VPWR _10175_ sky130_fd_sc_hd__buf_1
X_20773_ _07822_ _08060_ _08062_ _07868_ VGND VGND VPWR VPWR _08063_ sky130_fd_sc_hd__o211a_1
X_32759_ clknet_leaf_157_clk _04181_ VGND VGND VPWR VPWR datamem.data_ram\[15\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25300_ _10762_ net2205 _10887_ VGND VGND VPWR VPWR _10893_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23677__274 clknet_1_1__leaf__10193_ VGND VGND VPWR VPWR net400 sky130_fd_sc_hd__inv_2
X_22512_ rvcpu.dp.rf.reg_file_arr\[0\]\[10\] rvcpu.dp.rf.reg_file_arr\[1\]\[10\] rvcpu.dp.rf.reg_file_arr\[2\]\[10\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[10\] _09477_ _09466_ VGND VGND VPWR VPWR _09668_
+ sky130_fd_sc_hd__mux4_1
X_26280_ _11472_ VGND VGND VPWR VPWR _03097_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_174_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25231_ _10764_ net2259 _10848_ VGND VGND VPWR VPWR _10855_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_138_Left_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22443_ _09596_ _09598_ _09601_ _09412_ _09413_ VGND VGND VPWR VPWR _09602_ sky130_fd_sc_hd__a221o_1
XFILLER_0_134_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25162_ _10814_ net3050 net58 VGND VGND VPWR VPWR _10815_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22374_ _09429_ _09533_ _09536_ _09438_ VGND VGND VPWR VPWR _09537_ sky130_fd_sc_hd__a211o_1
XFILLER_0_115_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21325_ _08581_ rvcpu.dp.plde.RdE\[1\] rvcpu.dp.plde.RdE\[4\] _08509_ _08586_ VGND
+ VGND VPWR VPWR _08587_ sky130_fd_sc_hd__o221a_1
X_25093_ _10600_ _10778_ VGND VGND VPWR VPWR _10779_ sky130_fd_sc_hd__nor2_2
XFILLER_0_32_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29970_ net340 _01705_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[15\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_206_1278 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28921_ _12700_ net2698 _12959_ VGND VGND VPWR VPWR _12966_ sky130_fd_sc_hd__mux2_1
Xhold450 datamem.data_ram\[23\]\[2\] VGND VGND VPWR VPWR net1600 sky130_fd_sc_hd__dlygate4sd3_1
X_21256_ rvcpu.dp.plfd.InstrD\[16\] VGND VGND VPWR VPWR _08518_ sky130_fd_sc_hd__buf_4
Xhold461 datamem.data_ram\[23\]\[5\] VGND VGND VPWR VPWR net1611 sky130_fd_sc_hd__dlygate4sd3_1
Xhold472 datamem.data_ram\[6\]\[2\] VGND VGND VPWR VPWR net1622 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold483 datamem.data_ram\[63\]\[0\] VGND VGND VPWR VPWR net1633 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_221_5801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20207_ datamem.data_ram\[53\]\[11\] _06722_ _06695_ datamem.data_ram\[48\]\[11\]
+ _07499_ VGND VGND VPWR VPWR _07500_ sky130_fd_sc_hd__o221a_1
Xhold494 datamem.data_ram\[63\]\[7\] VGND VGND VPWR VPWR net1644 sky130_fd_sc_hd__dlygate4sd3_1
X_28852_ _12929_ VGND VGND VPWR VPWR _04212_ sky130_fd_sc_hd__clkbuf_1
X_21187_ _08473_ VGND VGND VPWR VPWR _04445_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_216_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_1243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27803_ _12343_ VGND VGND VPWR VPWR _03749_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_147_Left_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20138_ datamem.data_ram\[33\]\[27\] _06782_ _07427_ _07430_ VGND VGND VPWR VPWR
+ _07431_ sky130_fd_sc_hd__o211a_1
XFILLER_0_216_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25995_ net11 _11317_ VGND VGND VPWR VPWR _11322_ sky130_fd_sc_hd__or2_1
X_28783_ _12762_ net3224 _12887_ VGND VGND VPWR VPWR _12893_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_69_clk clknet_5_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_69_clk sky130_fd_sc_hd__clkbuf_8
X_23310__951 clknet_1_0__leaf__10133_ VGND VGND VPWR VPWR net1077 sky130_fd_sc_hd__inv_2
X_24946_ _10448_ net2973 _10687_ VGND VGND VPWR VPWR _10692_ sky130_fd_sc_hd__mux2_1
X_20069_ datamem.data_ram\[55\]\[26\] _06704_ _07242_ datamem.data_ram\[49\]\[26\]
+ _07362_ VGND VGND VPWR VPWR _07363_ sky130_fd_sc_hd__o221a_1
X_27734_ _12095_ net1960 net49 VGND VGND VPWR VPWR _12306_ sky130_fd_sc_hd__mux2_1
Xhold1150 datamem.data_ram\[61\]\[25\] VGND VGND VPWR VPWR net2300 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1161 datamem.data_ram\[54\]\[10\] VGND VGND VPWR VPWR net2311 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1172 datamem.data_ram\[36\]\[19\] VGND VGND VPWR VPWR net2322 sky130_fd_sc_hd__dlygate4sd3_1
X_24877_ _10474_ net2721 net92 VGND VGND VPWR VPWR _10655_ sky130_fd_sc_hd__mux2_1
X_27665_ _12157_ net2519 net79 VGND VGND VPWR VPWR _12269_ sky130_fd_sc_hd__mux2_1
Xhold1183 datamem.data_ram\[39\]\[15\] VGND VGND VPWR VPWR net2333 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_301 _13931_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1194 datamem.data_ram\[16\]\[22\] VGND VGND VPWR VPWR net2344 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_219_5741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_219_5752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29404_ clknet_leaf_0_clk _01139_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD2E\[15\] sky130_fd_sc_hd__dfxtp_1
X_14630_ _13206_ VGND VGND VPWR VPWR _13207_ sky130_fd_sc_hd__buf_4
XANTENNA_312 _14177_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_219_5763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_212_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23828_ _10209_ _09301_ _09361_ VGND VGND VPWR VPWR _10210_ sky130_fd_sc_hd__a21oi_4
XANTENNA_323 _14447_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26616_ _10822_ net2630 _11650_ VGND VGND VPWR VPWR _11656_ sky130_fd_sc_hd__mux2_1
X_27596_ _12140_ net2256 _12224_ VGND VGND VPWR VPWR _12232_ sky130_fd_sc_hd__mux2_1
XANTENNA_334 _14459_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_200_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_345 _14478_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_185_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_356 rvcpu.dp.SrcBFW_Mux.y\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26547_ _11517_ net1833 _11608_ _11617_ VGND VGND VPWR VPWR _03219_ sky130_fd_sc_hd__a31o_1
XANTENNA_367 rvcpu.dp.plde.ImmExtE\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29335_ clknet_leaf_266_clk _01070_ VGND VGND VPWR VPWR datamem.data_ram\[62\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_215_5649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_172_4620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_378 rvcpu.dp.plmw.ReadDataW\[29\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_389 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_4631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_156_Left_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16300_ net4339 _14466_ _14511_ VGND VGND VPWR VPWR _14513_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17280_ _04901_ VGND VGND VPWR VPWR _04902_ sky130_fd_sc_hd__clkbuf_4
X_26478_ _08620_ _08621_ _06562_ VGND VGND VPWR VPWR _11597_ sky130_fd_sc_hd__a21o_1
X_29266_ _09278_ net3625 _13150_ VGND VGND VPWR VPWR _13154_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16231_ net2295 _14472_ _14464_ VGND VGND VPWR VPWR _14473_ sky130_fd_sc_hd__mux2_1
X_25429_ _10751_ net3646 _10970_ VGND VGND VPWR VPWR _10971_ sky130_fd_sc_hd__mux2_1
X_28217_ _12577_ VGND VGND VPWR VPWR _03929_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__10078_ _10078_ VGND VGND VPWR VPWR clknet_0__10078_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_180_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29197_ _13116_ VGND VGND VPWR VPWR _04370_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_183_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload309 clknet_1_1__leaf__10194_ VGND VGND VPWR VPWR clkload309/Y sky130_fd_sc_hd__clkinvlp_4
X_16162_ _13186_ VGND VGND VPWR VPWR _14426_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_134_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28148_ _12540_ VGND VGND VPWR VPWR _03897_ sky130_fd_sc_hd__clkbuf_1
Xclkload17 clknet_5_21__leaf_clk VGND VGND VPWR VPWR clkload17/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload28 clknet_leaf_16_clk VGND VGND VPWR VPWR clkload28/Y sky130_fd_sc_hd__inv_6
X_15113_ _13282_ _13305_ VGND VGND VPWR VPWR _13658_ sky130_fd_sc_hd__and2b_1
Xclkload39 clknet_leaf_23_clk VGND VGND VPWR VPWR clkload39/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_140_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28079_ _12435_ net3836 _12501_ VGND VGND VPWR VPWR _12504_ sky130_fd_sc_hd__mux2_1
X_16093_ _14388_ VGND VGND VPWR VPWR _01977_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30110_ net472 _01845_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[10\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_71_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15044_ _13374_ _13416_ _13465_ _13590_ VGND VGND VPWR VPWR _13591_ sky130_fd_sc_hd__or4_1
X_19921_ datamem.data_ram\[62\]\[17\] _06682_ _06790_ datamem.data_ram\[57\]\[17\]
+ _06810_ VGND VGND VPWR VPWR _07216_ sky130_fd_sc_hd__o221a_1
X_31090_ clknet_leaf_101_clk _02825_ VGND VGND VPWR VPWR datamem.data_ram\[21\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_166_4468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_4479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_165_Left_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30041_ net403 _01776_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[13\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_19852_ datamem.data_ram\[62\]\[1\] _07127_ _06970_ datamem.data_ram\[61\]\[1\] VGND
+ VGND VPWR VPWR _07147_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18803_ _06132_ _06133_ _06150_ VGND VGND VPWR VPWR rvcpu.ALUResultE\[16\] sky130_fd_sc_hd__o21ai_2
XFILLER_0_78_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_5_6__f_clk clknet_2_0_0_clk VGND VGND VPWR VPWR clknet_5_6__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_19783_ datamem.data_ram\[44\]\[9\] _06688_ _06701_ datamem.data_ram\[41\]\[9\] VGND
+ VGND VPWR VPWR _07078_ sky130_fd_sc_hd__o22a_1
XFILLER_0_78_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16995_ net2449 _14478_ _04742_ VGND VGND VPWR VPWR _04750_ sky130_fd_sc_hd__mux2_1
XFILLER_0_223_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18734_ _05324_ _05332_ VGND VGND VPWR VPWR _06085_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_30_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15946_ net2252 _13278_ _14274_ VGND VGND VPWR VPWR _14309_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31992_ clknet_leaf_127_clk _03414_ VGND VGND VPWR VPWR datamem.data_ram\[31\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_0_clk clknet_5_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_69_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_3486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30943_ clknet_leaf_97_clk _02678_ VGND VGND VPWR VPWR datamem.data_ram\[3\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_18665_ _05599_ _05601_ _06017_ _06018_ VGND VGND VPWR VPWR _06020_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_125_3497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23088__768 clknet_1_1__leaf__10102_ VGND VGND VPWR VPWR net894 sky130_fd_sc_hd__inv_2
X_15877_ rvcpu.dp.plmw.RdW\[3\] _13176_ _13174_ VGND VGND VPWR VPWR _14271_ sky130_fd_sc_hd__or3b_4
XFILLER_0_149_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17616_ _05079_ VGND VGND VPWR VPWR _01229_ sky130_fd_sc_hd__clkbuf_1
X_14828_ _13380_ _13369_ VGND VGND VPWR VPWR _13381_ sky130_fd_sc_hd__nor2_2
X_30874_ clknet_leaf_57_clk _02609_ VGND VGND VPWR VPWR datamem.data_ram\[42\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_18596_ _05361_ _05404_ _05356_ VGND VGND VPWR VPWR _05954_ sky130_fd_sc_hd__a21oi_1
X_23819__402 clknet_1_1__leaf__10207_ VGND VGND VPWR VPWR net528 sky130_fd_sc_hd__inv_2
XFILLER_0_153_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32613_ clknet_leaf_78_clk _04035_ VGND VGND VPWR VPWR datamem.data_ram\[20\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_138_3814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17547_ _13275_ net2128 _05009_ VGND VGND VPWR VPWR _05043_ sky130_fd_sc_hd__mux2_1
X_14759_ _13311_ VGND VGND VPWR VPWR _13312_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_15_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32544_ clknet_leaf_171_clk _03966_ VGND VGND VPWR VPWR datamem.data_ram\[23\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_28_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17478_ _05006_ VGND VGND VPWR VPWR _01302_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_229_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19217_ _06521_ _06524_ VGND VGND VPWR VPWR _06525_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_60_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16429_ net2913 _14459_ _14572_ VGND VGND VPWR VPWR _14581_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_99_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32475_ clknet_leaf_247_clk _03897_ VGND VGND VPWR VPWR datamem.data_ram\[26\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_568 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19148_ rvcpu.dp.plde.ImmExtE\[17\] rvcpu.dp.plde.PCE\[17\] VGND VGND VPWR VPWR _06464_
+ sky130_fd_sc_hd__nand2_1
X_31426_ clknet_leaf_59_clk _03129_ VGND VGND VPWR VPWR datamem.data_ram\[44\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19079_ _06402_ _06403_ VGND VGND VPWR VPWR _06404_ sky130_fd_sc_hd__xnor2_1
X_31357_ clknet_leaf_22_clk _03060_ VGND VGND VPWR VPWR rvcpu.dp.plde.ImmExtE\[6\]
+ sky130_fd_sc_hd__dfxtp_2
Xclkbuf_1_0__f__10205_ clknet_0__10205_ VGND VGND VPWR VPWR clknet_1_0__leaf__10205_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_124_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21110_ datamem.data_ram\[22\]\[7\] _06950_ _06919_ datamem.data_ram\[21\]\[7\] _08398_
+ VGND VGND VPWR VPWR _08399_ sky130_fd_sc_hd__a221o_1
XFILLER_0_160_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30308_ net654 _02043_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[5\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22090_ _09303_ VGND VGND VPWR VPWR _01076_ sky130_fd_sc_hd__clkbuf_1
X_31288_ clknet_leaf_109_clk _02991_ VGND VGND VPWR VPWR datamem.data_ram\[34\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f__10136_ clknet_0__10136_ VGND VGND VPWR VPWR clknet_1_0__leaf__10136_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_58_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21041_ datamem.data_ram\[8\]\[31\] _06644_ _08326_ _06917_ _08329_ VGND VGND VPWR
+ VPWR _08330_ sky130_fd_sc_hd__o221a_1
X_30239_ net593 _01974_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[7\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24800_ _10613_ VGND VGND VPWR VPWR _02476_ sky130_fd_sc_hd__clkbuf_1
X_23032__734 clknet_1_1__leaf__10088_ VGND VGND VPWR VPWR net860 sky130_fd_sc_hd__inv_2
XFILLER_0_226_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25780_ net1376 _11144_ _11147_ _11176_ VGND VGND VPWR VPWR _02893_ sky130_fd_sc_hd__o211a_1
X_24731_ _10574_ VGND VGND VPWR VPWR _02446_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21943_ _08842_ _09175_ VGND VGND VPWR VPWR _09176_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27450_ _12152_ VGND VGND VPWR VPWR _03587_ sky130_fd_sc_hd__clkbuf_1
X_24662_ _10412_ net1541 _10531_ _10536_ VGND VGND VPWR VPWR _02415_ sky130_fd_sc_hd__a31o_1
XFILLER_0_132_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21874_ rvcpu.dp.rf.reg_file_arr\[20\]\[26\] rvcpu.dp.rf.reg_file_arr\[21\]\[26\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[26\] rvcpu.dp.rf.reg_file_arr\[23\]\[26\] _08778_
+ _08825_ VGND VGND VPWR VPWR _09110_ sky130_fd_sc_hd__mux4_1
X_26401_ _06398_ _11522_ _11526_ _11164_ _11543_ VGND VGND VPWR VPWR _11544_ sky130_fd_sc_hd__a221o_1
XFILLER_0_210_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27381_ _10729_ net4115 net86 VGND VGND VPWR VPWR _12110_ sky130_fd_sc_hd__mux2_1
X_20825_ datamem.data_ram\[10\]\[30\] datamem.data_ram\[11\]\[30\] _07827_ VGND VGND
+ VPWR VPWR _08115_ sky130_fd_sc_hd__mux2_1
X_24593_ _10497_ VGND VGND VPWR VPWR _02385_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26332_ _11104_ VGND VGND VPWR VPWR _11501_ sky130_fd_sc_hd__buf_2
X_29120_ _13075_ VGND VGND VPWR VPWR _04334_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20756_ datamem.data_ram\[6\]\[6\] datamem.data_ram\[7\]\[6\] _07828_ VGND VGND VPWR
+ VPWR _08046_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29051_ _10075_ _13031_ VGND VGND VPWR VPWR _13039_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_210_5524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26263_ _11463_ VGND VGND VPWR VPWR _03089_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_635 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_210_5535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20687_ datamem.data_ram\[55\]\[5\] _06993_ _07977_ VGND VGND VPWR VPWR _07978_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_210_5546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25214_ _10824_ net3267 _10839_ VGND VGND VPWR VPWR _10846_ sky130_fd_sc_hd__mux2_1
X_28002_ _09290_ VGND VGND VPWR VPWR _12462_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_165_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22426_ rvcpu.dp.rf.reg_file_arr\[0\]\[6\] rvcpu.dp.rf.reg_file_arr\[1\]\[6\] rvcpu.dp.rf.reg_file_arr\[2\]\[6\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[6\] _09417_ _09585_ VGND VGND VPWR VPWR _09586_ sky130_fd_sc_hd__mux4_1
XFILLER_0_208_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26194_ _11434_ VGND VGND VPWR VPWR _03049_ sky130_fd_sc_hd__clkbuf_1
X_25145_ _10756_ net3062 _10802_ VGND VGND VPWR VPWR _10805_ sky130_fd_sc_hd__mux2_1
X_22357_ rvcpu.dp.rf.reg_file_arr\[28\]\[3\] rvcpu.dp.rf.reg_file_arr\[30\]\[3\] rvcpu.dp.rf.reg_file_arr\[29\]\[3\]
+ rvcpu.dp.rf.reg_file_arr\[31\]\[3\] _09446_ _09402_ VGND VGND VPWR VPWR _09520_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_5_590 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21308_ _08569_ VGND VGND VPWR VPWR _08570_ sky130_fd_sc_hd__buf_6
X_29953_ net323 _01688_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[15\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_25076_ _10769_ VGND VGND VPWR VPWR _02596_ sky130_fd_sc_hd__clkbuf_1
X_22288_ _09423_ VGND VGND VPWR VPWR _09453_ sky130_fd_sc_hd__buf_4
X_28904_ _12747_ net4250 net68 VGND VGND VPWR VPWR _12957_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_208_5486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold280 datamem.data_ram\[30\]\[4\] VGND VGND VPWR VPWR net1430 sky130_fd_sc_hd__dlygate4sd3_1
X_21239_ datamem.data_ram\[53\]\[8\] datamem.data_ram\[52\]\[8\] datamem.data_ram\[52\]\[1\]
+ datamem.data_ram\[53\]\[1\] VGND VGND VPWR VPWR _08502_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_208_5497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold291 datamem.data_ram\[32\]\[0\] VGND VGND VPWR VPWR net1441 sky130_fd_sc_hd__dlygate4sd3_1
X_29884_ net262 _01619_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[17\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28835_ _12920_ VGND VGND VPWR VPWR _04204_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_161_4354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_161_4365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23465__114 clknet_1_1__leaf__10157_ VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__inv_2
XFILLER_0_205_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15800_ _14189_ net2537 _14221_ VGND VGND VPWR VPWR _14230_ sky130_fd_sc_hd__mux2_1
X_16780_ _04636_ VGND VGND VPWR VPWR _01654_ sky130_fd_sc_hd__clkbuf_1
X_28766_ _12883_ VGND VGND VPWR VPWR _04172_ sky130_fd_sc_hd__clkbuf_1
X_25978_ _11146_ VGND VGND VPWR VPWR _11312_ sky130_fd_sc_hd__buf_2
XFILLER_0_217_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15731_ _14191_ net4015 _14173_ VGND VGND VPWR VPWR _14192_ sky130_fd_sc_hd__mux2_1
X_23994__528 clknet_1_1__leaf__10240_ VGND VGND VPWR VPWR net654 sky130_fd_sc_hd__inv_2
X_27717_ _12157_ net3494 net50 VGND VGND VPWR VPWR _12297_ sky130_fd_sc_hd__mux2_1
X_24929_ _10474_ net3795 net91 VGND VGND VPWR VPWR _10683_ sky130_fd_sc_hd__mux2_1
XFILLER_0_217_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28697_ _12745_ net3599 net42 VGND VGND VPWR VPWR _12847_ sky130_fd_sc_hd__mux2_1
XFILLER_0_217_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18450_ _05810_ _05791_ _05812_ VGND VGND VPWR VPWR _05813_ sky130_fd_sc_hd__a21oi_1
XANTENNA_120 _07203_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27648_ _12259_ VGND VGND VPWR VPWR _03678_ sky130_fd_sc_hd__clkbuf_1
X_15662_ _13203_ VGND VGND VPWR VPWR _14145_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_64_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_131 _07821_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17401_ _14183_ net3997 _04960_ VGND VGND VPWR VPWR _04966_ sky130_fd_sc_hd__mux2_1
XANTENNA_142 _07836_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_200_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14613_ rvcpu.dp.plmw.ALUResultW\[27\] rvcpu.dp.plmw.ReadDataW\[27\] rvcpu.dp.plmw.PCPlus4W\[27\]
+ rvcpu.dp.plmw.lAuiPCW\[27\] _13192_ _13193_ VGND VGND VPWR VPWR _13194_ sky130_fd_sc_hd__mux4_2
XFILLER_0_150_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_3372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_153 _07912_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18381_ _05742_ _05744_ VGND VGND VPWR VPWR _05745_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_120_3383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15593_ _14104_ VGND VGND VPWR VPWR _02209_ sky130_fd_sc_hd__clkbuf_1
X_23009__714 clknet_1_0__leaf__10085_ VGND VGND VPWR VPWR net840 sky130_fd_sc_hd__inv_2
XANTENNA_164 _08653_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_175 _08809_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27579_ _12095_ net2635 net82 VGND VGND VPWR VPWR _12223_ sky130_fd_sc_hd__mux2_1
XFILLER_0_200_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_186 _09163_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_185_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29318_ clknet_leaf_11_clk _01053_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD1E\[25\] sky130_fd_sc_hd__dfxtp_1
X_17332_ _04929_ VGND VGND VPWR VPWR _01379_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_197 _09410_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_30590_ clknet_leaf_117_clk _02325_ VGND VGND VPWR VPWR datamem.data_ram\[53\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29249_ _09243_ net2870 _13141_ VGND VGND VPWR VPWR _13145_ sky130_fd_sc_hd__mux2_1
X_17263_ _04892_ VGND VGND VPWR VPWR _01411_ sky130_fd_sc_hd__clkbuf_1
X_24031__562 clknet_1_0__leaf__10243_ VGND VGND VPWR VPWR net688 sky130_fd_sc_hd__inv_2
XFILLER_0_187_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_183_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19002_ _05298_ _05558_ VGND VGND VPWR VPWR _06336_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16214_ _13240_ VGND VGND VPWR VPWR _14461_ sky130_fd_sc_hd__buf_4
XFILLER_0_180_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17194_ _14181_ net2755 _04851_ VGND VGND VPWR VPWR _04856_ sky130_fd_sc_hd__mux2_1
X_32260_ clknet_leaf_256_clk _03682_ VGND VGND VPWR VPWR datamem.data_ram\[34\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload106 clknet_leaf_160_clk VGND VGND VPWR VPWR clkload106/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_0_84_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_871 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload117 clknet_leaf_96_clk VGND VGND VPWR VPWR clkload117/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_148_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_168_4519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload128 clknet_leaf_256_clk VGND VGND VPWR VPWR clkload128/Y sky130_fd_sc_hd__clkinv_4
X_31211_ clknet_leaf_42_clk net1680 VGND VGND VPWR VPWR rvcpu.dp.plfd.PCD\[0\] sky130_fd_sc_hd__dfxtp_1
X_16145_ _14415_ VGND VGND VPWR VPWR _01952_ sky130_fd_sc_hd__clkbuf_1
Xclkload139 clknet_leaf_244_clk VGND VGND VPWR VPWR clkload139/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_94_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32191_ clknet_leaf_270_clk _03613_ VGND VGND VPWR VPWR datamem.data_ram\[37\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_94_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22994__700 clknet_1_1__leaf__10084_ VGND VGND VPWR VPWR net826 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_173_Left_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31142_ clknet_leaf_66_clk rvcpu.ALUResultE\[1\] VGND VGND VPWR VPWR rvcpu.dp.plem.ALUResultM\[1\]
+ sky130_fd_sc_hd__dfxtp_4
X_23317__957 clknet_1_1__leaf__10134_ VGND VGND VPWR VPWR net1083 sky130_fd_sc_hd__inv_2
X_16076_ net2027 _13266_ _14371_ VGND VGND VPWR VPWR _14379_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_90_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15027_ _13397_ _13414_ VGND VGND VPWR VPWR _13574_ sky130_fd_sc_hd__nand2_1
X_19904_ datamem.data_ram\[11\]\[17\] _06863_ _07020_ datamem.data_ram\[15\]\[17\]
+ _06602_ VGND VGND VPWR VPWR _07199_ sky130_fd_sc_hd__o221a_1
XFILLER_0_121_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31073_ clknet_leaf_164_clk _02808_ VGND VGND VPWR VPWR datamem.data_ram\[9\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2609 datamem.data_ram\[62\]\[8\] VGND VGND VPWR VPWR net3759 sky130_fd_sc_hd__dlygate4sd3_1
X_30024_ net386 _01759_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[13\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19835_ datamem.data_ram\[33\]\[1\] _06997_ _07124_ _07129_ VGND VGND VPWR VPWR _07130_
+ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_127_3537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_3548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1908 datamem.data_ram\[17\]\[9\] VGND VGND VPWR VPWR net3058 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1919 datamem.data_ram\[18\]\[21\] VGND VGND VPWR VPWR net3069 sky130_fd_sc_hd__dlygate4sd3_1
X_19766_ datamem.data_ram\[18\]\[25\] _06692_ _06779_ datamem.data_ram\[16\]\[25\]
+ VGND VGND VPWR VPWR _07061_ sky130_fd_sc_hd__o22a_1
XFILLER_0_21_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16978_ net2191 _14461_ _04731_ VGND VGND VPWR VPWR _04741_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_223_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18717_ _05410_ _05419_ _06039_ _05608_ VGND VGND VPWR VPWR _06069_ sky130_fd_sc_hd__o31ai_2
X_15929_ _14300_ VGND VGND VPWR VPWR _02061_ sky130_fd_sc_hd__clkbuf_1
X_19697_ _06925_ VGND VGND VPWR VPWR _06993_ sky130_fd_sc_hd__buf_4
XFILLER_0_189_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31975_ clknet_leaf_155_clk _03397_ VGND VGND VPWR VPWR datamem.data_ram\[53\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_88_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_182_Left_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30926_ clknet_leaf_155_clk _02661_ VGND VGND VPWR VPWR datamem.data_ram\[40\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_18648_ _05789_ VGND VGND VPWR VPWR _06004_ sky130_fd_sc_hd__buf_2
XFILLER_0_149_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23363__999 clknet_1_0__leaf__10138_ VGND VGND VPWR VPWR net1125 sky130_fd_sc_hd__inv_2
XFILLER_0_47_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_308 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18579_ _05358_ _05664_ _05802_ _05689_ VGND VGND VPWR VPWR _05938_ sky130_fd_sc_hd__o211a_1
X_30857_ clknet_leaf_152_clk _02592_ VGND VGND VPWR VPWR datamem.data_ram\[43\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20610_ datamem.data_ram\[42\]\[13\] _06804_ _07037_ datamem.data_ram\[45\]\[13\]
+ VGND VGND VPWR VPWR _07901_ sky130_fd_sc_hd__o22a_1
XFILLER_0_163_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21590_ _08673_ VGND VGND VPWR VPWR _08842_ sky130_fd_sc_hd__clkbuf_4
X_30788_ clknet_leaf_135_clk _02523_ VGND VGND VPWR VPWR datamem.data_ram\[46\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20541_ _07831_ VGND VGND VPWR VPWR _07832_ sky130_fd_sc_hd__buf_6
XFILLER_0_172_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32527_ clknet_leaf_274_clk _03949_ VGND VGND VPWR VPWR datamem.data_ram\[24\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20472_ datamem.data_ram\[38\]\[20\] _06628_ _07230_ datamem.data_ram\[36\]\[20\]
+ VGND VGND VPWR VPWR _07764_ sky130_fd_sc_hd__o22a_1
XFILLER_0_6_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32458_ clknet_leaf_239_clk _03880_ VGND VGND VPWR VPWR datamem.data_ram\[26\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_191_Left_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22211_ _09378_ VGND VGND VPWR VPWR _01122_ sky130_fd_sc_hd__clkbuf_1
X_31409_ clknet_leaf_27_clk _03112_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCE\[26\] sky130_fd_sc_hd__dfxtp_1
X_23191_ _10116_ VGND VGND VPWR VPWR _01364_ sky130_fd_sc_hd__clkbuf_1
X_32389_ clknet_leaf_232_clk _03811_ VGND VGND VPWR VPWR datamem.data_ram\[29\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22142_ _09340_ VGND VGND VPWR VPWR _01091_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_219_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26950_ _11827_ _11854_ VGND VGND VPWR VPWR _11857_ sky130_fd_sc_hd__and2_1
X_22073_ _09288_ net2180 _09270_ VGND VGND VPWR VPWR _09289_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25901_ _13368_ _11268_ VGND VGND VPWR VPWR _11269_ sky130_fd_sc_hd__nand2_1
X_21024_ datamem.data_ram\[30\]\[31\] datamem.data_ram\[31\]\[31\] _07912_ VGND VGND
+ VPWR VPWR _08313_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26881_ _11795_ net1412 _11809_ _11812_ VGND VGND VPWR VPWR _03358_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_203_5361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28620_ _12806_ VGND VGND VPWR VPWR _04103_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_203_5372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25832_ _11217_ VGND VGND VPWR VPWR _02904_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28551_ _12769_ VGND VGND VPWR VPWR _04071_ sky130_fd_sc_hd__clkbuf_1
X_25763_ _11149_ _11163_ VGND VGND VPWR VPWR _11164_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_195_5173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27502_ _12182_ VGND VGND VPWR VPWR _03609_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_195_5184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24714_ _10472_ net4012 net59 VGND VGND VPWR VPWR _10565_ sky130_fd_sc_hd__mux2_1
X_21926_ _08623_ _09151_ _09155_ _09159_ VGND VGND VPWR VPWR _09160_ sky130_fd_sc_hd__and4_1
XFILLER_0_96_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25694_ _11089_ _11113_ VGND VGND VPWR VPWR _11119_ sky130_fd_sc_hd__and2_1
X_28482_ _11965_ _12724_ VGND VGND VPWR VPWR _12725_ sky130_fd_sc_hd__and2_1
XFILLER_0_139_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27433_ _12140_ net2130 _12126_ VGND VGND VPWR VPWR _12141_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24645_ _10526_ VGND VGND VPWR VPWR _02408_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21857_ _09092_ _09093_ _08743_ VGND VGND VPWR VPWR _09094_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20808_ datamem.data_ram\[46\]\[30\] datamem.data_ram\[47\]\[30\] _07826_ VGND VGND
+ VPWR VPWR _08098_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24576_ _10488_ VGND VGND VPWR VPWR _02377_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27364_ _12100_ VGND VGND VPWR VPWR _03553_ sky130_fd_sc_hd__clkbuf_1
X_21788_ _08795_ _09024_ _09026_ _09028_ VGND VGND VPWR VPWR _09029_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_148_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29103_ _13066_ VGND VGND VPWR VPWR _04326_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26315_ _11490_ VGND VGND VPWR VPWR _03114_ sky130_fd_sc_hd__clkbuf_1
X_23527_ clknet_1_1__leaf__10152_ VGND VGND VPWR VPWR _10171_ sky130_fd_sc_hd__buf_1
XFILLER_0_37_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27295_ _12036_ net1611 _12053_ _12060_ VGND VGND VPWR VPWR _03524_ sky130_fd_sc_hd__a31o_1
X_20739_ datamem.data_ram\[33\]\[6\] _06997_ _08024_ _07636_ _08028_ VGND VGND VPWR
+ VPWR _08029_ sky130_fd_sc_hd__a221o_1
XFILLER_0_167_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_4180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_4191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29034_ _10932_ _10778_ VGND VGND VPWR VPWR _13029_ sky130_fd_sc_hd__or2_1
X_26246_ _11438_ _11458_ _11459_ _09482_ VGND VGND VPWR VPWR _03076_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_162_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23575__197 clknet_1_0__leaf__10176_ VGND VGND VPWR VPWR net323 sky130_fd_sc_hd__inv_2
XFILLER_0_34_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_150_4088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_4099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22409_ _09461_ _09567_ _09569_ _09474_ VGND VGND VPWR VPWR _09570_ sky130_fd_sc_hd__o211a_1
XFILLER_0_162_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26177_ _11425_ VGND VGND VPWR VPWR _03041_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_180_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23389_ _10145_ VGND VGND VPWR VPWR _01533_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25128_ _10470_ net3942 net87 VGND VGND VPWR VPWR _10796_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_163_4405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_163_4416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25059_ _09243_ VGND VGND VPWR VPWR _10758_ sky130_fd_sc_hd__buf_2
X_17950_ _05321_ rvcpu.dp.plde.ImmExtE\[13\] VGND VGND VPWR VPWR _05322_ sky130_fd_sc_hd__nand2_1
X_29936_ net306 _01671_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[16\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16901_ _04700_ VGND VGND VPWR VPWR _01589_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_178_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24061__588 clknet_1_0__leaf__10247_ VGND VGND VPWR VPWR net714 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_168_Right_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17881_ rvcpu.dp.plde.Rs1E\[0\] rvcpu.dp.plmw.RegWriteW VGND VGND VPWR VPWR _05254_
+ sky130_fd_sc_hd__or2b_1
X_29867_ net245 _01602_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[18\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_228_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19620_ _06753_ VGND VGND VPWR VPWR _06916_ sky130_fd_sc_hd__buf_4
X_16832_ net2750 _14451_ _04659_ VGND VGND VPWR VPWR _04664_ sky130_fd_sc_hd__mux2_1
X_28818_ _12911_ VGND VGND VPWR VPWR _04196_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_217_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29798_ clknet_leaf_208_clk _01533_ VGND VGND VPWR VPWR datamem.data_ram\[59\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_205_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_3412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19551_ datamem.data_ram\[17\]\[24\] _06658_ _06843_ _06846_ VGND VGND VPWR VPWR
+ _06847_ sky130_fd_sc_hd__o211a_1
XFILLER_0_221_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_122_3423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16763_ _04627_ VGND VGND VPWR VPWR _01662_ sky130_fd_sc_hd__clkbuf_1
X_28749_ _12874_ VGND VGND VPWR VPWR _04164_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_122_3434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18502_ _05862_ _05863_ VGND VGND VPWR VPWR _05864_ sky130_fd_sc_hd__or2_2
XFILLER_0_214_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15714_ _14180_ VGND VGND VPWR VPWR _02164_ sky130_fd_sc_hd__clkbuf_1
X_31760_ clknet_leaf_105_clk _03214_ VGND VGND VPWR VPWR datamem.data_ram\[18\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_19482_ _06646_ VGND VGND VPWR VPWR _06778_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_186_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16694_ _14158_ net4249 _04587_ VGND VGND VPWR VPWR _04591_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18433_ _05689_ _05685_ VGND VGND VPWR VPWR _05796_ sky130_fd_sc_hd__nand2_1
X_30711_ clknet_leaf_192_clk _02446_ VGND VGND VPWR VPWR datamem.data_ram\[49\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_15645_ _14133_ net4161 _14131_ VGND VGND VPWR VPWR _14134_ sky130_fd_sc_hd__mux2_1
X_31691_ clknet_leaf_33_clk _03149_ VGND VGND VPWR VPWR rvcpu.dp.pcreg.q\[9\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_180_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30642_ clknet_leaf_139_clk _02377_ VGND VGND VPWR VPWR datamem.data_ram\[51\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_18364_ _05236_ _05659_ VGND VGND VPWR VPWR _05729_ sky130_fd_sc_hd__nor2_2
XFILLER_0_12_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15576_ _14095_ VGND VGND VPWR VPWR _02217_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17315_ _04920_ VGND VGND VPWR VPWR _01387_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_185_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18295_ rvcpu.dp.plde.ALUControlE\[2\] _05659_ rvcpu.dp.plde.ALUControlE\[3\] VGND
+ VGND VPWR VPWR _05660_ sky130_fd_sc_hd__or3b_4
XTAP_TAPCELL_ROW_96_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30573_ clknet_leaf_181_clk _02308_ VGND VGND VPWR VPWR datamem.data_ram\[54\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23061__760 clknet_1_0__leaf__10091_ VGND VGND VPWR VPWR net886 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_21_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32312_ clknet_leaf_276_clk _03734_ VGND VGND VPWR VPWR datamem.data_ram\[32\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17246_ _04883_ VGND VGND VPWR VPWR _01419_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32243_ clknet_leaf_211_clk _03665_ VGND VGND VPWR VPWR datamem.data_ram\[34\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17177_ _14164_ net4341 _04840_ VGND VGND VPWR VPWR _04847_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16128_ _14406_ VGND VGND VPWR VPWR _01960_ sky130_fd_sc_hd__clkbuf_1
X_32174_ clknet_leaf_215_clk _03596_ VGND VGND VPWR VPWR datamem.data_ram\[37\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31125_ clknet_leaf_125_clk _02860_ VGND VGND VPWR VPWR datamem.data_ram\[25\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3107 rvcpu.dp.rf.reg_file_arr\[8\]\[14\] VGND VGND VPWR VPWR net4257 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3118 rvcpu.dp.rf.reg_file_arr\[24\]\[10\] VGND VGND VPWR VPWR net4268 sky130_fd_sc_hd__dlygate4sd3_1
X_16059_ net1881 _13241_ _14360_ VGND VGND VPWR VPWR _14370_ sky130_fd_sc_hd__mux2_1
Xhold3129 datamem.data_ram\[57\]\[18\] VGND VGND VPWR VPWR net4279 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2406 datamem.data_ram\[13\]\[13\] VGND VGND VPWR VPWR net3556 sky130_fd_sc_hd__dlygate4sd3_1
X_31056_ clknet_leaf_115_clk _02791_ VGND VGND VPWR VPWR datamem.data_ram\[38\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2417 datamem.data_ram\[14\]\[19\] VGND VGND VPWR VPWR net3567 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_135_Right_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2428 datamem.data_ram\[55\]\[14\] VGND VGND VPWR VPWR net3578 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2439 datamem.data_ram\[29\]\[19\] VGND VGND VPWR VPWR net3589 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1705 rvcpu.dp.rf.reg_file_arr\[7\]\[6\] VGND VGND VPWR VPWR net2855 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1716 rvcpu.dp.rf.reg_file_arr\[15\]\[29\] VGND VGND VPWR VPWR net2866 sky130_fd_sc_hd__dlygate4sd3_1
X_19818_ datamem.data_ram\[24\]\[9\] _06647_ _06782_ datamem.data_ram\[25\]\[9\] VGND
+ VGND VPWR VPWR _07113_ sky130_fd_sc_hd__o22a_1
X_30007_ clknet_leaf_265_clk _01742_ VGND VGND VPWR VPWR datamem.data_ram\[59\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1727 datamem.data_ram\[13\]\[19\] VGND VGND VPWR VPWR net2877 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1738 datamem.data_ram\[58\]\[13\] VGND VGND VPWR VPWR net2888 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1749 datamem.data_ram\[28\]\[29\] VGND VGND VPWR VPWR net2899 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19749_ datamem.data_ram\[45\]\[25\] _06723_ _06807_ datamem.data_ram\[40\]\[25\]
+ _07043_ VGND VGND VPWR VPWR _07044_ sky130_fd_sc_hd__o221a_1
XFILLER_0_154_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22760_ rvcpu.dp.rf.reg_file_arr\[24\]\[24\] rvcpu.dp.rf.reg_file_arr\[25\]\[24\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[24\] rvcpu.dp.rf.reg_file_arr\[27\]\[24\] _09406_
+ _09395_ VGND VGND VPWR VPWR _09902_ sky130_fd_sc_hd__mux4_2
X_31958_ clknet_leaf_133_clk _03380_ VGND VGND VPWR VPWR datamem.data_ram\[55\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_480 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21711_ _08725_ _08955_ VGND VGND VPWR VPWR _08956_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_49_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30909_ clknet_leaf_263_clk _02644_ VGND VGND VPWR VPWR datamem.data_ram\[41\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_49_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22691_ rvcpu.dp.rf.reg_file_arr\[24\]\[20\] rvcpu.dp.rf.reg_file_arr\[25\]\[20\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[20\] rvcpu.dp.rf.reg_file_arr\[27\]\[20\] _09392_
+ _09394_ VGND VGND VPWR VPWR _09837_ sky130_fd_sc_hd__mux4_1
X_31889_ clknet_leaf_113_clk _03343_ VGND VGND VPWR VPWR datamem.data_ram\[36\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24430_ _09287_ VGND VGND VPWR VPWR _10398_ sky130_fd_sc_hd__buf_2
X_21642_ rvcpu.dp.rf.reg_file_arr\[0\]\[13\] rvcpu.dp.rf.reg_file_arr\[1\]\[13\] rvcpu.dp.rf.reg_file_arr\[2\]\[13\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[13\] _08810_ _08811_ VGND VGND VPWR VPWR _08891_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_192_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24361_ _10358_ VGND VGND VPWR VPWR _02292_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_192_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_191_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_20 _06615_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21573_ _08552_ VGND VGND VPWR VPWR _08825_ sky130_fd_sc_hd__buf_4
X_23494__140 clknet_1_0__leaf__10160_ VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__inv_2
XFILLER_0_7_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_31 _06645_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26100_ net1571 _11372_ VGND VGND VPWR VPWR _11385_ sky130_fd_sc_hd__and2_1
XANTENNA_42 _06678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27080_ _11153_ _11146_ VGND VGND VPWR VPWR _11933_ sky130_fd_sc_hd__nor2_1
X_20524_ datamem.data_ram\[23\]\[21\] _07021_ _06659_ datamem.data_ram\[17\]\[21\]
+ VGND VGND VPWR VPWR _07815_ sky130_fd_sc_hd__o22a_1
XFILLER_0_144_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_53 _06702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_64 _06752_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24292_ _10319_ VGND VGND VPWR VPWR _02262_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_75 _06776_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26031_ _11121_ net1746 _11339_ _11342_ VGND VGND VPWR VPWR _02978_ sky130_fd_sc_hd__a31o_1
XFILLER_0_160_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_86 _06784_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_97 _06815_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20455_ _06680_ _07739_ _07741_ _07746_ VGND VGND VPWR VPWR _07747_ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20386_ datamem.data_ram\[50\]\[28\] _06803_ _07674_ _07677_ VGND VGND VPWR VPWR
+ _07678_ sky130_fd_sc_hd__o211a_1
XFILLER_0_179_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_219_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22125_ _09331_ VGND VGND VPWR VPWR _01083_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_282_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_282_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_205_5412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_1298 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_205_5423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27982_ _12447_ net3922 net76 VGND VGND VPWR VPWR _12449_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29721_ net1067 _01456_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[22\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_26933_ _11831_ net1489 _11841_ _11846_ VGND VGND VPWR VPWR _03376_ sky130_fd_sc_hd__a31o_1
X_22056_ _09275_ VGND VGND VPWR VPWR _09276_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_201_5309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_102_Right_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_197_5213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2940 rvcpu.dp.rf.reg_file_arr\[20\]\[11\] VGND VGND VPWR VPWR net4090 sky130_fd_sc_hd__dlygate4sd3_1
X_21007_ _08287_ _08289_ _08291_ _08295_ VGND VGND VPWR VPWR _08296_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_197_5224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29652_ net998 _01387_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[24\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_26864_ _11684_ _11798_ VGND VGND VPWR VPWR _11802_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_197_5235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2951 datamem.data_ram\[9\]\[22\] VGND VGND VPWR VPWR net4101 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2962 datamem.data_ram\[59\]\[13\] VGND VGND VPWR VPWR net4112 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2973 datamem.data_ram\[15\]\[18\] VGND VGND VPWR VPWR net4123 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2984 datamem.data_ram\[4\]\[18\] VGND VGND VPWR VPWR net4134 sky130_fd_sc_hd__dlygate4sd3_1
X_28603_ _12797_ VGND VGND VPWR VPWR _04095_ sky130_fd_sc_hd__clkbuf_1
X_25815_ rvcpu.dp.pcreg.q\[20\] _11200_ VGND VGND VPWR VPWR _11203_ sky130_fd_sc_hd__nand2_1
Xhold2995 rvcpu.dp.rf.reg_file_arr\[5\]\[30\] VGND VGND VPWR VPWR net4145 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29583_ net937 _01318_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[26\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_26795_ _07191_ _11725_ _11494_ VGND VGND VPWR VPWR _11760_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_3_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28534_ _09243_ VGND VGND VPWR VPWR _12758_ sky130_fd_sc_hd__buf_2
X_25746_ net1660 _11144_ _11147_ _11150_ VGND VGND VPWR VPWR _02885_ sky130_fd_sc_hd__o211a_1
Xmax_cap44 _12592_ VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__buf_4
Xmax_cap55 _10857_ VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__buf_4
XFILLER_0_97_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_186_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap66 _13020_ VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__buf_4
X_21909_ _09143_ VGND VGND VPWR VPWR _01055_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap77 _12382_ VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__buf_4
Xmax_cap88 _10784_ VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__buf_4
X_28465_ _12450_ net3562 _12713_ VGND VGND VPWR VPWR _12715_ sky130_fd_sc_hd__mux2_1
X_25677_ _11064_ _11098_ VGND VGND VPWR VPWR _11108_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_156_4231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22889_ _09380_ _10023_ VGND VGND VPWR VPWR _10024_ sky130_fd_sc_hd__or2_1
Xmax_cap99 _12188_ VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_156_4242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15430_ _13958_ _13960_ VGND VGND VPWR VPWR _13961_ sky130_fd_sc_hd__nor2_1
X_27416_ _12129_ VGND VGND VPWR VPWR _03576_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_214_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24628_ _10450_ net3317 _10511_ VGND VGND VPWR VPWR _10517_ sky130_fd_sc_hd__mux2_1
X_28396_ _12674_ VGND VGND VPWR VPWR _04011_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_14_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15361_ _13370_ _13862_ _13858_ _13442_ VGND VGND VPWR VPWR _13896_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_152_4139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27347_ _12089_ net4215 _12081_ VGND VGND VPWR VPWR _12090_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24559_ _10478_ net2691 net60 VGND VGND VPWR VPWR _10479_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17100_ _04806_ VGND VGND VPWR VPWR _01488_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15292_ _13643_ _13829_ _13581_ VGND VGND VPWR VPWR _13830_ sky130_fd_sc_hd__a21oi_1
X_18080_ _05416_ VGND VGND VPWR VPWR _05448_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27278_ _12050_ VGND VGND VPWR VPWR _03517_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17031_ net2475 _14445_ _04768_ VGND VGND VPWR VPWR _04770_ sky130_fd_sc_hd__mux2_1
X_29017_ _10141_ _11020_ _12977_ VGND VGND VPWR VPWR _13020_ sky130_fd_sc_hd__a21oi_2
X_26229_ _11453_ VGND VGND VPWR VPWR _11454_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_115_3260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_468 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_5_31__f_clk clknet_2_3_0_clk VGND VGND VPWR VPWR clknet_5_31__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_22_945 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_186_4950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_186_4961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_3168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_273_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_273_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_104_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18982_ _06314_ _06315_ _06316_ _06317_ VGND VGND VPWR VPWR _06318_ sky130_fd_sc_hd__or4b_1
XFILLER_0_21_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_182_4858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_182_4869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17933_ rvcpu.dp.plde.RD1E\[14\] _05293_ _05263_ VGND VGND VPWR VPWR _05306_ sky130_fd_sc_hd__and3_1
X_29919_ net289 _01654_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[16\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32930_ clknet_leaf_156_clk _04352_ VGND VGND VPWR VPWR datamem.data_ram\[7\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_17864_ _05237_ VGND VGND VPWR VPWR _00003_ sky130_fd_sc_hd__buf_2
XFILLER_0_205_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_178_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19603_ datamem.data_ram\[18\]\[8\] _06804_ _06806_ datamem.data_ram\[20\]\[8\] _06898_
+ VGND VGND VPWR VPWR _06899_ sky130_fd_sc_hd__o221a_1
XFILLER_0_17_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16815_ net1865 _14434_ _04648_ VGND VGND VPWR VPWR _04655_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32861_ clknet_leaf_55_clk _04283_ VGND VGND VPWR VPWR datamem.data_ram\[11\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17795_ rvcpu.dp.plem.ALUResultM\[3\] _05175_ _05188_ _05189_ VGND VGND VPWR VPWR
+ _05190_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_85_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_85_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31812_ clknet_leaf_109_clk _03266_ VGND VGND VPWR VPWR datamem.data_ram\[17\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19534_ datamem.data_ram\[38\]\[24\] _06718_ _06686_ datamem.data_ram\[36\]\[24\]
+ VGND VGND VPWR VPWR _06830_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_141_3876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16746_ _04618_ VGND VGND VPWR VPWR _01670_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_141_3887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32792_ clknet_leaf_283_clk _04214_ VGND VGND VPWR VPWR datamem.data_ram\[14\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19465_ _06760_ VGND VGND VPWR VPWR _06761_ sky130_fd_sc_hd__clkbuf_8
X_31743_ net128 _03201_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[9\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16677_ _14141_ net3707 _04576_ VGND VGND VPWR VPWR _04582_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18416_ _05778_ _05779_ _05677_ VGND VGND VPWR VPWR _05780_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15628_ _14122_ VGND VGND VPWR VPWR _02192_ sky130_fd_sc_hd__clkbuf_1
X_31674_ clknet_leaf_29_clk net1279 VGND VGND VPWR VPWR rvcpu.dp.plmw.ALUResultW\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19396_ _06691_ VGND VGND VPWR VPWR _06692_ sky130_fd_sc_hd__buf_8
XFILLER_0_57_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24111__618 clknet_1_0__leaf__10259_ VGND VGND VPWR VPWR net744 sky130_fd_sc_hd__inv_2
XFILLER_0_1_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18347_ _05671_ _05708_ _05710_ _05286_ _05711_ VGND VGND VPWR VPWR _05712_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_44_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30625_ clknet_leaf_178_clk _02360_ VGND VGND VPWR VPWR datamem.data_ram\[52\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_15559_ _13301_ _13767_ _13481_ _13797_ _14082_ VGND VGND VPWR VPWR _14083_ sky130_fd_sc_hd__o32a_1
XFILLER_0_5_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_100_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18278_ _05300_ VGND VGND VPWR VPWR _05643_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30556_ clknet_leaf_177_clk _02291_ VGND VGND VPWR VPWR datamem.data_ram\[55\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_204_Right_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_226_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17229_ _04874_ VGND VGND VPWR VPWR _01427_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30487_ clknet_leaf_198_clk _02222_ VGND VGND VPWR VPWR datamem.data_ram\[57\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold802 datamem.data_ram\[44\]\[23\] VGND VGND VPWR VPWR net1952 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20240_ datamem.data_ram\[55\]\[3\] _06927_ _07532_ _06967_ VGND VGND VPWR VPWR _07533_
+ sky130_fd_sc_hd__a211o_1
X_32226_ clknet_leaf_87_clk _03648_ VGND VGND VPWR VPWR datamem.data_ram\[35\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold813 rvcpu.dp.rf.reg_file_arr\[7\]\[9\] VGND VGND VPWR VPWR net1963 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold824 rvcpu.dp.rf.reg_file_arr\[6\]\[19\] VGND VGND VPWR VPWR net1974 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold835 rvcpu.dp.rf.reg_file_arr\[10\]\[20\] VGND VGND VPWR VPWR net1985 sky130_fd_sc_hd__dlygate4sd3_1
Xhold846 datamem.data_ram\[4\]\[31\] VGND VGND VPWR VPWR net1996 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_264_clk clknet_5_17__leaf_clk VGND VGND VPWR VPWR clknet_leaf_264_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold857 rvcpu.dp.rf.reg_file_arr\[5\]\[11\] VGND VGND VPWR VPWR net2007 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32157_ clknet_leaf_167_clk _03579_ VGND VGND VPWR VPWR datamem.data_ram\[38\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_20171_ datamem.data_ram\[30\]\[11\] _06764_ _06761_ datamem.data_ram\[31\]\[11\]
+ VGND VGND VPWR VPWR _07464_ sky130_fd_sc_hd__o22a_1
Xhold868 rvcpu.dp.rf.reg_file_arr\[10\]\[0\] VGND VGND VPWR VPWR net2018 sky130_fd_sc_hd__dlygate4sd3_1
Xhold879 datamem.data_ram\[2\]\[31\] VGND VGND VPWR VPWR net2029 sky130_fd_sc_hd__dlygate4sd3_1
X_31108_ clknet_leaf_106_clk _02843_ VGND VGND VPWR VPWR datamem.data_ram\[19\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2203 datamem.data_ram\[16\]\[9\] VGND VGND VPWR VPWR net3353 sky130_fd_sc_hd__dlygate4sd3_1
X_32088_ clknet_leaf_73_clk _03510_ VGND VGND VPWR VPWR datamem.data_ram\[47\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2214 datamem.data_ram\[28\]\[17\] VGND VGND VPWR VPWR net3364 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2225 datamem.data_ram\[8\]\[8\] VGND VGND VPWR VPWR net3375 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2236 datamem.data_ram\[43\]\[26\] VGND VGND VPWR VPWR net3386 sky130_fd_sc_hd__dlygate4sd3_1
X_31039_ clknet_leaf_97_clk _02774_ VGND VGND VPWR VPWR datamem.data_ram\[41\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1502 rvcpu.dp.rf.reg_file_arr\[21\]\[7\] VGND VGND VPWR VPWR net2652 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2247 datamem.data_ram\[9\]\[28\] VGND VGND VPWR VPWR net3397 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1513 datamem.data_ram\[17\]\[19\] VGND VGND VPWR VPWR net2663 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2258 rvcpu.dp.rf.reg_file_arr\[19\]\[25\] VGND VGND VPWR VPWR net3408 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1524 rvcpu.dp.rf.reg_file_arr\[5\]\[2\] VGND VGND VPWR VPWR net2674 sky130_fd_sc_hd__dlygate4sd3_1
X_22972__680 clknet_1_0__leaf__10082_ VGND VGND VPWR VPWR net806 sky130_fd_sc_hd__inv_2
Xhold2269 datamem.data_ram\[48\]\[10\] VGND VGND VPWR VPWR net3419 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1535 rvcpu.dp.rf.reg_file_arr\[12\]\[11\] VGND VGND VPWR VPWR net2685 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_165_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1546 rvcpu.dp.rf.reg_file_arr\[16\]\[17\] VGND VGND VPWR VPWR net2696 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1557 rvcpu.dp.rf.reg_file_arr\[18\]\[6\] VGND VGND VPWR VPWR net2707 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1568 rvcpu.dp.rf.reg_file_arr\[28\]\[13\] VGND VGND VPWR VPWR net2718 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1579 rvcpu.dp.rf.reg_file_arr\[15\]\[25\] VGND VGND VPWR VPWR net2729 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25600_ _11057_ net1501 _11053_ _11063_ VGND VGND VPWR VPWR _02826_ sky130_fd_sc_hd__a31o_1
X_22812_ _09461_ _09949_ _09951_ _09489_ VGND VGND VPWR VPWR _09952_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_192_5110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26580_ _11635_ VGND VGND VPWR VPWR _03234_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_211_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0__10180_ _10180_ VGND VGND VPWR VPWR clknet_0__10180_ sky130_fd_sc_hd__clkbuf_16
X_22743_ rvcpu.dp.rf.reg_file_arr\[20\]\[23\] rvcpu.dp.rf.reg_file_arr\[21\]\[23\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[23\] rvcpu.dp.rf.reg_file_arr\[23\]\[23\] _09517_
+ _09577_ VGND VGND VPWR VPWR _09886_ sky130_fd_sc_hd__mux4_2
XFILLER_0_67_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25531_ _11023_ VGND VGND VPWR VPWR _02797_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__10080_ clknet_0__10080_ VGND VGND VPWR VPWR clknet_1_1__leaf__10080_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_177_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_211_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25462_ _10408_ _10985_ VGND VGND VPWR VPWR _10987_ sky130_fd_sc_hd__and2_1
XFILLER_0_137_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28250_ _12452_ net4243 net44 VGND VGND VPWR VPWR _12595_ sky130_fd_sc_hd__mux2_1
XFILLER_0_220_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22674_ _09399_ _09820_ _09523_ VGND VGND VPWR VPWR _09821_ sky130_fd_sc_hd__o21a_1
XFILLER_0_191_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27201_ _12005_ net1432 _12007_ _12010_ VGND VGND VPWR VPWR _03480_ sky130_fd_sc_hd__a31o_1
XFILLER_0_30_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24413_ _10385_ datamem.data_ram\[53\]\[8\] _10386_ VGND VGND VPWR VPWR _10387_ sky130_fd_sc_hd__mux2_1
XFILLER_0_191_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21625_ _08541_ _08874_ VGND VGND VPWR VPWR _08875_ sky130_fd_sc_hd__and2_1
X_25393_ _10405_ _10950_ VGND VGND VPWR VPWR _10951_ sky130_fd_sc_hd__and2_1
X_28181_ _12435_ net4375 _12555_ VGND VGND VPWR VPWR _12558_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_1246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27132_ _11965_ _11966_ VGND VGND VPWR VPWR _11967_ sky130_fd_sc_hd__and2_1
XFILLER_0_152_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24344_ _10349_ VGND VGND VPWR VPWR _02284_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_192_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21556_ _08795_ _08797_ _08802_ _08807_ _08808_ VGND VGND VPWR VPWR _08809_ sky130_fd_sc_hd__a311o_1
XFILLER_0_173_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_209_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27063_ _10142_ _11112_ _11898_ VGND VGND VPWR VPWR _11924_ sky130_fd_sc_hd__and3_1
X_20507_ datamem.data_ram\[48\]\[21\] _07191_ _07182_ datamem.data_ram\[52\]\[21\]
+ _07797_ VGND VGND VPWR VPWR _07798_ sky130_fd_sc_hd__o221a_1
X_24275_ _10310_ VGND VGND VPWR VPWR _02254_ sky130_fd_sc_hd__clkbuf_1
X_23730__322 clknet_1_1__leaf__10198_ VGND VGND VPWR VPWR net448 sky130_fd_sc_hd__inv_2
X_21487_ _08742_ VGND VGND VPWR VPWR _08743_ sky130_fd_sc_hd__buf_4
XFILLER_0_200_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26014_ net1315 _11329_ _11325_ _11332_ VGND VGND VPWR VPWR _02971_ sky130_fd_sc_hd__o211a_1
XFILLER_0_209_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20438_ datamem.data_ram\[26\]\[12\] _06610_ _06821_ datamem.data_ram\[24\]\[12\]
+ VGND VGND VPWR VPWR _07730_ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_255_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_255_clk
+ sky130_fd_sc_hd__clkbuf_8
X_20369_ datamem.data_ram\[37\]\[28\] _06722_ _07659_ _07660_ VGND VGND VPWR VPWR
+ _07661_ sky130_fd_sc_hd__o211a_1
XFILLER_0_30_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22108_ _09317_ VGND VGND VPWR VPWR _09318_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_224_5865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_224_5876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27965_ _09243_ VGND VGND VPWR VPWR _12437_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_8_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29704_ net1050 _01439_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[22\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_14930_ _13322_ _13478_ VGND VGND VPWR VPWR _13479_ sky130_fd_sc_hd__or2_1
X_26916_ _10072_ VGND VGND VPWR VPWR _11835_ sky130_fd_sc_hd__buf_2
X_22039_ _09261_ VGND VGND VPWR VPWR _01067_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_175_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27896_ _10066_ _12394_ VGND VGND VPWR VPWR _12399_ sky130_fd_sc_hd__and2_1
XFILLER_0_227_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29635_ clknet_leaf_139_clk _01370_ VGND VGND VPWR VPWR datamem.data_ram\[5\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2770 datamem.data_ram\[63\]\[28\] VGND VGND VPWR VPWR net3920 sky130_fd_sc_hd__dlygate4sd3_1
X_26847_ _11781_ net1483 _11785_ _11791_ VGND VGND VPWR VPWR _03345_ sky130_fd_sc_hd__a31o_1
X_14861_ _13412_ _13385_ VGND VGND VPWR VPWR _13413_ sky130_fd_sc_hd__nor2_2
Xhold2781 datamem.data_ram\[32\]\[30\] VGND VGND VPWR VPWR net3931 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2792 datamem.data_ram\[42\]\[26\] VGND VGND VPWR VPWR net3942 sky130_fd_sc_hd__dlygate4sd3_1
X_16600_ _04541_ VGND VGND VPWR VPWR _01739_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_215_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29566_ net920 _01301_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[26\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_17580_ _13223_ net2662 _05057_ VGND VGND VPWR VPWR _05061_ sky130_fd_sc_hd__mux2_1
X_26778_ _11735_ net1633 _11748_ _11750_ VGND VGND VPWR VPWR _03317_ sky130_fd_sc_hd__a31o_1
X_14792_ _13280_ _13286_ VGND VGND VPWR VPWR _13345_ sky130_fd_sc_hd__or2b_1
XFILLER_0_216_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16531_ _04504_ VGND VGND VPWR VPWR _01779_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28517_ _12746_ VGND VGND VPWR VPWR _04060_ sky130_fd_sc_hd__clkbuf_1
X_25729_ _11138_ VGND VGND VPWR VPWR _02880_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_80_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29497_ net859 _01232_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[28\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19250_ rvcpu.dp.plde.ImmExtE\[30\] rvcpu.dp.plde.PCE\[30\] VGND VGND VPWR VPWR _06553_
+ sky130_fd_sc_hd__and2_1
X_28448_ _12433_ net3495 _12704_ VGND VGND VPWR VPWR _12706_ sky130_fd_sc_hd__mux2_1
X_16462_ net2170 _14420_ _04467_ VGND VGND VPWR VPWR _04468_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_175_4684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23891__451 clknet_1_0__leaf__10222_ VGND VGND VPWR VPWR net577 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_175_4695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_1302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18201_ _05506_ VGND VGND VPWR VPWR _05566_ sky130_fd_sc_hd__inv_2
XFILLER_0_156_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15413_ _13392_ _13348_ _13796_ _13513_ VGND VGND VPWR VPWR _13945_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_117_3300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19181_ _06492_ rvcpu.dp.plde.ImmExtE\[20\] _06493_ VGND VGND VPWR VPWR _06494_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_117_3311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_182_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28379_ _12367_ net3887 _12659_ VGND VGND VPWR VPWR _12665_ sky130_fd_sc_hd__mux2_1
X_16393_ _14562_ VGND VGND VPWR VPWR _01843_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_183_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18132_ _05488_ _05497_ VGND VGND VPWR VPWR _05498_ sky130_fd_sc_hd__and2_1
X_30410_ net748 _02145_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[31\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_15344_ _13387_ _13750_ VGND VGND VPWR VPWR _13880_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31390_ clknet_leaf_40_clk _03093_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCE\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_113_3208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_207_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18063_ net102 _05430_ VGND VGND VPWR VPWR _05431_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_41_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30341_ net687 _02076_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[4\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_15275_ _13385_ _13812_ _13813_ _13783_ VGND VGND VPWR VPWR _13814_ sky130_fd_sc_hd__a31o_1
XFILLER_0_124_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_184_4909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold109 rvcpu.dp.plde.RdE\[4\] VGND VGND VPWR VPWR net1259 sky130_fd_sc_hd__dlygate4sd3_1
X_17014_ net2523 _14428_ _04757_ VGND VGND VPWR VPWR _04761_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30272_ net626 _02007_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[6\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_24067__594 clknet_1_1__leaf__10247_ VGND VGND VPWR VPWR net720 sky130_fd_sc_hd__inv_2
XFILLER_0_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32011_ clknet_leaf_128_clk _03433_ VGND VGND VPWR VPWR datamem.data_ram\[27\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_246_clk clknet_5_17__leaf_clk VGND VGND VPWR VPWR clknet_leaf_246_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_111_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18965_ _05775_ _05906_ _06285_ _05275_ VGND VGND VPWR VPWR _06302_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17916_ _05286_ _05287_ VGND VGND VPWR VPWR _05289_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_37_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18896_ _05240_ _06226_ _06229_ _06237_ VGND VGND VPWR VPWR rvcpu.ALUResultE\[22\]
+ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_143_3927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32913_ clknet_leaf_156_clk _04335_ VGND VGND VPWR VPWR datamem.data_ram\[0\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_33_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17847_ rvcpu.dp.plde.RD2E\[13\] _05195_ _05225_ VGND VGND VPWR VPWR _05226_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_179_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32844_ clknet_leaf_96_clk _04266_ VGND VGND VPWR VPWR datamem.data_ram\[7\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_17778_ _05175_ VGND VGND VPWR VPWR _05176_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19517_ datamem.data_ram\[56\]\[24\] _06811_ _06812_ datamem.data_ram\[59\]\[24\]
+ VGND VGND VPWR VPWR _06813_ sky130_fd_sc_hd__o22a_1
XFILLER_0_159_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16729_ _14193_ net3899 _04575_ VGND VGND VPWR VPWR _04609_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_46_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32775_ clknet_leaf_212_clk _04197_ VGND VGND VPWR VPWR datamem.data_ram\[14\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_792 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31726_ net175 _03184_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[9\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19448_ _06743_ VGND VGND VPWR VPWR _06744_ sky130_fd_sc_hd__buf_6
XFILLER_0_186_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23141__816 clknet_1_0__leaf__10107_ VGND VGND VPWR VPWR net942 sky130_fd_sc_hd__inv_2
XFILLER_0_29_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31657_ clknet_leaf_63_clk net1626 VGND VGND VPWR VPWR rvcpu.dp.plmw.ALUResultW\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_19379_ _06585_ rvcpu.dp.plem.ALUResultM\[5\] VGND VGND VPWR VPWR _06675_ sky130_fd_sc_hd__nand2_1
XFILLER_0_174_666 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21410_ _08572_ _08669_ VGND VGND VPWR VPWR _08670_ sky130_fd_sc_hd__or2_1
X_30608_ clknet_leaf_218_clk _02343_ VGND VGND VPWR VPWR datamem.data_ram\[52\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_22390_ _09392_ VGND VGND VPWR VPWR _09552_ sky130_fd_sc_hd__buf_4
XFILLER_0_45_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31588_ clknet_leaf_57_clk net1187 VGND VGND VPWR VPWR rvcpu.dp.plmw.PCPlus4W\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21341_ rvcpu.ALUResultE\[10\] rvcpu.ALUResultE\[12\] rvcpu.ALUResultE\[16\] _08602_
+ VGND VGND VPWR VPWR _08603_ sky130_fd_sc_hd__or4_1
X_23256__903 clknet_1_0__leaf__10127_ VGND VGND VPWR VPWR net1029 sky130_fd_sc_hd__inv_2
XFILLER_0_5_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30539_ clknet_leaf_195_clk _02274_ VGND VGND VPWR VPWR datamem.data_ram\[55\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold610 datamem.data_ram\[30\]\[0\] VGND VGND VPWR VPWR net1760 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21272_ _08533_ VGND VGND VPWR VPWR _08534_ sky130_fd_sc_hd__buf_6
XFILLER_0_102_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold621 datamem.data_ram\[8\]\[4\] VGND VGND VPWR VPWR net1771 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_229_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold632 datamem.data_ram\[16\]\[0\] VGND VGND VPWR VPWR net1782 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_237_clk clknet_5_20__leaf_clk VGND VGND VPWR VPWR clknet_leaf_237_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold643 datamem.data_ram\[8\]\[0\] VGND VGND VPWR VPWR net1793 sky130_fd_sc_hd__dlygate4sd3_1
X_20223_ datamem.data_ram\[16\]\[3\] _07138_ _07514_ _07515_ VGND VGND VPWR VPWR _07516_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_124_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32209_ clknet_leaf_241_clk _03631_ VGND VGND VPWR VPWR datamem.data_ram\[36\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold654 datamem.data_ram\[26\]\[5\] VGND VGND VPWR VPWR net1804 sky130_fd_sc_hd__dlygate4sd3_1
Xhold665 rvcpu.dp.plfd.PCD\[16\] VGND VGND VPWR VPWR net1815 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold676 datamem.data_ram\[34\]\[5\] VGND VGND VPWR VPWR net1826 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_204_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_228_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold687 datamem.data_ram\[52\]\[0\] VGND VGND VPWR VPWR net1837 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold698 datamem.data_ram\[52\]\[5\] VGND VGND VPWR VPWR net1848 sky130_fd_sc_hd__dlygate4sd3_1
X_20154_ datamem.data_ram\[52\]\[27\] _07230_ _07443_ _07446_ VGND VGND VPWR VPWR
+ _07447_ sky130_fd_sc_hd__o211a_1
Xhold2000 datamem.data_ram\[25\]\[8\] VGND VGND VPWR VPWR net3150 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2011 datamem.data_ram\[16\]\[8\] VGND VGND VPWR VPWR net3161 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2022 datamem.data_ram\[31\]\[27\] VGND VGND VPWR VPWR net3172 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27750_ _12314_ VGND VGND VPWR VPWR _03725_ sky130_fd_sc_hd__clkbuf_1
Xhold2033 rvcpu.dp.rf.reg_file_arr\[26\]\[11\] VGND VGND VPWR VPWR net3183 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2044 datamem.data_ram\[26\]\[21\] VGND VGND VPWR VPWR net3194 sky130_fd_sc_hd__dlygate4sd3_1
X_24962_ _10700_ VGND VGND VPWR VPWR _02551_ sky130_fd_sc_hd__clkbuf_1
X_20085_ datamem.data_ram\[53\]\[10\] _06823_ _06670_ datamem.data_ram\[55\]\[10\]
+ VGND VGND VPWR VPWR _07379_ sky130_fd_sc_hd__o22a_1
XFILLER_0_176_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2055 rvcpu.dp.rf.reg_file_arr\[12\]\[26\] VGND VGND VPWR VPWR net3205 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1310 datamem.data_ram\[63\]\[27\] VGND VGND VPWR VPWR net2460 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1321 rvcpu.dp.rf.reg_file_arr\[15\]\[21\] VGND VGND VPWR VPWR net2471 sky130_fd_sc_hd__dlygate4sd3_1
X_26701_ _11705_ VGND VGND VPWR VPWR _03285_ sky130_fd_sc_hd__clkbuf_1
Xhold2066 datamem.data_ram\[3\]\[12\] VGND VGND VPWR VPWR net3216 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2077 datamem.data_ram\[48\]\[24\] VGND VGND VPWR VPWR net3227 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1332 datamem.data_ram\[60\]\[29\] VGND VGND VPWR VPWR net2482 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1343 rvcpu.dp.rf.reg_file_arr\[4\]\[23\] VGND VGND VPWR VPWR net2493 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2088 rvcpu.dp.rf.reg_file_arr\[29\]\[5\] VGND VGND VPWR VPWR net3238 sky130_fd_sc_hd__dlygate4sd3_1
X_27681_ _12277_ VGND VGND VPWR VPWR _03693_ sky130_fd_sc_hd__clkbuf_1
X_24893_ _10663_ VGND VGND VPWR VPWR _02519_ sky130_fd_sc_hd__clkbuf_1
Xhold1354 rvcpu.dp.rf.reg_file_arr\[27\]\[5\] VGND VGND VPWR VPWR net2504 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_212_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2099 datamem.data_ram\[25\]\[28\] VGND VGND VPWR VPWR net3249 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29420_ clknet_leaf_12_clk _01155_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD2E\[31\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__10201_ clknet_0__10201_ VGND VGND VPWR VPWR clknet_1_1__leaf__10201_
+ sky130_fd_sc_hd__clkbuf_16
Xhold1365 datamem.data_ram\[57\]\[24\] VGND VGND VPWR VPWR net2515 sky130_fd_sc_hd__dlygate4sd3_1
X_26632_ _07808_ _10946_ _11494_ VGND VGND VPWR VPWR _11661_ sky130_fd_sc_hd__or3_1
Xhold1376 rvcpu.dp.rf.reg_file_arr\[7\]\[16\] VGND VGND VPWR VPWR net2526 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1387 rvcpu.dp.rf.reg_file_arr\[31\]\[3\] VGND VGND VPWR VPWR net2537 sky130_fd_sc_hd__dlygate4sd3_1
X_23844_ _10218_ VGND VGND VPWR VPWR _01915_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_505 _11946_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1398 datamem.data_ram\[34\]\[20\] VGND VGND VPWR VPWR net2548 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_516 _13223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_185_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_527 _13319_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29351_ clknet_leaf_145_clk _01086_ VGND VGND VPWR VPWR datamem.data_ram\[61\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__10132_ clknet_0__10132_ VGND VGND VPWR VPWR clknet_1_1__leaf__10132_
+ sky130_fd_sc_hd__clkbuf_16
X_26563_ _11626_ VGND VGND VPWR VPWR _03226_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_538 clknet_1_1__leaf__10087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20987_ datamem.data_ram\[9\]\[15\] _06653_ _08275_ _06597_ VGND VGND VPWR VPWR _08276_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_549 _06790_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_212_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28302_ _12624_ VGND VGND VPWR VPWR _03967_ sky130_fd_sc_hd__clkbuf_1
X_25514_ _10991_ net1502 _11009_ _11013_ VGND VGND VPWR VPWR _02790_ sky130_fd_sc_hd__a31o_1
XFILLER_0_165_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22726_ _09636_ _09867_ _09869_ _09510_ VGND VGND VPWR VPWR _09870_ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29282_ _13162_ VGND VGND VPWR VPWR _04409_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_211_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_644 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28233_ _12435_ net2876 _12583_ VGND VGND VPWR VPWR _12586_ sky130_fd_sc_hd__mux2_1
XFILLER_0_193_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25445_ _07122_ VGND VGND VPWR VPWR _10979_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_137_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22657_ _09412_ _09800_ _09802_ _09804_ _09413_ VGND VGND VPWR VPWR _09805_ sky130_fd_sc_hd__a221o_1
XFILLER_0_211_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_188_5009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21608_ _08682_ _08855_ _08858_ VGND VGND VPWR VPWR _08859_ sky130_fd_sc_hd__a21o_1
XFILLER_0_153_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28164_ _12361_ net3835 _12546_ VGND VGND VPWR VPWR _12549_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_213_5599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25376_ _10410_ _10936_ VGND VGND VPWR VPWR _10940_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_170_4570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22588_ rvcpu.dp.rf.reg_file_arr\[0\]\[14\] rvcpu.dp.rf.reg_file_arr\[1\]\[14\] rvcpu.dp.rf.reg_file_arr\[2\]\[14\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[14\] _09477_ _09466_ VGND VGND VPWR VPWR _09740_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_170_4581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27115_ _11918_ VGND VGND VPWR VPWR _11956_ sky130_fd_sc_hd__buf_2
XFILLER_0_62_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24327_ _09236_ net4236 _10338_ VGND VGND VPWR VPWR _10340_ sky130_fd_sc_hd__mux2_1
X_21539_ _08572_ _08792_ VGND VGND VPWR VPWR _08793_ sky130_fd_sc_hd__or2_1
X_28095_ _12512_ VGND VGND VPWR VPWR _03872_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15060_ _13397_ _13387_ _13390_ VGND VGND VPWR VPWR _13607_ sky130_fd_sc_hd__and3_2
X_27046_ _11904_ net1850 _11910_ _11913_ VGND VGND VPWR VPWR _03422_ sky130_fd_sc_hd__a31o_1
X_24258_ _10301_ VGND VGND VPWR VPWR _02246_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_226_5916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_226_5927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_147_4016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_228_clk clknet_5_20__leaf_clk VGND VGND VPWR VPWR clknet_leaf_228_clk
+ sky130_fd_sc_hd__clkbuf_8
X_22979__686 clknet_1_0__leaf__10083_ VGND VGND VPWR VPWR net812 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_147_4027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_222_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28997_ _07077_ _10932_ _10918_ VGND VGND VPWR VPWR _13008_ sky130_fd_sc_hd__or3_1
X_18750_ _05782_ _05936_ _05950_ _05776_ _06100_ VGND VGND VPWR VPWR _06101_ sky130_fd_sc_hd__o221a_1
X_27948_ _12426_ VGND VGND VPWR VPWR _03811_ sky130_fd_sc_hd__clkbuf_1
X_15962_ net2347 _13201_ _14311_ VGND VGND VPWR VPWR _14318_ sky130_fd_sc_hd__mux2_1
XFILLER_0_219_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_218_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold3290 rvcpu.dp.rf.reg_file_arr\[24\]\[6\] VGND VGND VPWR VPWR net4440 sky130_fd_sc_hd__dlygate4sd3_1
X_17701_ _13201_ net2354 _05118_ VGND VGND VPWR VPWR _05125_ sky130_fd_sc_hd__mux2_1
X_14913_ _13365_ VGND VGND VPWR VPWR _13463_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_222_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18681_ _05239_ _06016_ _06021_ _06035_ VGND VGND VPWR VPWR rvcpu.ALUResultE\[9\]
+ sky130_fd_sc_hd__a211o_2
XTAP_TAPCELL_ROW_106_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27879_ _12388_ VGND VGND VPWR VPWR _03780_ sky130_fd_sc_hd__clkbuf_1
X_15893_ _14281_ VGND VGND VPWR VPWR _02078_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_106_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17632_ _05088_ VGND VGND VPWR VPWR _01222_ sky130_fd_sc_hd__clkbuf_1
X_29618_ net972 _01353_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[25\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_14844_ _13296_ VGND VGND VPWR VPWR _13397_ sky130_fd_sc_hd__buf_4
X_30890_ clknet_leaf_216_clk _02625_ VGND VGND VPWR VPWR datamem.data_ram\[42\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_177_4735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_177_4746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17563_ _13198_ net3741 _05046_ VGND VGND VPWR VPWR _05052_ sky130_fd_sc_hd__mux2_1
X_29549_ net903 _01284_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[27\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_14775_ _13282_ VGND VGND VPWR VPWR _13328_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_67_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19302_ _06597_ VGND VGND VPWR VPWR _06598_ sky130_fd_sc_hd__buf_6
X_16514_ net2739 _14474_ _04489_ VGND VGND VPWR VPWR _04495_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32560_ clknet_leaf_183_clk _03982_ VGND VGND VPWR VPWR datamem.data_ram\[22\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17494_ _05015_ VGND VGND VPWR VPWR _01295_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23737__328 clknet_1_0__leaf__10199_ VGND VGND VPWR VPWR net454 sky130_fd_sc_hd__inv_2
XFILLER_0_168_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31511_ clknet_leaf_52_clk net1183 VGND VGND VPWR VPWR rvcpu.dp.plem.PCPlus4M\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_19233_ _06538_ rvcpu.dp.plde.ImmExtE\[27\] _06493_ VGND VGND VPWR VPWR _06539_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16445_ _04457_ VGND VGND VPWR VPWR _01818_ sky130_fd_sc_hd__clkbuf_1
X_32491_ clknet_leaf_79_clk _03913_ VGND VGND VPWR VPWR datamem.data_ram\[25\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19164_ _06478_ net4363 _06419_ VGND VGND VPWR VPWR _06479_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_136_3753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31442_ clknet_leaf_5_clk rvcpu.dp.SrcBFW_Mux.y\[0\] VGND VGND VPWR VPWR rvcpu.dp.plem.WriteDataM\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_136_3764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16376_ net2129 _14474_ _14547_ VGND VGND VPWR VPWR _14553_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18115_ _05461_ _05467_ _05473_ _05481_ VGND VGND VPWR VPWR _05482_ sky130_fd_sc_hd__and4_1
XFILLER_0_143_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15327_ _13608_ _13578_ VGND VGND VPWR VPWR _13864_ sky130_fd_sc_hd__nand2_1
X_19095_ _06415_ _06417_ VGND VGND VPWR VPWR _06418_ sky130_fd_sc_hd__xnor2_1
X_31373_ clknet_leaf_18_clk _03076_ VGND VGND VPWR VPWR rvcpu.dp.plde.ImmExtE\[22\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f__10221_ clknet_0__10221_ VGND VGND VPWR VPWR clknet_1_0__leaf__10221_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18046_ rvcpu.dp.plde.ImmExtE\[10\] rvcpu.dp.SrcBFW_Mux.y\[10\] _05278_ VGND VGND
+ VPWR VPWR _05415_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30324_ net670 _02059_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[4\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_15258_ _13291_ _13337_ _13797_ VGND VGND VPWR VPWR _13798_ sky130_fd_sc_hd__or3b_1
Xclkbuf_1_0__f__10152_ clknet_0__10152_ VGND VGND VPWR VPWR clknet_1_0__leaf__10152_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_111_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_219_clk clknet_5_21__leaf_clk VGND VGND VPWR VPWR clknet_leaf_219_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_112_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30255_ net609 _01990_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[6\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_15189_ _13726_ _13727_ _13730_ _13731_ VGND VGND VPWR VPWR _13732_ sky130_fd_sc_hd__or4_1
XFILLER_0_22_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__10083_ clknet_0__10083_ VGND VGND VPWR VPWR clknet_1_0__leaf__10083_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_39_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19997_ datamem.data_ram\[17\]\[2\] _06947_ _07290_ _06851_ VGND VGND VPWR VPWR _07291_
+ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_35_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30186_ net540 _01921_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[8\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_226_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_225_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18948_ _05548_ _05785_ VGND VGND VPWR VPWR _06286_ sky130_fd_sc_hd__nor2_1
X_23286__929 clknet_1_1__leaf__10131_ VGND VGND VPWR VPWR net1055 sky130_fd_sc_hd__inv_2
XFILLER_0_225_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18879_ _06136_ _05937_ VGND VGND VPWR VPWR _06222_ sky130_fd_sc_hd__nor2_1
XFILLER_0_146_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23898__457 clknet_1_0__leaf__10223_ VGND VGND VPWR VPWR net583 sky130_fd_sc_hd__inv_2
XFILLER_0_94_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20910_ datamem.data_ram\[17\]\[22\] _07833_ _07840_ VGND VGND VPWR VPWR _08200_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_146_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21890_ _09117_ _09121_ _09125_ _08624_ VGND VGND VPWR VPWR _01054_ sky130_fd_sc_hd__o31a_1
XFILLER_0_179_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24117__624 clknet_1_1__leaf__10259_ VGND VGND VPWR VPWR net750 sky130_fd_sc_hd__inv_2
XFILLER_0_179_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32827_ clknet_leaf_164_clk _04249_ VGND VGND VPWR VPWR datamem.data_ram\[12\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_20841_ datamem.data_ram\[26\]\[14\] _07203_ _07077_ datamem.data_ram\[27\]\[14\]
+ _08130_ VGND VGND VPWR VPWR _08131_ sky130_fd_sc_hd__o221a_1
XFILLER_0_178_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20772_ datamem.data_ram\[62\]\[6\] _07833_ _08061_ _07840_ VGND VGND VPWR VPWR _08062_
+ sky130_fd_sc_hd__a211o_1
X_32758_ clknet_leaf_160_clk _04180_ VGND VGND VPWR VPWR datamem.data_ram\[15\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_193_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22511_ rvcpu.dp.rf.reg_file_arr\[4\]\[10\] rvcpu.dp.rf.reg_file_arr\[5\]\[10\] rvcpu.dp.rf.reg_file_arr\[6\]\[10\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[10\] _09478_ _09479_ VGND VGND VPWR VPWR _09667_
+ sky130_fd_sc_hd__mux4_1
X_31709_ clknet_leaf_31_clk _03167_ VGND VGND VPWR VPWR rvcpu.dp.pcreg.q\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32689_ clknet_leaf_251_clk _04111_ VGND VGND VPWR VPWR datamem.data_ram\[18\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_175_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25230_ _10854_ VGND VGND VPWR VPWR _02665_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22442_ _09599_ _09600_ _09380_ VGND VGND VPWR VPWR _09601_ sky130_fd_sc_hd__mux2_2
XFILLER_0_73_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25161_ _09305_ VGND VGND VPWR VPWR _10814_ sky130_fd_sc_hd__buf_2
XFILLER_0_190_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22373_ _09534_ _09535_ VGND VGND VPWR VPWR _09536_ sky130_fd_sc_hd__and2_1
XFILLER_0_161_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_206_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21324_ _08580_ rvcpu.dp.plde.RdE\[0\] _08582_ rvcpu.dp.plfd.InstrD\[18\] VGND VGND
+ VPWR VPWR _08586_ sky130_fd_sc_hd__o22a_1
XFILLER_0_66_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25092_ _10777_ _10051_ VGND VGND VPWR VPWR _10778_ sky130_fd_sc_hd__nand2_4
XFILLER_0_5_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_206_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28920_ _12965_ VGND VGND VPWR VPWR _04244_ sky130_fd_sc_hd__clkbuf_1
Xhold440 datamem.data_ram\[49\]\[2\] VGND VGND VPWR VPWR net1590 sky130_fd_sc_hd__dlygate4sd3_1
X_21255_ _08516_ VGND VGND VPWR VPWR _08517_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_41_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold451 datamem.data_ram\[7\]\[0\] VGND VGND VPWR VPWR net1601 sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 datamem.data_ram\[29\]\[0\] VGND VGND VPWR VPWR net1612 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold473 rvcpu.dp.plfd.PCPlus4D\[6\] VGND VGND VPWR VPWR net1623 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20206_ datamem.data_ram\[54\]\[11\] _06743_ _07242_ datamem.data_ram\[49\]\[11\]
+ VGND VGND VPWR VPWR _07499_ sky130_fd_sc_hd__o22a_1
Xhold484 datamem.data_ram\[32\]\[4\] VGND VGND VPWR VPWR net1634 sky130_fd_sc_hd__dlygate4sd3_1
X_28851_ _12745_ net2982 _12923_ VGND VGND VPWR VPWR _12929_ sky130_fd_sc_hd__mux2_1
Xhold495 datamem.data_ram\[16\]\[6\] VGND VGND VPWR VPWR net1645 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_221_5802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21186_ _08471_ _08472_ VGND VGND VPWR VPWR _08473_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_217_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27802_ _12138_ net2269 _12336_ VGND VGND VPWR VPWR _12343_ sky130_fd_sc_hd__mux2_1
X_20137_ datamem.data_ram\[37\]\[27\] _06815_ _07428_ _07429_ VGND VGND VPWR VPWR
+ _07430_ sky130_fd_sc_hd__o211a_1
X_28782_ _12892_ VGND VGND VPWR VPWR _04179_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25994_ _08572_ _11315_ _11312_ _11321_ VGND VGND VPWR VPWR _02962_ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_216_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27733_ _12305_ VGND VGND VPWR VPWR _03717_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_216_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24945_ _10691_ VGND VGND VPWR VPWR _02543_ sky130_fd_sc_hd__clkbuf_1
X_20068_ datamem.data_ram\[54\]\[26\] _06625_ _06631_ datamem.data_ram\[51\]\[26\]
+ VGND VGND VPWR VPWR _07362_ sky130_fd_sc_hd__o22a_1
Xhold1140 datamem.data_ram\[60\]\[27\] VGND VGND VPWR VPWR net2290 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1151 datamem.data_ram\[38\]\[26\] VGND VGND VPWR VPWR net2301 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1162 rvcpu.dp.rf.reg_file_arr\[2\]\[31\] VGND VGND VPWR VPWR net2312 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1173 rvcpu.dp.rf.reg_file_arr\[9\]\[25\] VGND VGND VPWR VPWR net2323 sky130_fd_sc_hd__dlygate4sd3_1
X_27664_ _12268_ VGND VGND VPWR VPWR _03685_ sky130_fd_sc_hd__clkbuf_1
X_24876_ _10654_ VGND VGND VPWR VPWR _02511_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_213_854 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1184 datamem.data_ram\[40\]\[15\] VGND VGND VPWR VPWR net2334 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29403_ clknet_leaf_0_clk _01138_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD2E\[14\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_302 _14127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1195 rvcpu.dp.rf.reg_file_arr\[4\]\[16\] VGND VGND VPWR VPWR net2345 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_219_5742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26615_ _11655_ VGND VGND VPWR VPWR _03249_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_313 _14177_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_219_5753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23827_ _07136_ VGND VGND VPWR VPWR _10209_ sky130_fd_sc_hd__buf_8
XANTENNA_324 _14447_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_206_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27595_ _12231_ VGND VGND VPWR VPWR _03653_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_335 _14461_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_346 clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_200_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_184_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_357 rvcpu.dp.SrcBFW_Mux.y\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29334_ clknet_leaf_176_clk _01069_ VGND VGND VPWR VPWR datamem.data_ram\[62\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_26546_ _11091_ _11610_ VGND VGND VPWR VPWR _11617_ sky130_fd_sc_hd__and2_1
XANTENNA_368 rvcpu.dp.plde.ImmExtE\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_379 rvcpu.dp.plmw.ReadDataW\[29\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_4621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_4632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29265_ _13153_ VGND VGND VPWR VPWR _04401_ sky130_fd_sc_hd__clkbuf_1
X_22709_ _09495_ _09853_ VGND VGND VPWR VPWR _09854_ sky130_fd_sc_hd__nor2_1
X_26477_ net1823 _11268_ _11596_ _10041_ VGND VGND VPWR VPWR _03170_ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23689_ clknet_1_0__leaf__10192_ VGND VGND VPWR VPWR _10195_ sky130_fd_sc_hd__buf_1
XFILLER_0_165_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16230_ _13256_ VGND VGND VPWR VPWR _14472_ sky130_fd_sc_hd__buf_4
X_28216_ _12361_ net3772 net45 VGND VGND VPWR VPWR _12577_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25428_ _10520_ _10630_ _10828_ VGND VGND VPWR VPWR _10970_ sky130_fd_sc_hd__a21oi_4
X_29196_ _09313_ net3519 _13112_ VGND VGND VPWR VPWR _13116_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28147_ _12452_ net3681 net73 VGND VGND VPWR VPWR _12540_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16161_ _14425_ VGND VGND VPWR VPWR _01946_ sky130_fd_sc_hd__clkbuf_1
X_25359_ _10876_ net1409 _10920_ _10928_ VGND VGND VPWR VPWR _02720_ sky130_fd_sc_hd__a31o_1
Xclkload18 clknet_5_22__leaf_clk VGND VGND VPWR VPWR clkload18/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload29 clknet_leaf_19_clk VGND VGND VPWR VPWR clkload29/Y sky130_fd_sc_hd__inv_6
X_15112_ _13348_ _13656_ VGND VGND VPWR VPWR _13657_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_499 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28078_ _12503_ VGND VGND VPWR VPWR _03864_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_131_3650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16092_ net2310 _13187_ _14385_ VGND VGND VPWR VPWR _14388_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27029_ _11829_ _11899_ VGND VGND VPWR VPWR _11903_ sky130_fd_sc_hd__and2_1
X_15043_ _13336_ _13472_ _13589_ VGND VGND VPWR VPWR _13590_ sky130_fd_sc_hd__a21oi_2
X_19920_ datamem.data_ram\[61\]\[17\] _07037_ _06837_ datamem.data_ram\[56\]\[17\]
+ VGND VGND VPWR VPWR _07215_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_71_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_166_4469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19851_ _07143_ _07145_ VGND VGND VPWR VPWR _07146_ sky130_fd_sc_hd__or2_1
X_30040_ net402 _01775_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[13\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23423__75 clknet_1_1__leaf__10154_ VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__inv_2
X_23170__842 clknet_1_0__leaf__10110_ VGND VGND VPWR VPWR net968 sky130_fd_sc_hd__inv_2
XFILLER_0_208_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18802_ _06134_ _05809_ _06135_ _06149_ VGND VGND VPWR VPWR _06150_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_101_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19782_ _06863_ VGND VGND VPWR VPWR _07077_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_207_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16994_ _04749_ VGND VGND VPWR VPWR _01545_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_129_3590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18733_ _06055_ _06070_ _06076_ _06084_ VGND VGND VPWR VPWR rvcpu.ALUResultE\[12\]
+ sky130_fd_sc_hd__a211o_1
X_15945_ _14308_ VGND VGND VPWR VPWR _02053_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_30_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31991_ clknet_leaf_127_clk _03413_ VGND VGND VPWR VPWR datamem.data_ram\[31\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_223_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30942_ clknet_leaf_96_clk _02677_ VGND VGND VPWR VPWR datamem.data_ram\[3\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_18664_ _05997_ _05599_ _06017_ _06018_ VGND VGND VPWR VPWR _06019_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_125_3487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15876_ _14270_ VGND VGND VPWR VPWR _02084_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_125_3498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17615_ _13275_ net3686 _05045_ VGND VGND VPWR VPWR _05079_ sky130_fd_sc_hd__mux2_1
X_14827_ _13286_ _13288_ VGND VGND VPWR VPWR _13380_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30873_ clknet_leaf_57_clk _02608_ VGND VGND VPWR VPWR datamem.data_ram\[42\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_18595_ _05886_ _05932_ _05953_ VGND VGND VPWR VPWR rvcpu.ALUResultE\[5\] sky130_fd_sc_hd__o21ai_4
XFILLER_0_99_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23971__507 clknet_1_0__leaf__10238_ VGND VGND VPWR VPWR net633 sky130_fd_sc_hd__inv_2
X_32612_ clknet_leaf_80_clk _04034_ VGND VGND VPWR VPWR datamem.data_ram\[20\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17546_ _05042_ VGND VGND VPWR VPWR _01270_ sky130_fd_sc_hd__clkbuf_1
X_14758_ rvcpu.dp.pcreg.q\[8\] VGND VGND VPWR VPWR _13311_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_138_3815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32543_ clknet_leaf_85_clk _03965_ VGND VGND VPWR VPWR datamem.data_ram\[23\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_28_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_184_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17477_ _14191_ net4284 _04996_ VGND VGND VPWR VPWR _05006_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14689_ net2059 _13251_ _13245_ VGND VGND VPWR VPWR _13252_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19216_ _06522_ _06523_ VGND VGND VPWR VPWR _06524_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16428_ _14580_ VGND VGND VPWR VPWR _01826_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_60_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32474_ clknet_leaf_258_clk _03896_ VGND VGND VPWR VPWR datamem.data_ram\[26\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_60_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_536 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19147_ rvcpu.dp.plde.ImmExtE\[17\] rvcpu.dp.plde.PCE\[17\] VGND VGND VPWR VPWR _06463_
+ sky130_fd_sc_hd__nor2_1
X_31425_ clknet_leaf_60_clk _03128_ VGND VGND VPWR VPWR datamem.data_ram\[44\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16359_ net3783 _14457_ _14536_ VGND VGND VPWR VPWR _14544_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19078_ _06396_ _06397_ _06394_ VGND VGND VPWR VPWR _06403_ sky130_fd_sc_hd__o21ai_2
X_31356_ clknet_leaf_22_clk _03059_ VGND VGND VPWR VPWR rvcpu.dp.plde.ImmExtE\[5\]
+ sky130_fd_sc_hd__dfxtp_2
Xclkbuf_1_0__f__10204_ clknet_0__10204_ VGND VGND VPWR VPWR clknet_1_0__leaf__10204_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_112_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18029_ _05398_ _05382_ VGND VGND VPWR VPWR _05399_ sky130_fd_sc_hd__nor2_1
X_30307_ net653 _02042_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[5\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31287_ clknet_leaf_108_clk _02990_ VGND VGND VPWR VPWR datamem.data_ram\[34\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__10135_ clknet_0__10135_ VGND VGND VPWR VPWR clknet_1_0__leaf__10135_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_58_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21040_ _07838_ _08327_ _08328_ VGND VGND VPWR VPWR _08329_ sky130_fd_sc_hd__or3_1
XFILLER_0_199_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30238_ net592 _01973_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[7\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_226_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30169_ net531 _01904_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[0\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_226_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24730_ _10444_ net4058 _10571_ VGND VGND VPWR VPWR _10574_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21942_ rvcpu.dp.rf.reg_file_arr\[8\]\[29\] rvcpu.dp.rf.reg_file_arr\[10\]\[29\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[29\] rvcpu.dp.rf.reg_file_arr\[11\]\[29\] _08649_
+ _08561_ VGND VGND VPWR VPWR _09175_ sky130_fd_sc_hd__mux4_1
XFILLER_0_59_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24661_ _10413_ _10532_ VGND VGND VPWR VPWR _10536_ sky130_fd_sc_hd__and2_1
X_23147__822 clknet_1_1__leaf__10107_ VGND VGND VPWR VPWR net948 sky130_fd_sc_hd__inv_2
X_21873_ rvcpu.dp.rf.reg_file_arr\[16\]\[26\] rvcpu.dp.rf.reg_file_arr\[17\]\[26\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[26\] rvcpu.dp.rf.reg_file_arr\[19\]\[26\] _08631_
+ _08632_ VGND VGND VPWR VPWR _09109_ sky130_fd_sc_hd__mux4_1
X_26400_ _11535_ rvcpu.ALUResultE\[7\] VGND VGND VPWR VPWR _11543_ sky130_fd_sc_hd__and2_1
XFILLER_0_221_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20824_ _08112_ _08113_ _07837_ VGND VGND VPWR VPWR _08114_ sky130_fd_sc_hd__a21o_1
X_27380_ _12109_ VGND VGND VPWR VPWR _03560_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_171_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24592_ _10396_ net3149 _10491_ VGND VGND VPWR VPWR _10497_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26331_ _11353_ net1718 _11496_ _11500_ VGND VGND VPWR VPWR _03120_ sky130_fd_sc_hd__a31o_1
XFILLER_0_147_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20755_ _08041_ _08043_ _08044_ VGND VGND VPWR VPWR _08045_ sky130_fd_sc_hd__or3_2
XFILLER_0_9_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23340__978 clknet_1_0__leaf__10136_ VGND VGND VPWR VPWR net1104 sky130_fd_sc_hd__inv_2
XFILLER_0_108_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29050_ _13018_ net1730 _13030_ _13038_ VGND VGND VPWR VPWR _04301_ sky130_fd_sc_hd__a31o_1
X_26262_ net1284 _11432_ VGND VGND VPWR VPWR _11463_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_210_5525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20686_ datamem.data_ram\[52\]\[5\] _06955_ _06948_ datamem.data_ram\[49\]\[5\] VGND
+ VGND VPWR VPWR _07977_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_718 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_210_5536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_210_5547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28001_ _12461_ VGND VGND VPWR VPWR _03829_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25213_ _10845_ VGND VGND VPWR VPWR _02657_ sky130_fd_sc_hd__clkbuf_1
X_22425_ _09418_ VGND VGND VPWR VPWR _09585_ sky130_fd_sc_hd__clkbuf_4
X_26193_ rvcpu.ALUControl\[2\] _11432_ VGND VGND VPWR VPWR _11434_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25144_ _10804_ VGND VGND VPWR VPWR _02629_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_149_Right_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22356_ _09516_ _09518_ VGND VGND VPWR VPWR _09519_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21307_ _08568_ VGND VGND VPWR VPWR _08569_ sky130_fd_sc_hd__buf_4
XFILLER_0_14_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29952_ net322 _01687_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[15\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_25075_ _10724_ net2781 net89 VGND VGND VPWR VPWR _10769_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22287_ _09451_ VGND VGND VPWR VPWR _09452_ sky130_fd_sc_hd__buf_4
XFILLER_0_104_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28903_ _12956_ VGND VGND VPWR VPWR _04236_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_208_5476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold270 datamem.data_ram\[21\]\[3\] VGND VGND VPWR VPWR net1420 sky130_fd_sc_hd__dlygate4sd3_1
X_21238_ datamem.data_ram\[52\]\[5\] datamem.data_ram\[53\]\[5\] _08499_ _08500_ VGND
+ VGND VPWR VPWR _08501_ sky130_fd_sc_hd__or4b_2
XFILLER_0_104_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29883_ net261 _01618_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[17\]\[14\] sky130_fd_sc_hd__dfxtp_1
Xhold281 datamem.data_ram\[30\]\[2\] VGND VGND VPWR VPWR net1431 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_208_5487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_208_5498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold292 datamem.data_ram\[12\]\[7\] VGND VGND VPWR VPWR net1442 sky130_fd_sc_hd__dlygate4sd3_1
X_28834_ _12762_ net3541 _12914_ VGND VGND VPWR VPWR _12920_ sky130_fd_sc_hd__mux2_1
X_23234__883 clknet_1_1__leaf__10125_ VGND VGND VPWR VPWR net1009 sky130_fd_sc_hd__inv_2
X_21169_ _06917_ _08457_ VGND VGND VPWR VPWR _08458_ sky130_fd_sc_hd__or2_1
XFILLER_0_218_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_161_4355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_4366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28765_ _12698_ net3173 _12877_ VGND VGND VPWR VPWR _12883_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_205_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25977_ net1762 _11302_ _11300_ _11311_ VGND VGND VPWR VPWR _02955_ sky130_fd_sc_hd__o211a_1
X_15730_ _13271_ VGND VGND VPWR VPWR _14191_ sky130_fd_sc_hd__buf_4
X_27716_ _12296_ VGND VGND VPWR VPWR _03709_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24928_ _10682_ VGND VGND VPWR VPWR _02535_ sky130_fd_sc_hd__clkbuf_1
X_28696_ _12846_ VGND VGND VPWR VPWR _04139_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_217_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27647_ _12140_ net2498 _12251_ VGND VGND VPWR VPWR _12259_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15661_ _14144_ VGND VGND VPWR VPWR _02181_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_110 _07031_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24859_ _10645_ VGND VGND VPWR VPWR _02503_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_213_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_185_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_121 _07226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17400_ _04965_ VGND VGND VPWR VPWR _01339_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_132 _07831_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_201_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14612_ _13170_ VGND VGND VPWR VPWR _13193_ sky130_fd_sc_hd__buf_4
XANTENNA_143 _07840_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18380_ rvcpu.dp.plde.unsignE _05284_ VGND VGND VPWR VPWR _05744_ sky130_fd_sc_hd__or2_1
XANTENNA_154 _08353_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15592_ net2066 _13213_ _14103_ VGND VGND VPWR VPWR _14104_ sky130_fd_sc_hd__mux2_1
X_27578_ _12222_ VGND VGND VPWR VPWR _03645_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_120_3384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_165 _08656_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_176 _08827_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29317_ clknet_leaf_11_clk _01052_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD1E\[24\] sky130_fd_sc_hd__dfxtp_1
X_17331_ net2280 _13256_ _04924_ VGND VGND VPWR VPWR _04929_ sky130_fd_sc_hd__mux2_1
XANTENNA_187 _09181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26529_ _11372_ _11606_ _02993_ VGND VGND VPWR VPWR _03212_ sky130_fd_sc_hd__a21o_1
XANTENNA_198 _09453_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_200_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0__10129_ _10129_ VGND VGND VPWR VPWR clknet_0__10129_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_154_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29248_ _13144_ VGND VGND VPWR VPWR _04393_ sky130_fd_sc_hd__clkbuf_1
X_17262_ _14181_ net2612 _04887_ VGND VGND VPWR VPWR _04892_ sky130_fd_sc_hd__mux2_1
XFILLER_0_193_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_181_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19001_ _05288_ _05289_ VGND VGND VPWR VPWR _06335_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16213_ _14460_ VGND VGND VPWR VPWR _01929_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_23_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29179_ _09243_ net3421 net63 VGND VGND VPWR VPWR _13107_ sky130_fd_sc_hd__mux2_1
X_17193_ _04855_ VGND VGND VPWR VPWR _01444_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_47 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload107 clknet_leaf_161_clk VGND VGND VPWR VPWR clkload107/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_141_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload118 clknet_leaf_100_clk VGND VGND VPWR VPWR clkload118/Y sky130_fd_sc_hd__inv_6
XFILLER_0_183_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31210_ clknet_leaf_33_clk _02913_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCPlus4D\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16144_ net3678 _13266_ _14407_ VGND VGND VPWR VPWR _14415_ sky130_fd_sc_hd__mux2_1
Xclkload129 clknet_leaf_257_clk VGND VGND VPWR VPWR clkload129/Y sky130_fd_sc_hd__clkinvlp_4
XPHY_EDGE_ROW_116_Right_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32190_ clknet_leaf_271_clk _03612_ VGND VGND VPWR VPWR datamem.data_ram\[37\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_94_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24146__650 clknet_1_1__leaf__10262_ VGND VGND VPWR VPWR net776 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_94_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23552__176 clknet_1_0__leaf__10174_ VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__inv_2
X_31141_ clknet_leaf_68_clk rvcpu.ALUResultE\[0\] VGND VGND VPWR VPWR rvcpu.dp.plem.ALUResultM\[0\]
+ sky130_fd_sc_hd__dfxtp_4
X_16075_ _14378_ VGND VGND VPWR VPWR _01985_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_224_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15026_ _13513_ VGND VGND VPWR VPWR _13573_ sky130_fd_sc_hd__clkbuf_4
X_19903_ datamem.data_ram\[14\]\[17\] _06683_ _06648_ datamem.data_ram\[8\]\[17\]
+ VGND VGND VPWR VPWR _07198_ sky130_fd_sc_hd__o22a_1
X_31072_ clknet_leaf_163_clk _02807_ VGND VGND VPWR VPWR datamem.data_ram\[9\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_30023_ net385 _01758_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[13\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_19834_ datamem.data_ram\[39\]\[1\] _07125_ _07126_ _07128_ VGND VGND VPWR VPWR _07129_
+ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_127_3538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_127_3549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1909 datamem.data_ram\[40\]\[21\] VGND VGND VPWR VPWR net3059 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16977_ _04740_ VGND VGND VPWR VPWR _01553_ sky130_fd_sc_hd__clkbuf_1
X_19765_ datamem.data_ram\[21\]\[25\] _06865_ _06672_ datamem.data_ram\[23\]\[25\]
+ _07059_ VGND VGND VPWR VPWR _07060_ sky130_fd_sc_hd__o221a_1
XFILLER_0_208_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_217_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18716_ _05239_ _06054_ _06068_ VGND VGND VPWR VPWR rvcpu.ALUResultE\[11\] sky130_fd_sc_hd__a21o_1
X_15928_ net1915 _13251_ _14297_ VGND VGND VPWR VPWR _14300_ sky130_fd_sc_hd__mux2_1
X_19696_ datamem.data_ram\[10\]\[0\] _06989_ _06990_ datamem.data_ram\[8\]\[0\] _06991_
+ VGND VGND VPWR VPWR _06992_ sky130_fd_sc_hd__a221o_1
XFILLER_0_190_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31974_ clknet_leaf_130_clk _03396_ VGND VGND VPWR VPWR datamem.data_ram\[54\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18647_ _05775_ _05780_ _06002_ _05805_ VGND VGND VPWR VPWR _06003_ sky130_fd_sc_hd__a211oi_1
X_30925_ clknet_leaf_155_clk _02660_ VGND VGND VPWR VPWR datamem.data_ram\[40\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_15859_ net1945 _13254_ _14258_ VGND VGND VPWR VPWR _14262_ sky130_fd_sc_hd__mux2_1
XFILLER_0_189_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18578_ _05935_ _05936_ _05696_ VGND VGND VPWR VPWR _05937_ sky130_fd_sc_hd__mux2_1
X_30856_ clknet_leaf_155_clk _02591_ VGND VGND VPWR VPWR datamem.data_ram\[43\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_188_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17529_ _13248_ net2733 _05032_ VGND VGND VPWR VPWR _05034_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30787_ clknet_leaf_134_clk _02522_ VGND VGND VPWR VPWR datamem.data_ram\[46\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_528 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20540_ _06944_ VGND VGND VPWR VPWR _07831_ sky130_fd_sc_hd__buf_6
X_32526_ clknet_leaf_250_clk _03948_ VGND VGND VPWR VPWR datamem.data_ram\[24\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20471_ datamem.data_ram\[43\]\[20\] _06635_ _07759_ _07762_ VGND VGND VPWR VPWR
+ _07763_ sky130_fd_sc_hd__o211a_1
X_32457_ clknet_leaf_230_clk _03879_ VGND VGND VPWR VPWR datamem.data_ram\[26\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_229_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22210_ _09288_ net2555 _09371_ VGND VGND VPWR VPWR _09378_ sky130_fd_sc_hd__mux2_1
X_31408_ clknet_leaf_31_clk _03111_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCE\[25\] sky130_fd_sc_hd__dfxtp_1
X_23190_ _09224_ net4318 _10115_ VGND VGND VPWR VPWR _10116_ sky130_fd_sc_hd__mux2_1
X_23177__848 clknet_1_1__leaf__10111_ VGND VGND VPWR VPWR net974 sky130_fd_sc_hd__inv_2
XFILLER_0_14_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32388_ clknet_leaf_232_clk _03810_ VGND VGND VPWR VPWR datamem.data_ram\[29\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22141_ _09260_ net4269 _09332_ VGND VGND VPWR VPWR _09340_ sky130_fd_sc_hd__mux2_1
X_31339_ clknet_leaf_13_clk _03042_ VGND VGND VPWR VPWR rvcpu.dp.plde.Rs1E\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_1052 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22072_ _09287_ VGND VGND VPWR VPWR _09288_ sky130_fd_sc_hd__buf_2
XFILLER_0_227_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25900_ _11155_ VGND VGND VPWR VPWR _11268_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21023_ datamem.data_ram\[27\]\[31\] _06729_ _06654_ datamem.data_ram\[25\]\[31\]
+ VGND VGND VPWR VPWR _08312_ sky130_fd_sc_hd__o22a_1
XFILLER_0_199_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26880_ _11679_ _11810_ VGND VGND VPWR VPWR _11812_ sky130_fd_sc_hd__and2_1
XFILLER_0_226_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25831_ _11206_ _11207_ _11216_ VGND VGND VPWR VPWR _11217_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_203_5362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23529__156 clknet_1_1__leaf__10171_ VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__inv_2
XFILLER_0_227_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_203_5373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28550_ _12687_ net4056 _12768_ VGND VGND VPWR VPWR _12769_ sky130_fd_sc_hd__mux2_1
X_25762_ _13463_ _13876_ _11162_ VGND VGND VPWR VPWR _11163_ sky130_fd_sc_hd__a21o_1
XFILLER_0_184_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27501_ _12147_ net3771 _12179_ VGND VGND VPWR VPWR _12182_ sky130_fd_sc_hd__mux2_1
X_24713_ _10564_ VGND VGND VPWR VPWR _02438_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_195_5174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28481_ _06997_ _10049_ _10921_ VGND VGND VPWR VPWR _12724_ sky130_fd_sc_hd__and3_2
X_21925_ _08817_ _09156_ _09158_ _08699_ VGND VGND VPWR VPWR _09159_ sky130_fd_sc_hd__a211o_1
X_25693_ _11105_ net1712 _11111_ _11118_ VGND VGND VPWR VPWR _02864_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_195_5185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27432_ _09259_ VGND VGND VPWR VPWR _12140_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_132_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_210_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24644_ _10394_ net3411 _10521_ VGND VGND VPWR VPWR _10526_ sky130_fd_sc_hd__mux2_1
X_21856_ rvcpu.dp.rf.reg_file_arr\[20\]\[25\] rvcpu.dp.rf.reg_file_arr\[21\]\[25\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[25\] rvcpu.dp.rf.reg_file_arr\[23\]\[25\] _08778_
+ _08825_ VGND VGND VPWR VPWR _09093_ sky130_fd_sc_hd__mux4_1
XFILLER_0_78_873 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_218_Right_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20807_ datamem.data_ram\[44\]\[30\] datamem.data_ram\[45\]\[30\] _07826_ VGND VGND
+ VPWR VPWR _08097_ sky130_fd_sc_hd__mux2_1
X_27363_ _12085_ net4106 _12097_ VGND VGND VPWR VPWR _12100_ sky130_fd_sc_hd__mux2_1
X_24575_ _10450_ net4143 _10482_ VGND VGND VPWR VPWR _10488_ sky130_fd_sc_hd__mux2_1
X_24015__547 clknet_1_1__leaf__10242_ VGND VGND VPWR VPWR net673 sky130_fd_sc_hd__inv_2
X_21787_ _08686_ _09027_ _08748_ VGND VGND VPWR VPWR _09028_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_203_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29102_ _09329_ net2177 _13058_ VGND VGND VPWR VPWR _13066_ sky130_fd_sc_hd__mux2_1
X_26314_ net1588 _11436_ VGND VGND VPWR VPWR _11490_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_203_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27294_ _11976_ _12054_ VGND VGND VPWR VPWR _12060_ sky130_fd_sc_hd__and2_1
X_20738_ datamem.data_ram\[32\]\[6\] _07122_ _08027_ _07868_ VGND VGND VPWR VPWR _08028_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_154_4181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_154_4192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29033_ _13028_ VGND VGND VPWR VPWR _04294_ sky130_fd_sc_hd__clkbuf_1
X_26245_ _11438_ _11458_ _11459_ _09479_ VGND VGND VPWR VPWR _03075_ sky130_fd_sc_hd__a2bb2o_1
X_20669_ datamem.data_ram\[53\]\[29\] _06823_ _06733_ _07959_ VGND VGND VPWR VPWR
+ _07960_ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_150_4089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22408_ _09469_ _09568_ VGND VGND VPWR VPWR _09569_ sky130_fd_sc_hd__or2_1
X_26176_ rvcpu.dp.plfd.InstrD\[24\] _11362_ VGND VGND VPWR VPWR _11425_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23388_ _09306_ net2476 _10143_ VGND VGND VPWR VPWR _10145_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_626 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25127_ _10795_ VGND VGND VPWR VPWR _02621_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22339_ rvcpu.dp.rf.reg_file_arr\[0\]\[2\] rvcpu.dp.rf.reg_file_arr\[1\]\[2\] rvcpu.dp.rf.reg_file_arr\[2\]\[2\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[2\] _09463_ _09466_ VGND VGND VPWR VPWR _09503_ sky130_fd_sc_hd__mux4_1
XFILLER_0_108_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_163_4406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_163_4417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25058_ _10757_ VGND VGND VPWR VPWR _02590_ sky130_fd_sc_hd__clkbuf_1
X_29935_ net305 _01670_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[16\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_16900_ net3674 _14451_ _04695_ VGND VGND VPWR VPWR _04700_ sky130_fd_sc_hd__mux2_1
X_17880_ rvcpu.dp.plde.Rs1E\[3\] rvcpu.dp.plmw.RdW\[3\] VGND VGND VPWR VPWR _05253_
+ sky130_fd_sc_hd__xor2_1
X_29866_ net244 _01601_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[18\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_228_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16831_ _04663_ VGND VGND VPWR VPWR _01622_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28817_ _12698_ net3230 _12905_ VGND VGND VPWR VPWR _12911_ sky130_fd_sc_hd__mux2_1
X_29797_ clknet_leaf_218_clk _01532_ VGND VGND VPWR VPWR datamem.data_ram\[59\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_219_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19550_ datamem.data_ram\[20\]\[24\] _06687_ _06844_ _06845_ VGND VGND VPWR VPWR
+ _06846_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_122_3413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16762_ net2838 _14449_ _04623_ VGND VGND VPWR VPWR _04627_ sky130_fd_sc_hd__mux2_1
X_28748_ _12745_ net2441 net41 VGND VGND VPWR VPWR _12874_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_122_3424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18501_ _05688_ _05684_ _05398_ VGND VGND VPWR VPWR _05863_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_122_3435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15713_ _14179_ net4185 _14173_ VGND VGND VPWR VPWR _14180_ sky130_fd_sc_hd__mux2_1
X_19481_ _06776_ VGND VGND VPWR VPWR _06777_ sky130_fd_sc_hd__buf_8
X_28679_ _12837_ VGND VGND VPWR VPWR _04131_ sky130_fd_sc_hd__clkbuf_1
X_16693_ _04590_ VGND VGND VPWR VPWR _01695_ sky130_fd_sc_hd__clkbuf_1
X_18432_ _05795_ VGND VGND VPWR VPWR rvcpu.ALUResultE\[0\] sky130_fd_sc_hd__buf_1
X_30710_ clknet_leaf_148_clk _02445_ VGND VGND VPWR VPWR datamem.data_ram\[49\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_15644_ _13183_ VGND VGND VPWR VPWR _14133_ sky130_fd_sc_hd__buf_4
XFILLER_0_38_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31690_ clknet_leaf_41_clk _03148_ VGND VGND VPWR VPWR rvcpu.dp.pcreg.q\[8\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_180_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_14_Left_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18363_ _05727_ VGND VGND VPWR VPWR _05728_ sky130_fd_sc_hd__clkbuf_4
X_30641_ clknet_leaf_192_clk _02376_ VGND VGND VPWR VPWR datamem.data_ram\[51\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15575_ net2008 _13187_ _14092_ VGND VGND VPWR VPWR _14095_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17314_ net4426 _13231_ _04913_ VGND VGND VPWR VPWR _04920_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18294_ rvcpu.dp.plde.ALUControlE\[0\] rvcpu.dp.plde.ALUControlE\[1\] VGND VGND VPWR
+ VPWR _05659_ sky130_fd_sc_hd__nand2_1
X_30572_ clknet_leaf_146_clk _02307_ VGND VGND VPWR VPWR datamem.data_ram\[54\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_23935__490 clknet_1_0__leaf__10227_ VGND VGND VPWR VPWR net616 sky130_fd_sc_hd__inv_2
XFILLER_0_12_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32311_ clknet_leaf_269_clk _03733_ VGND VGND VPWR VPWR datamem.data_ram\[32\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17245_ _14164_ net3885 _04876_ VGND VGND VPWR VPWR _04883_ sky130_fd_sc_hd__mux2_1
XFILLER_0_226_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_1063 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32242_ clknet_leaf_229_clk _03664_ VGND VGND VPWR VPWR datamem.data_ram\[34\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_17176_ _04846_ VGND VGND VPWR VPWR _01452_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16127_ net2851 _13241_ _14396_ VGND VGND VPWR VPWR _14406_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32173_ clknet_leaf_227_clk _03595_ VGND VGND VPWR VPWR datamem.data_ram\[37\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_23_Left_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31124_ clknet_leaf_109_clk _02859_ VGND VGND VPWR VPWR datamem.data_ram\[35\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_55_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3108 rvcpu.dp.rf.reg_file_arr\[11\]\[0\] VGND VGND VPWR VPWR net4258 sky130_fd_sc_hd__dlygate4sd3_1
X_16058_ _14369_ VGND VGND VPWR VPWR _01993_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3119 datamem.data_ram\[61\]\[23\] VGND VGND VPWR VPWR net4269 sky130_fd_sc_hd__dlygate4sd3_1
X_15009_ _13504_ _13551_ _13555_ _13556_ VGND VGND VPWR VPWR _13557_ sky130_fd_sc_hd__a211o_1
XFILLER_0_20_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31055_ clknet_leaf_93_clk _02790_ VGND VGND VPWR VPWR datamem.data_ram\[38\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2407 datamem.data_ram\[47\]\[10\] VGND VGND VPWR VPWR net3557 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2418 datamem.data_ram\[6\]\[20\] VGND VGND VPWR VPWR net3568 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2429 rvcpu.dp.rf.reg_file_arr\[28\]\[5\] VGND VGND VPWR VPWR net3579 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30006_ clknet_leaf_175_clk _01741_ VGND VGND VPWR VPWR datamem.data_ram\[59\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1706 rvcpu.dp.rf.reg_file_arr\[0\]\[29\] VGND VGND VPWR VPWR net2856 sky130_fd_sc_hd__dlygate4sd3_1
X_19817_ datamem.data_ram\[30\]\[9\] _06629_ _06620_ datamem.data_ram\[28\]\[9\] VGND
+ VGND VPWR VPWR _07112_ sky130_fd_sc_hd__o22a_1
Xhold1717 datamem.data_ram\[33\]\[12\] VGND VGND VPWR VPWR net2867 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1728 rvcpu.dp.rf.reg_file_arr\[20\]\[7\] VGND VGND VPWR VPWR net2878 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1739 rvcpu.dp.rf.reg_file_arr\[18\]\[11\] VGND VGND VPWR VPWR net2889 sky130_fd_sc_hd__dlygate4sd3_1
X_23977__513 clknet_1_1__leaf__10238_ VGND VGND VPWR VPWR net639 sky130_fd_sc_hd__inv_2
XFILLER_0_223_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19748_ datamem.data_ram\[47\]\[25\] _06725_ _06765_ datamem.data_ram\[44\]\[25\]
+ VGND VGND VPWR VPWR _07043_ sky130_fd_sc_hd__o22a_1
XFILLER_0_79_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_195_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19679_ datamem.data_ram\[53\]\[0\] _06970_ _06972_ _06974_ VGND VGND VPWR VPWR _06975_
+ sky130_fd_sc_hd__a211o_1
X_31957_ clknet_leaf_133_clk _03379_ VGND VGND VPWR VPWR datamem.data_ram\[55\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_32_Left_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_204_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21710_ rvcpu.dp.rf.reg_file_arr\[28\]\[17\] rvcpu.dp.rf.reg_file_arr\[30\]\[17\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[17\] rvcpu.dp.rf.reg_file_arr\[31\]\[17\] _08629_
+ _08683_ VGND VGND VPWR VPWR _08955_ sky130_fd_sc_hd__mux4_1
XFILLER_0_133_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22690_ rvcpu.dp.rf.reg_file_arr\[28\]\[20\] rvcpu.dp.rf.reg_file_arr\[30\]\[20\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[20\] rvcpu.dp.rf.reg_file_arr\[31\]\[20\] _09381_
+ _09423_ VGND VGND VPWR VPWR _09836_ sky130_fd_sc_hd__mux4_1
X_30908_ clknet_leaf_194_clk _02643_ VGND VGND VPWR VPWR datamem.data_ram\[41\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_31888_ clknet_leaf_113_clk _03342_ VGND VGND VPWR VPWR datamem.data_ram\[36\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21641_ _08795_ _08883_ _08885_ _08889_ _08808_ VGND VGND VPWR VPWR _08890_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_190_5060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30839_ clknet_leaf_241_clk _02574_ VGND VGND VPWR VPWR datamem.data_ram\[44\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_23795__380 clknet_1_0__leaf__10205_ VGND VGND VPWR VPWR net506 sky130_fd_sc_hd__inv_2
XFILLER_0_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21572_ rvcpu.dp.rf.reg_file_arr\[16\]\[10\] rvcpu.dp.rf.reg_file_arr\[17\]\[10\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[10\] rvcpu.dp.rf.reg_file_arr\[19\]\[10\] _08703_
+ _08721_ VGND VGND VPWR VPWR _08824_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_16_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24360_ _09298_ net3528 net61 VGND VGND VPWR VPWR _10358_ sky130_fd_sc_hd__mux2_1
XANTENNA_10 _06600_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_21 _06615_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_191_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_32 _06646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20523_ datamem.data_ram\[22\]\[21\] _07028_ _07182_ datamem.data_ram\[20\]\[21\]
+ VGND VGND VPWR VPWR _07814_ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_43 _06678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_54 _06702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32509_ clknet_leaf_245_clk _03931_ VGND VGND VPWR VPWR datamem.data_ram\[24\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24291_ _09276_ net3789 _10316_ VGND VGND VPWR VPWR _10319_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_65 _06760_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_76 _06776_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26030_ _11081_ _11340_ VGND VGND VPWR VPWR _11342_ sky130_fd_sc_hd__and2_1
XANTENNA_87 _06784_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20454_ _06742_ _07743_ _07745_ VGND VGND VPWR VPWR _07746_ sky130_fd_sc_hd__and3_1
XANTENNA_98 _06837_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_41_Left_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23173_ clknet_1_1__leaf__10108_ VGND VGND VPWR VPWR _10111_ sky130_fd_sc_hd__buf_1
XFILLER_0_28_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20385_ datamem.data_ram\[52\]\[28\] _06685_ _07675_ _07676_ VGND VGND VPWR VPWR
+ _07677_ sky130_fd_sc_hd__o211a_1
XFILLER_0_70_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22124_ _09330_ net2613 _09302_ VGND VGND VPWR VPWR _09331_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_205_5413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27981_ _12178_ _12345_ _12356_ VGND VGND VPWR VPWR _12448_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_219_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_205_5424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29720_ net1066 _01455_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[22\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_26932_ _11829_ _11842_ VGND VGND VPWR VPWR _11846_ sky130_fd_sc_hd__and2_1
X_22055_ rvcpu.dp.plem.WriteDataM\[2\] _09264_ _09265_ rvcpu.dp.plem.WriteDataM\[10\]
+ VGND VGND VPWR VPWR _09275_ sky130_fd_sc_hd__a22o_4
X_21006_ datamem.data_ram\[17\]\[15\] _06653_ _08293_ _08294_ VGND VGND VPWR VPWR
+ _08295_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_197_5214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2930 rvcpu.dp.rf.reg_file_arr\[17\]\[26\] VGND VGND VPWR VPWR net4080 sky130_fd_sc_hd__dlygate4sd3_1
X_29651_ net997 _01386_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[24\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26863_ _11795_ net1608 _11797_ _11801_ VGND VGND VPWR VPWR _03351_ sky130_fd_sc_hd__a31o_1
Xhold2941 datamem.data_ram\[8\]\[12\] VGND VGND VPWR VPWR net4091 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_197_5225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2952 datamem.data_ram\[17\]\[15\] VGND VGND VPWR VPWR net4102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2963 datamem.data_ram\[35\]\[25\] VGND VGND VPWR VPWR net4113 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_214_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28602_ _12687_ net3337 _12796_ VGND VGND VPWR VPWR _12797_ sky130_fd_sc_hd__mux2_1
X_25814_ net1765 _11181_ _11177_ _11202_ VGND VGND VPWR VPWR _02901_ sky130_fd_sc_hd__o211a_1
Xhold2974 rvcpu.dp.rf.reg_file_arr\[29\]\[23\] VGND VGND VPWR VPWR net4124 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2985 rvcpu.dp.rf.reg_file_arr\[13\]\[10\] VGND VGND VPWR VPWR net4135 sky130_fd_sc_hd__dlygate4sd3_1
X_29582_ net936 _01317_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[26\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_214_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26794_ _11753_ net1644 _11748_ _11759_ VGND VGND VPWR VPWR _03324_ sky130_fd_sc_hd__a31o_1
Xhold2996 rvcpu.dp.rf.reg_file_arr\[12\]\[0\] VGND VGND VPWR VPWR net4146 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28533_ _12757_ VGND VGND VPWR VPWR _04065_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_3_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_50_Left_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25745_ _13391_ _11149_ VGND VGND VPWR VPWR _11150_ sky130_fd_sc_hd__nand2_1
Xmax_cap45 _12574_ VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__buf_4
Xmax_cap56 _10839_ VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__buf_4
Xmax_cap67 _12978_ VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__buf_4
X_28464_ _12714_ VGND VGND VPWR VPWR _04039_ sky130_fd_sc_hd__clkbuf_1
X_23346__984 clknet_1_1__leaf__10136_ VGND VGND VPWR VPWR net1110 sky130_fd_sc_hd__inv_2
X_21908_ _08623_ _09134_ _09138_ _09142_ VGND VGND VPWR VPWR _09143_ sky130_fd_sc_hd__and4_1
X_25676_ _11105_ net1557 _11097_ _11107_ VGND VGND VPWR VPWR _02858_ sky130_fd_sc_hd__a31o_1
XFILLER_0_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_156_4232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap89 _10768_ VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__buf_4
X_23503__148 clknet_1_1__leaf__10161_ VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__inv_2
X_22888_ rvcpu.dp.rf.reg_file_arr\[16\]\[31\] rvcpu.dp.rf.reg_file_arr\[17\]\[31\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[31\] rvcpu.dp.rf.reg_file_arr\[19\]\[31\] _09517_
+ _09513_ VGND VGND VPWR VPWR _10023_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_156_4243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1006 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27415_ _12128_ net2722 _12126_ VGND VGND VPWR VPWR _12129_ sky130_fd_sc_hd__mux2_1
XFILLER_0_214_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_194_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24627_ _10516_ VGND VGND VPWR VPWR _02400_ sky130_fd_sc_hd__clkbuf_1
X_28395_ _12439_ net3523 _12669_ VGND VGND VPWR VPWR _12674_ sky130_fd_sc_hd__mux2_1
X_21839_ _08523_ _09076_ VGND VGND VPWR VPWR _09077_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23045__745 clknet_1_0__leaf__10090_ VGND VGND VPWR VPWR net871 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_14_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15360_ _13368_ _13498_ _13894_ rvcpu.dp.pcreg.q\[9\] VGND VGND VPWR VPWR _13895_
+ sky130_fd_sc_hd__o211a_1
X_27346_ _09317_ VGND VGND VPWR VPWR _12089_ sky130_fd_sc_hd__buf_2
XFILLER_0_81_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24558_ _09325_ VGND VGND VPWR VPWR _10478_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_38_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23509_ _09224_ net4373 _10162_ VGND VGND VPWR VPWR _10163_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15291_ _13430_ _13506_ _13447_ _13654_ VGND VGND VPWR VPWR _13829_ sky130_fd_sc_hd__or4_1
XFILLER_0_163_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27277_ _10824_ net2727 _12043_ VGND VGND VPWR VPWR _12050_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24489_ _09318_ datamem.data_ram\[52\]\[28\] _10430_ VGND VGND VPWR VPWR _10435_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29016_ _13018_ net1476 _13009_ _13019_ VGND VGND VPWR VPWR _04286_ sky130_fd_sc_hd__a31o_1
XFILLER_0_145_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17030_ _04769_ VGND VGND VPWR VPWR _01521_ sky130_fd_sc_hd__clkbuf_1
X_26228_ rvcpu.dp.plfd.InstrD\[31\] _11362_ _11452_ VGND VGND VPWR VPWR _11453_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_115_3250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_3261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_180_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26159_ _11416_ VGND VGND VPWR VPWR _03032_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_957 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_186_4951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_186_4962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_111_3169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18981_ _05305_ _05786_ _05776_ _05925_ VGND VGND VPWR VPWR _06317_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_182_4859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17932_ _05304_ VGND VGND VPWR VPWR _05305_ sky130_fd_sc_hd__buf_2
X_29918_ net288 _01653_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[16\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17863_ rvcpu.dp.plde.ALUControlE\[1\] _05236_ VGND VGND VPWR VPWR _05237_ sky130_fd_sc_hd__or2_1
XFILLER_0_139_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29849_ net227 _01584_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[18\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_89_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19602_ datamem.data_ram\[16\]\[8\] _06696_ _06731_ datamem.data_ram\[19\]\[8\] VGND
+ VGND VPWR VPWR _06898_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_145_3980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16814_ _04654_ VGND VGND VPWR VPWR _01630_ sky130_fd_sc_hd__clkbuf_1
X_32860_ clknet_leaf_54_clk _04282_ VGND VGND VPWR VPWR datamem.data_ram\[11\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_17794_ _13268_ _05154_ _05161_ net114 VGND VGND VPWR VPWR _05189_ sky130_fd_sc_hd__a31o_1
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_85_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31811_ clknet_leaf_109_clk _03265_ VGND VGND VPWR VPWR datamem.data_ram\[17\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_19533_ _06828_ VGND VGND VPWR VPWR _06829_ sky130_fd_sc_hd__buf_6
X_16745_ net4192 _14432_ _04612_ VGND VGND VPWR VPWR _04618_ sky130_fd_sc_hd__mux2_1
X_32791_ clknet_leaf_282_clk _04213_ VGND VGND VPWR VPWR datamem.data_ram\[14\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_141_3877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_3888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19464_ _06725_ VGND VGND VPWR VPWR _06760_ sky130_fd_sc_hd__buf_6
X_31742_ net127 _03200_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[9\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_16676_ _04581_ VGND VGND VPWR VPWR _01703_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18415_ _05603_ _05307_ _05437_ _05610_ _05683_ _05579_ VGND VGND VPWR VPWR _05779_
+ sky130_fd_sc_hd__mux4_1
X_15627_ net1910 _13266_ _14114_ VGND VGND VPWR VPWR _14122_ sky130_fd_sc_hd__mux2_1
X_31673_ clknet_leaf_69_clk net1285 VGND VGND VPWR VPWR rvcpu.dp.plmw.ALUResultW\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19395_ _06690_ VGND VGND VPWR VPWR _06691_ sky130_fd_sc_hd__buf_6
XFILLER_0_185_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23478__125 clknet_1_1__leaf__10159_ VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__inv_2
XFILLER_0_130_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18346_ _05274_ _05688_ _05684_ VGND VGND VPWR VPWR _05711_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_44_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30624_ clknet_leaf_188_clk _02359_ VGND VGND VPWR VPWR datamem.data_ram\[52\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_15558_ _13291_ _13414_ _13294_ VGND VGND VPWR VPWR _14082_ sky130_fd_sc_hd__and3_1
XFILLER_0_189_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18277_ rvcpu.dp.plde.RD1E\[29\] _05291_ _05295_ VGND VGND VPWR VPWR _05642_ sky130_fd_sc_hd__o21ai_2
X_30555_ clknet_leaf_177_clk _02290_ VGND VGND VPWR VPWR datamem.data_ram\[55\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_23558__182 clknet_1_1__leaf__10174_ VGND VGND VPWR VPWR net308 sky130_fd_sc_hd__inv_2
X_15489_ _13517_ _13308_ _14004_ _14017_ _13413_ VGND VGND VPWR VPWR _14018_ sky130_fd_sc_hd__o311a_1
XFILLER_0_4_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17228_ _14147_ net2396 _04865_ VGND VGND VPWR VPWR _04874_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30486_ clknet_leaf_207_clk _02221_ VGND VGND VPWR VPWR datamem.data_ram\[57\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32225_ clknet_leaf_169_clk _03647_ VGND VGND VPWR VPWR datamem.data_ram\[35\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold803 rvcpu.dp.rf.reg_file_arr\[2\]\[17\] VGND VGND VPWR VPWR net1953 sky130_fd_sc_hd__dlygate4sd3_1
X_17159_ _04837_ VGND VGND VPWR VPWR _01460_ sky130_fd_sc_hd__clkbuf_1
Xhold814 rvcpu.dp.rf.reg_file_arr\[5\]\[13\] VGND VGND VPWR VPWR net1964 sky130_fd_sc_hd__dlygate4sd3_1
Xhold825 rvcpu.dp.rf.reg_file_arr\[9\]\[28\] VGND VGND VPWR VPWR net1975 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold836 rvcpu.dp.plem.ALUResultM\[7\] VGND VGND VPWR VPWR net1986 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold847 datamem.data_ram\[30\]\[22\] VGND VGND VPWR VPWR net1997 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32156_ clknet_leaf_161_clk _03578_ VGND VGND VPWR VPWR datamem.data_ram\[38\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_20170_ datamem.data_ram\[28\]\[11\] _06688_ _06658_ datamem.data_ram\[25\]\[11\]
+ _07462_ VGND VGND VPWR VPWR _07463_ sky130_fd_sc_hd__o221a_1
Xhold858 rvcpu.dp.rf.reg_file_arr\[19\]\[29\] VGND VGND VPWR VPWR net2008 sky130_fd_sc_hd__dlygate4sd3_1
Xhold869 rvcpu.dp.rf.reg_file_arr\[3\]\[27\] VGND VGND VPWR VPWR net2019 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31107_ clknet_leaf_108_clk _02842_ VGND VGND VPWR VPWR datamem.data_ram\[19\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_24044__573 clknet_1_1__leaf__10245_ VGND VGND VPWR VPWR net699 sky130_fd_sc_hd__inv_2
X_32087_ clknet_leaf_84_clk _03509_ VGND VGND VPWR VPWR datamem.data_ram\[47\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_1141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2204 datamem.data_ram\[50\]\[28\] VGND VGND VPWR VPWR net3354 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2215 datamem.data_ram\[47\]\[20\] VGND VGND VPWR VPWR net3365 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2226 datamem.data_ram\[22\]\[24\] VGND VGND VPWR VPWR net3376 sky130_fd_sc_hd__dlygate4sd3_1
X_31038_ clknet_leaf_60_clk _02773_ VGND VGND VPWR VPWR datamem.data_ram\[41\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2237 rvcpu.dp.rf.reg_file_arr\[22\]\[23\] VGND VGND VPWR VPWR net3387 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1503 datamem.data_ram\[34\]\[26\] VGND VGND VPWR VPWR net2653 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_584 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2248 datamem.data_ram\[39\]\[24\] VGND VGND VPWR VPWR net3398 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1514 rvcpu.dp.rf.reg_file_arr\[23\]\[3\] VGND VGND VPWR VPWR net2664 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2259 datamem.data_ram\[62\]\[10\] VGND VGND VPWR VPWR net3409 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1525 datamem.data_ram\[25\]\[19\] VGND VGND VPWR VPWR net2675 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1536 rvcpu.dp.rf.reg_file_arr\[29\]\[13\] VGND VGND VPWR VPWR net2686 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1547 rvcpu.dp.rf.reg_file_arr\[12\]\[17\] VGND VGND VPWR VPWR net2697 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1558 datamem.data_ram\[39\]\[8\] VGND VGND VPWR VPWR net2708 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1569 datamem.data_ram\[38\]\[9\] VGND VGND VPWR VPWR net2719 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22811_ _09469_ _09950_ VGND VGND VPWR VPWR _09951_ sky130_fd_sc_hd__or2_1
XFILLER_0_224_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_192_5100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_192_5111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32989_ clknet_leaf_205_clk _04411_ VGND VGND VPWR VPWR datamem.data_ram\[62\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25530_ _10727_ net3957 net54 VGND VGND VPWR VPWR _11023_ sky130_fd_sc_hd__mux2_1
XFILLER_0_211_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22742_ _09511_ _09884_ VGND VGND VPWR VPWR _09885_ sky130_fd_sc_hd__or2_1
XFILLER_0_189_491 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_176_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25461_ _10954_ net1515 _10984_ _10986_ VGND VGND VPWR VPWR _02764_ sky130_fd_sc_hd__a31o_1
XFILLER_0_176_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22673_ rvcpu.dp.rf.reg_file_arr\[28\]\[19\] rvcpu.dp.rf.reg_file_arr\[30\]\[19\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[19\] rvcpu.dp.rf.reg_file_arr\[31\]\[19\] _09400_
+ _09484_ VGND VGND VPWR VPWR _09820_ sky130_fd_sc_hd__mux4_1
X_27200_ _11968_ _12008_ VGND VGND VPWR VPWR _12010_ sky130_fd_sc_hd__and2_1
XFILLER_0_168_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24412_ _10113_ _10347_ _10366_ VGND VGND VPWR VPWR _10386_ sky130_fd_sc_hd__a21oi_4
X_28180_ _12557_ VGND VGND VPWR VPWR _03912_ sky130_fd_sc_hd__clkbuf_1
X_21624_ rvcpu.dp.rf.reg_file_arr\[12\]\[12\] rvcpu.dp.rf.reg_file_arr\[13\]\[12\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[12\] rvcpu.dp.rf.reg_file_arr\[15\]\[12\] _08549_
+ _08553_ VGND VGND VPWR VPWR _08874_ sky130_fd_sc_hd__mux4_1
XFILLER_0_47_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25392_ _10946_ _10947_ VGND VGND VPWR VPWR _10950_ sky130_fd_sc_hd__nor2_1
XFILLER_0_192_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27131_ _10209_ _08059_ _11898_ VGND VGND VPWR VPWR _11966_ sky130_fd_sc_hd__and3_1
XFILLER_0_74_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24343_ _09267_ net4293 _10348_ VGND VGND VPWR VPWR _10349_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21555_ _08509_ VGND VGND VPWR VPWR _08808_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27062_ _11922_ VGND VGND VPWR VPWR _11923_ sky130_fd_sc_hd__clkbuf_2
X_20506_ datamem.data_ram\[55\]\[21\] _07021_ _06701_ datamem.data_ram\[49\]\[21\]
+ VGND VGND VPWR VPWR _07797_ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24274_ _09240_ net3732 _10307_ VGND VGND VPWR VPWR _10310_ sky130_fd_sc_hd__mux2_1
X_21486_ rvcpu.dp.plfd.InstrD\[17\] VGND VGND VPWR VPWR _08742_ sky130_fd_sc_hd__buf_2
XFILLER_0_160_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26013_ net20 _11152_ VGND VGND VPWR VPWR _11332_ sky130_fd_sc_hd__or2_1
XFILLER_0_205_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23225_ clknet_1_1__leaf__10108_ VGND VGND VPWR VPWR _10125_ sky130_fd_sc_hd__buf_1
X_20437_ datamem.data_ram\[18\]\[12\] _06611_ _07725_ _07728_ VGND VGND VPWR VPWR
+ _07729_ sky130_fd_sc_hd__o211a_1
XFILLER_0_30_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__11602_ clknet_0__11602_ VGND VGND VPWR VPWR clknet_1_1__leaf__11602_
+ sky130_fd_sc_hd__clkbuf_16
X_20368_ datamem.data_ram\[34\]\[28\] _06689_ _06729_ datamem.data_ram\[35\]\[28\]
+ _06676_ VGND VGND VPWR VPWR _07660_ sky130_fd_sc_hd__o221a_1
Xclkload290 clknet_1_0__leaf__10238_ VGND VGND VPWR VPWR clkload290/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_140_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_149_4080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_219_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22107_ rvcpu.dp.plem.WriteDataM\[28\] _09316_ _09214_ VGND VGND VPWR VPWR _09317_
+ sky130_fd_sc_hd__mux2_8
X_27964_ _12436_ VGND VGND VPWR VPWR _03817_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_224_5866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20299_ datamem.data_ram\[2\]\[19\] _06691_ _06737_ datamem.data_ram\[3\]\[19\] _06769_
+ VGND VGND VPWR VPWR _07592_ sky130_fd_sc_hd__o221a_1
XFILLER_0_105_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_224_5877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26915_ _11831_ net1666 _11821_ _11834_ VGND VGND VPWR VPWR _03370_ sky130_fd_sc_hd__a31o_1
X_22038_ _09260_ net4364 _09232_ VGND VGND VPWR VPWR _09261_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29703_ net1049 _01438_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[22\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_8_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27895_ _12391_ net1686 _12393_ _12398_ VGND VGND VPWR VPWR _03786_ sky130_fd_sc_hd__a31o_1
XFILLER_0_175_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2760 datamem.data_ram\[60\]\[10\] VGND VGND VPWR VPWR net3910 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26846_ _11645_ _11786_ VGND VGND VPWR VPWR _11791_ sky130_fd_sc_hd__and2_1
X_14860_ rvcpu.dp.pcreg.q\[8\] VGND VGND VPWR VPWR _13412_ sky130_fd_sc_hd__clkbuf_4
X_29634_ clknet_leaf_139_clk _01369_ VGND VGND VPWR VPWR datamem.data_ram\[5\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2771 datamem.data_ram\[9\]\[10\] VGND VGND VPWR VPWR net3921 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2782 rvcpu.dp.rf.reg_file_arr\[6\]\[10\] VGND VGND VPWR VPWR net3932 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2793 rvcpu.dp.rf.reg_file_arr\[21\]\[28\] VGND VGND VPWR VPWR net3943 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_1226 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29565_ net919 _01300_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[26\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_26777_ _11676_ _11749_ VGND VGND VPWR VPWR _11750_ sky130_fd_sc_hd__and2_1
X_14791_ _13341_ _13343_ VGND VGND VPWR VPWR _13344_ sky130_fd_sc_hd__nand2_2
XFILLER_0_225_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16530_ _14127_ net4296 _04503_ VGND VGND VPWR VPWR _04504_ sky130_fd_sc_hd__mux2_1
X_28516_ _12745_ net2656 _12735_ VGND VGND VPWR VPWR _12746_ sky130_fd_sc_hd__mux2_1
X_25728_ _10820_ net2513 _11133_ VGND VGND VPWR VPWR _11138_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24190__30 clknet_1_0__leaf__10266_ VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__inv_2
X_29496_ net858 _01231_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[28\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_196_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28447_ _12705_ VGND VGND VPWR VPWR _04031_ sky130_fd_sc_hd__clkbuf_1
X_16461_ _04466_ VGND VGND VPWR VPWR _04467_ sky130_fd_sc_hd__clkbuf_4
X_25659_ _11096_ VGND VGND VPWR VPWR _11097_ sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_191_clk clknet_5_28__leaf_clk VGND VGND VPWR VPWR clknet_leaf_191_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_175_4685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18200_ rvcpu.dp.plde.RD1E\[17\] _05564_ _05499_ VGND VGND VPWR VPWR _05565_ sky130_fd_sc_hd__o21ai_2
X_15412_ _13410_ _13942_ _13943_ _13608_ VGND VGND VPWR VPWR _13944_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_175_4696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19180_ rvcpu.dp.plde.luiE VGND VGND VPWR VPWR _06493_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_186_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28378_ _12664_ VGND VGND VPWR VPWR _04003_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16392_ net2193 _14420_ _14561_ VGND VGND VPWR VPWR _14562_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_117_3312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18131_ _05496_ VGND VGND VPWR VPWR _05497_ sky130_fd_sc_hd__clkbuf_2
X_15343_ _13668_ _13489_ _13374_ VGND VGND VPWR VPWR _13879_ sky130_fd_sc_hd__a21oi_1
X_27329_ _10782_ _12078_ _12079_ net1305 VGND VGND VPWR VPWR _03539_ sky130_fd_sc_hd__o22a_1
XFILLER_0_124_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_113_3209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18062_ rvcpu.dp.plde.ImmExtE\[9\] rvcpu.dp.SrcBFW_Mux.y\[9\] _05277_ VGND VGND VPWR
+ VPWR _05430_ sky130_fd_sc_hd__mux2_2
X_30340_ net686 _02075_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[4\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_15274_ _13300_ _13767_ _13488_ _13401_ VGND VGND VPWR VPWR _13813_ sky130_fd_sc_hd__or4_1
XFILLER_0_0_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17013_ _04760_ VGND VGND VPWR VPWR _01529_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_184_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30271_ net625 _02006_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[6\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32010_ clknet_leaf_127_clk _03432_ VGND VGND VPWR VPWR datamem.data_ram\[27\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_186_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18964_ _05775_ _05724_ _05906_ _06299_ _06300_ VGND VGND VPWR VPWR _06301_ sky130_fd_sc_hd__a311o_1
X_22956__665 clknet_1_0__leaf__10081_ VGND VGND VPWR VPWR net791 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_37_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17915_ _05286_ _05287_ VGND VGND VPWR VPWR _05288_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_37_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_143_3917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18895_ _06004_ _06232_ _06233_ _06236_ VGND VGND VPWR VPWR _06237_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_143_3928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32912_ clknet_leaf_278_clk _04334_ VGND VGND VPWR VPWR datamem.data_ram\[7\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17846_ _13237_ _05179_ _05180_ net114 VGND VGND VPWR VPWR _05225_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_33_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32843_ clknet_leaf_96_clk _04265_ VGND VGND VPWR VPWR datamem.data_ram\[7\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14989_ _13528_ _13536_ _13503_ VGND VGND VPWR VPWR _13537_ sky130_fd_sc_hd__o21a_1
X_17777_ _05174_ VGND VGND VPWR VPWR _05175_ sky130_fd_sc_hd__clkbuf_4
X_23900__459 clknet_1_1__leaf__10223_ VGND VGND VPWR VPWR net585 sky130_fd_sc_hd__inv_2
XFILLER_0_135_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19516_ _06729_ VGND VGND VPWR VPWR _06812_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_89_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16728_ _04608_ VGND VGND VPWR VPWR _01678_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_18_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32774_ clknet_leaf_237_clk _04196_ VGND VGND VPWR VPWR datamem.data_ram\[14\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_102_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_187_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16659_ _14191_ net3132 _04562_ VGND VGND VPWR VPWR _04572_ sky130_fd_sc_hd__mux2_1
X_31725_ net174 _03183_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[9\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_19447_ _06624_ VGND VGND VPWR VPWR _06743_ sky130_fd_sc_hd__clkbuf_8
Xclkbuf_leaf_182_clk clknet_5_22__leaf_clk VGND VGND VPWR VPWR clknet_leaf_182_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_14_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31656_ clknet_leaf_62_clk net4303 VGND VGND VPWR VPWR rvcpu.dp.plmw.ALUResultW\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_19378_ datamem.data_ram\[8\]\[16\] _06649_ _06659_ datamem.data_ram\[9\]\[16\] _06673_
+ VGND VGND VPWR VPWR _06674_ sky130_fd_sc_hd__o221a_1
XFILLER_0_57_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_174_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_846 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18329_ _05693_ VGND VGND VPWR VPWR _05694_ sky130_fd_sc_hd__buf_2
X_30607_ clknet_leaf_196_clk _02342_ VGND VGND VPWR VPWR datamem.data_ram\[52\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_23714__307 clknet_1_1__leaf__10197_ VGND VGND VPWR VPWR net433 sky130_fd_sc_hd__inv_2
X_31587_ clknet_leaf_52_clk net1236 VGND VGND VPWR VPWR rvcpu.dp.plmw.PCPlus4W\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21340_ rvcpu.ALUResultE\[8\] rvcpu.ALUResultE\[9\] _08601_ VGND VGND VPWR VPWR _08602_
+ sky130_fd_sc_hd__or3_1
X_30538_ clknet_leaf_217_clk _02273_ VGND VGND VPWR VPWR datamem.data_ram\[55\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23429__81 clknet_1_1__leaf__10154_ VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__inv_2
XFILLER_0_25_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21271_ rvcpu.dp.plfd.InstrD\[16\] VGND VGND VPWR VPWR _08533_ sky130_fd_sc_hd__clkbuf_8
Xhold600 datamem.data_ram\[7\]\[3\] VGND VGND VPWR VPWR net1750 sky130_fd_sc_hd__dlygate4sd3_1
X_30469_ net147 _02204_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[19\]\[16\] sky130_fd_sc_hd__dfxtp_1
Xhold611 rvcpu.dp.plfd.PCPlus4D\[20\] VGND VGND VPWR VPWR net1761 sky130_fd_sc_hd__dlygate4sd3_1
Xhold622 datamem.data_ram\[51\]\[6\] VGND VGND VPWR VPWR net1772 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20222_ datamem.data_ram\[18\]\[3\] _06931_ _06926_ datamem.data_ram\[23\]\[3\] _06742_
+ VGND VGND VPWR VPWR _07515_ sky130_fd_sc_hd__a221o_1
Xhold633 rvcpu.dp.plfd.PCD\[14\] VGND VGND VPWR VPWR net1783 sky130_fd_sc_hd__dlygate4sd3_1
X_23010_ clknet_1_1__leaf__10080_ VGND VGND VPWR VPWR _10086_ sky130_fd_sc_hd__buf_1
XFILLER_0_229_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold644 datamem.data_ram\[17\]\[1\] VGND VGND VPWR VPWR net1794 sky130_fd_sc_hd__dlygate4sd3_1
X_32208_ clknet_leaf_162_clk _03630_ VGND VGND VPWR VPWR datamem.data_ram\[36\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold655 datamem.data_ram\[34\]\[2\] VGND VGND VPWR VPWR net1805 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold666 datamem.data_ram\[26\]\[3\] VGND VGND VPWR VPWR net1816 sky130_fd_sc_hd__dlygate4sd3_1
Xhold677 datamem.data_ram\[36\]\[7\] VGND VGND VPWR VPWR net1827 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold688 rvcpu.dp.plfd.PCD\[12\] VGND VGND VPWR VPWR net1838 sky130_fd_sc_hd__dlygate4sd3_1
X_32139_ clknet_leaf_241_clk _03561_ VGND VGND VPWR VPWR datamem.data_ram\[39\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_20153_ datamem.data_ram\[49\]\[27\] _06781_ _07444_ _07445_ VGND VGND VPWR VPWR
+ _07446_ sky130_fd_sc_hd__o211a_1
XFILLER_0_100_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold699 rvcpu.dp.plfd.PCPlus4D\[29\] VGND VGND VPWR VPWR net1849 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2001 datamem.data_ram\[49\]\[20\] VGND VGND VPWR VPWR net3151 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2012 rvcpu.dp.rf.reg_file_arr\[13\]\[26\] VGND VGND VPWR VPWR net3162 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2023 datamem.data_ram\[15\]\[29\] VGND VGND VPWR VPWR net3173 sky130_fd_sc_hd__dlygate4sd3_1
X_20084_ _06602_ _07370_ _07372_ _07377_ VGND VGND VPWR VPWR _07378_ sky130_fd_sc_hd__a31o_1
X_24961_ _10392_ net2929 _10696_ VGND VGND VPWR VPWR _10700_ sky130_fd_sc_hd__mux2_1
XFILLER_0_228_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2034 datamem.data_ram\[44\]\[8\] VGND VGND VPWR VPWR net3184 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1300 rvcpu.dp.rf.reg_file_arr\[10\]\[27\] VGND VGND VPWR VPWR net2450 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2045 rvcpu.dp.rf.reg_file_arr\[29\]\[4\] VGND VGND VPWR VPWR net3195 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1311 datamem.data_ram\[47\]\[27\] VGND VGND VPWR VPWR net2461 sky130_fd_sc_hd__dlygate4sd3_1
X_26700_ _10811_ net3126 _11704_ VGND VGND VPWR VPWR _11705_ sky130_fd_sc_hd__mux2_1
Xhold2056 datamem.data_ram\[16\]\[25\] VGND VGND VPWR VPWR net3206 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1322 rvcpu.dp.rf.reg_file_arr\[20\]\[15\] VGND VGND VPWR VPWR net2472 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2067 rvcpu.dp.rf.reg_file_arr\[16\]\[21\] VGND VGND VPWR VPWR net3217 sky130_fd_sc_hd__dlygate4sd3_1
X_27680_ _12093_ net3328 _12270_ VGND VGND VPWR VPWR _12277_ sky130_fd_sc_hd__mux2_1
X_24892_ _10446_ net4054 _10659_ VGND VGND VPWR VPWR _10663_ sky130_fd_sc_hd__mux2_1
X_23760__349 clknet_1_1__leaf__10201_ VGND VGND VPWR VPWR net475 sky130_fd_sc_hd__inv_2
Xhold1333 rvcpu.dp.rf.reg_file_arr\[9\]\[29\] VGND VGND VPWR VPWR net2483 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2078 datamem.data_ram\[2\]\[30\] VGND VGND VPWR VPWR net3228 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1344 rvcpu.dp.rf.reg_file_arr\[14\]\[9\] VGND VGND VPWR VPWR net2494 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2089 datamem.data_ram\[6\]\[29\] VGND VGND VPWR VPWR net3239 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1355 datamem.data_ram\[6\]\[15\] VGND VGND VPWR VPWR net2505 sky130_fd_sc_hd__dlygate4sd3_1
X_26631_ _10783_ _11659_ _11660_ net1339 VGND VGND VPWR VPWR _03260_ sky130_fd_sc_hd__a22o_1
Xclkbuf_1_1__f__10200_ clknet_0__10200_ VGND VGND VPWR VPWR clknet_1_1__leaf__10200_
+ sky130_fd_sc_hd__clkbuf_16
Xhold1366 rvcpu.dp.rf.reg_file_arr\[28\]\[17\] VGND VGND VPWR VPWR net2516 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1377 rvcpu.dp.rf.reg_file_arr\[12\]\[10\] VGND VGND VPWR VPWR net2527 sky130_fd_sc_hd__dlygate4sd3_1
X_23843_ _09330_ net3758 _10210_ VGND VGND VPWR VPWR _10218_ sky130_fd_sc_hd__mux2_1
Xhold1388 datamem.data_ram\[38\]\[18\] VGND VGND VPWR VPWR net2538 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_506 _13209_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1399 rvcpu.dp.rf.reg_file_arr\[20\]\[31\] VGND VGND VPWR VPWR net2549 sky130_fd_sc_hd__dlygate4sd3_1
X_29350_ clknet_leaf_144_clk _01085_ VGND VGND VPWR VPWR datamem.data_ram\[61\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__10131_ clknet_0__10131_ VGND VGND VPWR VPWR clknet_1_1__leaf__10131_
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_517 _13223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_528 _13372_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_212_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26562_ _10822_ net3106 _11620_ VGND VGND VPWR VPWR _11626_ sky130_fd_sc_hd__mux2_1
XFILLER_0_192_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23875__436 clknet_1_0__leaf__10221_ VGND VGND VPWR VPWR net562 sky130_fd_sc_hd__inv_2
XANTENNA_539 _06600_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20986_ datamem.data_ram\[8\]\[15\] _06643_ _08272_ _06614_ _08274_ VGND VGND VPWR
+ VPWR _08275_ sky130_fd_sc_hd__o221a_1
X_28301_ _12447_ net3875 net72 VGND VGND VPWR VPWR _12624_ sky130_fd_sc_hd__mux2_1
X_25513_ _10410_ _11010_ VGND VGND VPWR VPWR _11013_ sky130_fd_sc_hd__and2_1
XFILLER_0_215_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22725_ _09516_ _09868_ VGND VGND VPWR VPWR _09869_ sky130_fd_sc_hd__or2_1
X_29281_ _09309_ net3348 _13159_ VGND VGND VPWR VPWR _13162_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_173_clk clknet_5_24__leaf_clk VGND VGND VPWR VPWR clknet_leaf_173_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_137_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_217_5692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28232_ _12585_ VGND VGND VPWR VPWR _03936_ sky130_fd_sc_hd__clkbuf_1
X_25444_ _10978_ VGND VGND VPWR VPWR _02755_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22656_ _09399_ _09803_ _09523_ VGND VGND VPWR VPWR _09804_ sky130_fd_sc_hd__o21a_1
XFILLER_0_165_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_192_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28163_ _12548_ VGND VGND VPWR VPWR _03904_ sky130_fd_sc_hd__clkbuf_1
X_21607_ _08813_ _08857_ _08689_ VGND VGND VPWR VPWR _08858_ sky130_fd_sc_hd__a21o_1
X_25375_ _10938_ net1527 _10934_ _10939_ VGND VGND VPWR VPWR _02725_ sky130_fd_sc_hd__a31o_1
XFILLER_0_192_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22587_ rvcpu.dp.rf.reg_file_arr\[4\]\[14\] rvcpu.dp.rf.reg_file_arr\[5\]\[14\] rvcpu.dp.rf.reg_file_arr\[6\]\[14\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[14\] _09464_ _09479_ VGND VGND VPWR VPWR _09739_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_170_4571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23654__254 clknet_1_1__leaf__10181_ VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__inv_2
XFILLER_0_8_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27114_ _11938_ net1784 _11952_ _11955_ VGND VGND VPWR VPWR _03448_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_170_4582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24326_ _10339_ VGND VGND VPWR VPWR _02276_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_211_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21538_ rvcpu.dp.rf.reg_file_arr\[8\]\[8\] rvcpu.dp.rf.reg_file_arr\[10\]\[8\] rvcpu.dp.rf.reg_file_arr\[9\]\[8\]
+ rvcpu.dp.rf.reg_file_arr\[11\]\[8\] _08649_ _08537_ VGND VGND VPWR VPWR _08792_
+ sky130_fd_sc_hd__mux4_1
X_28094_ _12450_ net3003 net75 VGND VGND VPWR VPWR _12512_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27045_ _11825_ _11911_ VGND VGND VPWR VPWR _11913_ sky130_fd_sc_hd__and2_1
X_24257_ _09310_ net3865 _10298_ VGND VGND VPWR VPWR _10301_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21469_ rvcpu.dp.rf.reg_file_arr\[28\]\[5\] rvcpu.dp.rf.reg_file_arr\[30\]\[5\] rvcpu.dp.rf.reg_file_arr\[29\]\[5\]
+ rvcpu.dp.rf.reg_file_arr\[31\]\[5\] _08635_ _08637_ VGND VGND VPWR VPWR _08726_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_226_5917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_226_5928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_147_4017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_147_4028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23139_ clknet_1_1__leaf__10087_ VGND VGND VPWR VPWR _10107_ sky130_fd_sc_hd__buf_1
XFILLER_0_222_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28996_ _13007_ VGND VGND VPWR VPWR _04278_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_179_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15961_ _14317_ VGND VGND VPWR VPWR _02046_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_179_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27947_ _12365_ net3393 _12421_ VGND VGND VPWR VPWR _12426_ sky130_fd_sc_hd__mux2_1
Xhold3280 rvcpu.dp.rf.reg_file_arr\[24\]\[23\] VGND VGND VPWR VPWR net4430 sky130_fd_sc_hd__dlygate4sd3_1
X_14912_ _13335_ _13434_ VGND VGND VPWR VPWR _13462_ sky130_fd_sc_hd__nor2_1
Xhold3291 datamem.data_ram\[52\]\[22\] VGND VGND VPWR VPWR net4441 sky130_fd_sc_hd__dlygate4sd3_1
X_17700_ _05124_ VGND VGND VPWR VPWR _01190_ sky130_fd_sc_hd__clkbuf_1
X_18680_ _06028_ _06032_ _06034_ VGND VGND VPWR VPWR _06035_ sky130_fd_sc_hd__or3b_1
X_27878_ _12153_ net3100 net77 VGND VGND VPWR VPWR _12388_ sky130_fd_sc_hd__mux2_1
X_15892_ net3520 _13198_ _14275_ VGND VGND VPWR VPWR _14281_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_106_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2590 datamem.data_ram\[35\]\[16\] VGND VGND VPWR VPWR net3740 sky130_fd_sc_hd__dlygate4sd3_1
X_14843_ _13370_ _13372_ _13374_ _13386_ _13395_ VGND VGND VPWR VPWR _13396_ sky130_fd_sc_hd__o311a_1
X_17631_ net2118 _13197_ _05082_ VGND VGND VPWR VPWR _05088_ sky130_fd_sc_hd__mux2_1
X_29617_ net971 _01352_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[25\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_26829_ _11767_ net1553 _11773_ _11780_ VGND VGND VPWR VPWR _03338_ sky130_fd_sc_hd__a31o_1
XFILLER_0_216_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_177_4736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_177_4747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17562_ _05051_ VGND VGND VPWR VPWR _01255_ sky130_fd_sc_hd__clkbuf_1
X_14774_ _13326_ VGND VGND VPWR VPWR _13327_ sky130_fd_sc_hd__clkbuf_4
X_29548_ net902 _01283_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[27\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19301_ _06585_ rvcpu.dp.plem.ALUResultM\[5\] VGND VGND VPWR VPWR _06597_ sky130_fd_sc_hd__and2_1
X_16513_ _04494_ VGND VGND VPWR VPWR _01787_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17493_ _13195_ net4063 _05010_ VGND VGND VPWR VPWR _05015_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_164_clk clknet_5_25__leaf_clk VGND VGND VPWR VPWR clknet_leaf_164_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_6_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29479_ net841 _01214_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[2\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_31510_ clknet_leaf_65_clk net1204 VGND VGND VPWR VPWR rvcpu.dp.plem.PCPlus4M\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_19232_ _06534_ _06537_ VGND VGND VPWR VPWR _06538_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_155_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16444_ net1983 _14474_ _04451_ VGND VGND VPWR VPWR _04457_ sky130_fd_sc_hd__mux2_1
X_32490_ clknet_leaf_81_clk _03912_ VGND VGND VPWR VPWR datamem.data_ram\[25\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19163_ _06476_ _06477_ VGND VGND VPWR VPWR _06478_ sky130_fd_sc_hd__and2_1
X_31441_ clknet_leaf_67_clk net1179 VGND VGND VPWR VPWR rvcpu.dp.plem.ResultSrcM\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_136_3754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16375_ _14552_ VGND VGND VPWR VPWR _01851_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_3765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18114_ _05479_ _05480_ VGND VGND VPWR VPWR _05481_ sky130_fd_sc_hd__nor2_2
X_15326_ _13798_ _13862_ _13442_ VGND VGND VPWR VPWR _13863_ sky130_fd_sc_hd__a21o_1
XFILLER_0_82_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19094_ _06407_ _06416_ VGND VGND VPWR VPWR _06417_ sky130_fd_sc_hd__or2_1
X_31372_ clknet_leaf_18_clk _03075_ VGND VGND VPWR VPWR rvcpu.dp.plde.ImmExtE\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__10220_ clknet_0__10220_ VGND VGND VPWR VPWR clknet_1_0__leaf__10220_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_53_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18045_ _05414_ VGND VGND VPWR VPWR rvcpu.dp.SrcBFW_Mux.y\[10\] sky130_fd_sc_hd__buf_1
X_30323_ net669 _02058_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[4\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15257_ _13369_ _13796_ VGND VGND VPWR VPWR _13797_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_227_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30254_ net608 _01989_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[6\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_15188_ _13465_ _13639_ _13640_ _13463_ VGND VGND VPWR VPWR _13731_ sky130_fd_sc_hd__o31a_1
XFILLER_0_10_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__10082_ clknet_0__10082_ VGND VGND VPWR VPWR clknet_1_0__leaf__10082_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_201_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30185_ net539 _01920_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[8\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_19996_ datamem.data_ram\[21\]\[2\] _06919_ _06953_ datamem.data_ram\[20\]\[2\] _07289_
+ VGND VGND VPWR VPWR _07290_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_35_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18947_ _06109_ _05863_ VGND VGND VPWR VPWR _06285_ sky130_fd_sc_hd__or2_1
XFILLER_0_225_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_193_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18878_ _05473_ _05728_ _06197_ _06220_ VGND VGND VPWR VPWR _06221_ sky130_fd_sc_hd__a211o_1
XFILLER_0_146_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17829_ rvcpu.dp.plem.ALUResultM\[23\] _05213_ _05177_ VGND VGND VPWR VPWR _05214_
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_6_Left_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_178_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32826_ clknet_leaf_156_clk _04248_ VGND VGND VPWR VPWR datamem.data_ram\[12\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_20840_ datamem.data_ram\[24\]\[14\] _06649_ _06701_ datamem.data_ram\[25\]\[14\]
+ _08129_ VGND VGND VPWR VPWR _08130_ sky130_fd_sc_hd__o221a_1
XFILLER_0_222_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20771_ _07635_ datamem.data_ram\[63\]\[6\] VGND VGND VPWR VPWR _08061_ sky130_fd_sc_hd__and2_1
XFILLER_0_162_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_155_clk clknet_5_28__leaf_clk VGND VGND VPWR VPWR clknet_leaf_155_clk
+ sky130_fd_sc_hd__clkbuf_8
X_32757_ clknet_leaf_164_clk _04179_ VGND VGND VPWR VPWR datamem.data_ram\[15\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22510_ _09461_ _09663_ _09665_ _09489_ VGND VGND VPWR VPWR _09666_ sky130_fd_sc_hd__o211a_1
X_31708_ clknet_leaf_31_clk _03166_ VGND VGND VPWR VPWR rvcpu.dp.pcreg.q\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32688_ clknet_leaf_172_clk _04110_ VGND VGND VPWR VPWR datamem.data_ram\[18\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_1331 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22441_ rvcpu.dp.rf.reg_file_arr\[20\]\[7\] rvcpu.dp.rf.reg_file_arr\[21\]\[7\] rvcpu.dp.rf.reg_file_arr\[22\]\[7\]
+ rvcpu.dp.rf.reg_file_arr\[23\]\[7\] _09512_ _09408_ VGND VGND VPWR VPWR _09600_
+ sky130_fd_sc_hd__mux4_1
X_31639_ clknet_leaf_68_clk net1152 VGND VGND VPWR VPWR rvcpu.dp.plmw.lAuiPCW\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25160_ _10813_ VGND VGND VPWR VPWR _02636_ sky130_fd_sc_hd__clkbuf_1
X_22372_ rvcpu.dp.rf.reg_file_arr\[12\]\[3\] rvcpu.dp.rf.reg_file_arr\[13\]\[3\] rvcpu.dp.rf.reg_file_arr\[14\]\[3\]
+ rvcpu.dp.rf.reg_file_arr\[15\]\[3\] _09434_ _09382_ VGND VGND VPWR VPWR _09535_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_115_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21323_ rvcpu.dp.plfd.InstrD\[17\] rvcpu.dp.plde.RdE\[2\] VGND VGND VPWR VPWR _08585_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25091_ _07136_ VGND VGND VPWR VPWR _10777_ sky130_fd_sc_hd__buf_8
XFILLER_0_142_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21254_ rvcpu.dp.plfd.InstrD\[15\] VGND VGND VPWR VPWR _08516_ sky130_fd_sc_hd__buf_6
Xhold430 datamem.data_ram\[18\]\[1\] VGND VGND VPWR VPWR net1580 sky130_fd_sc_hd__dlygate4sd3_1
Xhold441 datamem.data_ram\[1\]\[3\] VGND VGND VPWR VPWR net1591 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold452 datamem.data_ram\[24\]\[4\] VGND VGND VPWR VPWR net1602 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold463 datamem.data_ram\[63\]\[6\] VGND VGND VPWR VPWR net1613 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20205_ datamem.data_ram\[50\]\[11\] _06691_ _06760_ datamem.data_ram\[55\]\[11\]
+ VGND VGND VPWR VPWR _07498_ sky130_fd_sc_hd__o22a_1
Xhold474 datamem.data_ram\[57\]\[1\] VGND VGND VPWR VPWR net1624 sky130_fd_sc_hd__dlygate4sd3_1
X_21185_ _06910_ _06580_ _08468_ _06909_ VGND VGND VPWR VPWR _08472_ sky130_fd_sc_hd__o22ai_1
X_28850_ _12928_ VGND VGND VPWR VPWR _04211_ sky130_fd_sc_hd__clkbuf_1
Xhold485 datamem.data_ram\[57\]\[0\] VGND VGND VPWR VPWR net1635 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_221_5803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold496 datamem.data_ram\[37\]\[2\] VGND VGND VPWR VPWR net1646 sky130_fd_sc_hd__dlygate4sd3_1
X_27801_ _12342_ VGND VGND VPWR VPWR _03748_ sky130_fd_sc_hd__clkbuf_1
X_20136_ datamem.data_ram\[35\]\[27\] _06632_ _06704_ datamem.data_ram\[39\]\[27\]
+ _06677_ VGND VGND VPWR VPWR _07429_ sky130_fd_sc_hd__o221a_1
X_28781_ _12760_ net4189 _12887_ VGND VGND VPWR VPWR _12892_ sky130_fd_sc_hd__mux2_1
X_25993_ net10 _11317_ VGND VGND VPWR VPWR _11321_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27732_ _12093_ net3931 _12298_ VGND VGND VPWR VPWR _12305_ sky130_fd_sc_hd__mux2_1
X_24944_ _10446_ net3546 _10687_ VGND VGND VPWR VPWR _10691_ sky130_fd_sc_hd__mux2_1
X_20067_ datamem.data_ram\[48\]\[26\] _06645_ _06617_ datamem.data_ram\[52\]\[26\]
+ _07360_ VGND VGND VPWR VPWR _07361_ sky130_fd_sc_hd__o221a_1
Xhold1130 rvcpu.dp.rf.reg_file_arr\[24\]\[7\] VGND VGND VPWR VPWR net2280 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1141 datamem.data_ram\[29\]\[10\] VGND VGND VPWR VPWR net2291 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1152 datamem.data_ram\[29\]\[21\] VGND VGND VPWR VPWR net2302 sky130_fd_sc_hd__dlygate4sd3_1
X_27663_ _12155_ net3854 _12261_ VGND VGND VPWR VPWR _12268_ sky130_fd_sc_hd__mux2_1
X_24875_ _10472_ net3780 net92 VGND VGND VPWR VPWR _10654_ sky130_fd_sc_hd__mux2_1
Xhold1163 rvcpu.dp.rf.reg_file_arr\[11\]\[29\] VGND VGND VPWR VPWR net2313 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_217_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1174 datamem.data_ram\[6\]\[23\] VGND VGND VPWR VPWR net2324 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1185 rvcpu.dp.rf.reg_file_arr\[6\]\[28\] VGND VGND VPWR VPWR net2335 sky130_fd_sc_hd__dlygate4sd3_1
X_29402_ clknet_leaf_0_clk _01137_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD2E\[13\] sky130_fd_sc_hd__dfxtp_1
X_26614_ _10820_ net2503 _11650_ VGND VGND VPWR VPWR _11655_ sky130_fd_sc_hd__mux2_1
Xhold1196 rvcpu.dp.rf.reg_file_arr\[8\]\[22\] VGND VGND VPWR VPWR net2346 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_219_5743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_866 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_303 _14133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_219_5754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27594_ _12138_ net1895 _12224_ VGND VGND VPWR VPWR _12231_ sky130_fd_sc_hd__mux2_1
XANTENNA_314 _14177_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_325 _14447_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_213_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_206_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_185_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_336 _14461_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_347 datamem.data_ram\[52\]\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26545_ _11517_ net1603 _11608_ _11616_ VGND VGND VPWR VPWR _03218_ sky130_fd_sc_hd__a31o_1
X_29333_ clknet_leaf_267_clk _01068_ VGND VGND VPWR VPWR datamem.data_ram\[62\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_358 rvcpu.dp.SrcBFW_Mux.y\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_146_clk clknet_5_29__leaf_clk VGND VGND VPWR VPWR clknet_leaf_146_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_369 rvcpu.dp.plde.ImmExtE\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20969_ datamem.data_ram\[35\]\[15\] _06639_ VGND VGND VPWR VPWR _08258_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_172_4622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23124__801 clknet_1_0__leaf__10105_ VGND VGND VPWR VPWR net927 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_172_4633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29264_ _09275_ net4357 _13150_ VGND VGND VPWR VPWR _13153_ sky130_fd_sc_hd__mux2_1
X_22708_ rvcpu.dp.rf.reg_file_arr\[28\]\[21\] rvcpu.dp.rf.reg_file_arr\[30\]\[21\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[21\] rvcpu.dp.rf.reg_file_arr\[31\]\[21\] _09443_
+ _09453_ VGND VGND VPWR VPWR _09853_ sky130_fd_sc_hd__mux4_1
X_26476_ _11576_ _11249_ _11522_ _06558_ _11595_ VGND VGND VPWR VPWR _11596_ sky130_fd_sc_hd__a221o_1
XFILLER_0_177_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28215_ _12576_ VGND VGND VPWR VPWR _03928_ sky130_fd_sc_hd__clkbuf_1
X_25427_ _10969_ VGND VGND VPWR VPWR _02747_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_192_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22639_ rvcpu.dp.rf.reg_file_arr\[4\]\[17\] rvcpu.dp.rf.reg_file_arr\[5\]\[17\] rvcpu.dp.rf.reg_file_arr\[6\]\[17\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[17\] _09604_ _09716_ VGND VGND VPWR VPWR _09788_
+ sky130_fd_sc_hd__mux4_1
X_29195_ _13115_ VGND VGND VPWR VPWR _04369_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_192_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16160_ net3440 _14424_ _14422_ VGND VGND VPWR VPWR _14425_ sky130_fd_sc_hd__mux2_1
X_28146_ _12539_ VGND VGND VPWR VPWR _03896_ sky130_fd_sc_hd__clkbuf_1
X_25358_ _10067_ _10923_ VGND VGND VPWR VPWR _10928_ sky130_fd_sc_hd__and2_1
XFILLER_0_35_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload19 clknet_5_23__leaf_clk VGND VGND VPWR VPWR clkload19/Y sky130_fd_sc_hd__clkinvlp_4
X_15111_ _13303_ _13432_ VGND VGND VPWR VPWR _13656_ sky130_fd_sc_hd__nor2_1
XFILLER_0_140_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24309_ _09306_ net3813 _10328_ VGND VGND VPWR VPWR _10330_ sky130_fd_sc_hd__mux2_1
X_28077_ _12433_ net3601 _12501_ VGND VGND VPWR VPWR _12503_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_131_3640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16091_ _14387_ VGND VGND VPWR VPWR _01978_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_131_3651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25289_ _10741_ _10114_ _10828_ VGND VGND VPWR VPWR _10887_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_20_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15042_ _13387_ _13402_ VGND VGND VPWR VPWR _13589_ sky130_fd_sc_hd__nor2_2
X_27028_ _11889_ net1510 _11897_ _11902_ VGND VGND VPWR VPWR _03415_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_71_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_181_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19850_ datamem.data_ram\[51\]\[1\] _06966_ _06927_ datamem.data_ram\[55\]\[1\] _07144_
+ VGND VGND VPWR VPWR _07145_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18801_ _06136_ _05765_ _06140_ _06148_ VGND VGND VPWR VPWR _06149_ sky130_fd_sc_hd__o211ai_1
X_19781_ datamem.data_ram\[32\]\[9\] _06649_ _07072_ _07075_ VGND VGND VPWR VPWR _07076_
+ sky130_fd_sc_hd__o211a_1
X_28979_ _12995_ net1369 _12988_ _12998_ VGND VGND VPWR VPWR _04270_ sky130_fd_sc_hd__a31o_1
X_16993_ net2786 _14476_ _04742_ VGND VGND VPWR VPWR _04749_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_129_3580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18732_ _06077_ _06080_ _06083_ _05239_ VGND VGND VPWR VPWR _06084_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_129_3591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15944_ net2807 _13275_ _14274_ VGND VGND VPWR VPWR _14308_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31990_ clknet_leaf_117_clk _03412_ VGND VGND VPWR VPWR datamem.data_ram\[37\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_30_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23211__862 clknet_1_1__leaf__10112_ VGND VGND VPWR VPWR net988 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_30_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30941_ clknet_leaf_95_clk _02676_ VGND VGND VPWR VPWR datamem.data_ram\[3\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18663_ _05442_ _05444_ VGND VGND VPWR VPWR _06018_ sky130_fd_sc_hd__or2_1
X_15875_ net2087 _13278_ _14235_ VGND VGND VPWR VPWR _14270_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_125_3488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_3499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14826_ _13296_ _13378_ VGND VGND VPWR VPWR _13379_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17614_ _05078_ VGND VGND VPWR VPWR _01230_ sky130_fd_sc_hd__clkbuf_1
X_30872_ clknet_leaf_57_clk _02607_ VGND VGND VPWR VPWR datamem.data_ram\[42\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_18594_ _05933_ _05934_ _05952_ VGND VGND VPWR VPWR _05953_ sky130_fd_sc_hd__o21a_1
XFILLER_0_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32611_ clknet_leaf_78_clk _04033_ VGND VGND VPWR VPWR datamem.data_ram\[20\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_14757_ _13292_ _13294_ _13302_ _13309_ VGND VGND VPWR VPWR _13310_ sky130_fd_sc_hd__or4_1
X_17545_ _13272_ net2541 _05032_ VGND VGND VPWR VPWR _05042_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_137_clk clknet_5_30__leaf_clk VGND VGND VPWR VPWR clknet_leaf_137_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_138_3805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32542_ clknet_leaf_83_clk _03964_ VGND VGND VPWR VPWR datamem.data_ram\[23\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_17476_ _05005_ VGND VGND VPWR VPWR _01303_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14688_ _13250_ VGND VGND VPWR VPWR _13251_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_28_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19215_ rvcpu.dp.plde.ImmExtE\[25\] rvcpu.dp.plde.PCE\[25\] VGND VGND VPWR VPWR _06523_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16427_ net3728 _14457_ _14572_ VGND VGND VPWR VPWR _14580_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32473_ clknet_leaf_247_clk _03895_ VGND VGND VPWR VPWR datamem.data_ram\[26\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_60_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19146_ _06462_ VGND VGND VPWR VPWR rvcpu.dp.lAuiPCE\[16\] sky130_fd_sc_hd__clkbuf_1
X_31424_ clknet_leaf_60_clk _03127_ VGND VGND VPWR VPWR datamem.data_ram\[44\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_16358_ _14543_ VGND VGND VPWR VPWR _01859_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15309_ _13822_ _13828_ _13846_ VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__o21a_1
XFILLER_0_143_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31355_ clknet_leaf_17_clk _03058_ VGND VGND VPWR VPWR rvcpu.dp.plde.ImmExtE\[4\]
+ sky130_fd_sc_hd__dfxtp_4
X_19077_ _06400_ _06401_ VGND VGND VPWR VPWR _06402_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__10203_ clknet_0__10203_ VGND VGND VPWR VPWR clknet_1_0__leaf__10203_
+ sky130_fd_sc_hd__clkbuf_16
X_16289_ net2943 _14455_ _14500_ VGND VGND VPWR VPWR _14507_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30306_ net652 _02041_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[5\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_18028_ _05321_ rvcpu.dp.SrcBFW_Mux.y\[2\] _05379_ VGND VGND VPWR VPWR _05398_ sky130_fd_sc_hd__o21ai_2
X_31286_ clknet_leaf_108_clk _02989_ VGND VGND VPWR VPWR datamem.data_ram\[34\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__10134_ clknet_0__10134_ VGND VGND VPWR VPWR clknet_1_0__leaf__10134_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_199_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30237_ net591 _01972_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[7\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23826__408 clknet_1_0__leaf__10208_ VGND VGND VPWR VPWR net534 sky130_fd_sc_hd__inv_2
XFILLER_0_199_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_226_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30168_ net530 _01903_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[0\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19979_ datamem.data_ram\[18\]\[18\] _06612_ _07269_ _07272_ VGND VGND VPWR VPWR
+ _07273_ sky130_fd_sc_hd__o211a_1
XFILLER_0_226_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30099_ net461 _01834_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[11\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_21941_ rvcpu.dp.rf.reg_file_arr\[12\]\[29\] rvcpu.dp.rf.reg_file_arr\[13\]\[29\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[29\] rvcpu.dp.rf.reg_file_arr\[15\]\[29\] _08839_
+ _08840_ VGND VGND VPWR VPWR _09174_ sky130_fd_sc_hd__mux4_1
XFILLER_0_179_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24660_ _10412_ net1484 _10531_ _10535_ VGND VGND VPWR VPWR _02414_ sky130_fd_sc_hd__a31o_1
XFILLER_0_179_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21872_ _09100_ _09104_ _09108_ _08624_ VGND VGND VPWR VPWR _01053_ sky130_fd_sc_hd__o31a_1
XFILLER_0_167_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32809_ clknet_leaf_255_clk _04231_ VGND VGND VPWR VPWR datamem.data_ram\[13\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20823_ datamem.data_ram\[26\]\[30\] _06940_ _06934_ datamem.data_ram\[24\]\[30\]
+ VGND VGND VPWR VPWR _08113_ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_128_clk clknet_5_31__leaf_clk VGND VGND VPWR VPWR clknet_leaf_128_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_194_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24591_ _10496_ VGND VGND VPWR VPWR _02384_ sky130_fd_sc_hd__clkbuf_1
X_26330_ _11083_ _11497_ VGND VGND VPWR VPWR _11500_ sky130_fd_sc_hd__and2_1
XFILLER_0_119_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20754_ _07635_ datamem.data_ram\[10\]\[6\] datamem.data_ram\[11\]\[6\] _07833_ _07636_
+ VGND VGND VPWR VPWR _08044_ sky130_fd_sc_hd__o221a_1
XFILLER_0_33_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_214_5640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26261_ _11462_ VGND VGND VPWR VPWR _03088_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_210_5526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20685_ datamem.data_ram\[53\]\[5\] _06970_ _07137_ datamem.data_ram\[51\]\[5\] _06603_
+ VGND VGND VPWR VPWR _07976_ sky130_fd_sc_hd__a221o_1
X_28000_ _12460_ net3259 net76 VGND VGND VPWR VPWR _12461_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_210_5537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25212_ _10822_ net3978 net56 VGND VGND VPWR VPWR _10845_ sky130_fd_sc_hd__mux2_1
XFILLER_0_190_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22424_ _09510_ _09576_ _09579_ _09583_ _09525_ VGND VGND VPWR VPWR _09584_ sky130_fd_sc_hd__a311o_2
XFILLER_0_208_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26192_ _11433_ VGND VGND VPWR VPWR _03048_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25143_ _10754_ net2611 _10802_ VGND VGND VPWR VPWR _10804_ sky130_fd_sc_hd__mux2_1
X_22355_ rvcpu.dp.rf.reg_file_arr\[20\]\[3\] rvcpu.dp.rf.reg_file_arr\[21\]\[3\] rvcpu.dp.rf.reg_file_arr\[22\]\[3\]
+ rvcpu.dp.rf.reg_file_arr\[23\]\[3\] _09517_ _09513_ VGND VGND VPWR VPWR _09518_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_60_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21306_ _08552_ VGND VGND VPWR VPWR _08568_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_142_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25074_ _10741_ _10640_ _10705_ VGND VGND VPWR VPWR _10768_ sky130_fd_sc_hd__a21oi_4
X_29951_ net321 _01686_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[15\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22286_ _09398_ VGND VGND VPWR VPWR _09451_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_143_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23154__827 clknet_1_1__leaf__10109_ VGND VGND VPWR VPWR net953 sky130_fd_sc_hd__inv_2
X_28902_ _12745_ net3556 net68 VGND VGND VPWR VPWR _12956_ sky130_fd_sc_hd__mux2_1
Xhold260 datamem.data_ram\[30\]\[5\] VGND VGND VPWR VPWR net1410 sky130_fd_sc_hd__dlygate4sd3_1
X_21237_ datamem.data_ram\[52\]\[4\] datamem.data_ram\[53\]\[4\] datamem.data_ram\[52\]\[28\]
+ datamem.data_ram\[52\]\[20\] VGND VGND VPWR VPWR _08500_ sky130_fd_sc_hd__and4_1
XFILLER_0_104_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_208_5477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold271 datamem.data_ram\[28\]\[7\] VGND VGND VPWR VPWR net1421 sky130_fd_sc_hd__dlygate4sd3_1
X_29882_ net260 _01617_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[17\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_208_5488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold282 datamem.data_ram\[48\]\[1\] VGND VGND VPWR VPWR net1432 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_208_5499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold293 datamem.data_ram\[33\]\[1\] VGND VGND VPWR VPWR net1443 sky130_fd_sc_hd__dlygate4sd3_1
X_28833_ _12919_ VGND VGND VPWR VPWR _04203_ sky130_fd_sc_hd__clkbuf_1
X_21168_ datamem.data_ram\[12\]\[23\] datamem.data_ram\[13\]\[23\] _07824_ VGND VGND
+ VPWR VPWR _08457_ sky130_fd_sc_hd__mux2_1
XFILLER_0_218_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_176_1110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_4356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20119_ _07390_ _07412_ VGND VGND VPWR VPWR _07413_ sky130_fd_sc_hd__nor2_4
XFILLER_0_217_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21099_ datamem.data_ram\[14\]\[7\] datamem.data_ram\[15\]\[7\] _07824_ VGND VGND
+ VPWR VPWR _08388_ sky130_fd_sc_hd__mux2_1
X_25976_ net3 _11289_ VGND VGND VPWR VPWR _11311_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_161_4367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28764_ _12882_ VGND VGND VPWR VPWR _04171_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24927_ _10472_ net3825 net91 VGND VGND VPWR VPWR _10682_ sky130_fd_sc_hd__mux2_1
X_27715_ _12155_ net2084 net50 VGND VGND VPWR VPWR _12296_ sky130_fd_sc_hd__mux2_1
X_28695_ _12743_ net4017 net42 VGND VGND VPWR VPWR _12846_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15660_ _14143_ net4390 _14131_ VGND VGND VPWR VPWR _14144_ sky130_fd_sc_hd__mux2_1
X_27646_ _12258_ VGND VGND VPWR VPWR _03677_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_100 _06862_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24858_ _10392_ net2303 net93 VGND VGND VPWR VPWR _10645_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_111 _07077_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14611_ _13168_ VGND VGND VPWR VPWR _13192_ sky130_fd_sc_hd__clkbuf_8
XANTENNA_122 _07226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_133 _07831_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_212_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_119_clk clknet_5_27__leaf_clk VGND VGND VPWR VPWR clknet_leaf_119_clk
+ sky130_fd_sc_hd__clkbuf_8
X_15591_ _14091_ VGND VGND VPWR VPWR _14103_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_144 _07840_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27577_ _12093_ net2481 _12215_ VGND VGND VPWR VPWR _12222_ sky130_fd_sc_hd__mux2_1
XANTENNA_155 _08353_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24789_ _10474_ net3980 net94 VGND VGND VPWR VPWR _10607_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_120_3385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_166 _08667_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17330_ _04928_ VGND VGND VPWR VPWR _01380_ sky130_fd_sc_hd__clkbuf_1
X_26528_ _11374_ _06567_ _11367_ _11375_ VGND VGND VPWR VPWR _11606_ sky130_fd_sc_hd__a211o_1
X_29316_ clknet_leaf_11_clk _01051_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD1E\[23\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_177 _08937_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_188 _09195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_199 _09476_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0__10128_ _10128_ VGND VGND VPWR VPWR clknet_0__10128_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_3_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17261_ _04891_ VGND VGND VPWR VPWR _01412_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_78_Left_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26459_ net1859 _11573_ _11584_ _11570_ VGND VGND VPWR VPWR _03164_ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29247_ _09239_ net3252 _13141_ VGND VGND VPWR VPWR _13144_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_423 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19000_ _05240_ _06321_ _06322_ _06334_ VGND VGND VPWR VPWR rvcpu.ALUResultE\[29\]
+ sky130_fd_sc_hd__a31o_1
X_16212_ net2189 _14459_ _14443_ VGND VGND VPWR VPWR _14460_ sky130_fd_sc_hd__mux2_1
X_29178_ _13106_ VGND VGND VPWR VPWR _04361_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_23_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17192_ _14179_ net2744 _04851_ VGND VGND VPWR VPWR _04855_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_23_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_180_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload108 clknet_leaf_53_clk VGND VGND VPWR VPWR clkload108/Y sky130_fd_sc_hd__clkinvlp_2
XTAP_TAPCELL_ROW_12_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload119 clknet_leaf_101_clk VGND VGND VPWR VPWR clkload119/Y sky130_fd_sc_hd__clkinv_4
X_28129_ _12530_ VGND VGND VPWR VPWR _03888_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_12_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16143_ _14414_ VGND VGND VPWR VPWR _01953_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31140_ clknet_leaf_187_clk _02875_ VGND VGND VPWR VPWR datamem.data_ram\[4\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16074_ net2665 _13263_ _14371_ VGND VGND VPWR VPWR _14378_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_5_14__f_clk clknet_2_1_0_clk VGND VGND VPWR VPWR clknet_5_14__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_121_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15025_ _13521_ VGND VGND VPWR VPWR _13572_ sky130_fd_sc_hd__clkbuf_4
X_19902_ datamem.data_ram\[10\]\[17\] _06613_ _06665_ datamem.data_ram\[13\]\[17\]
+ VGND VGND VPWR VPWR _07197_ sky130_fd_sc_hd__o22a_1
XFILLER_0_220_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31071_ clknet_leaf_177_clk _02806_ VGND VGND VPWR VPWR datamem.data_ram\[9\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_23094__774 clknet_1_0__leaf__10102_ VGND VGND VPWR VPWR net900 sky130_fd_sc_hd__inv_2
X_30022_ net384 _01757_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[13\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_19833_ datamem.data_ram\[38\]\[1\] _07127_ _06966_ datamem.data_ram\[35\]\[1\] _06967_
+ VGND VGND VPWR VPWR _07128_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_87_Left_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_209_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_194_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_127_3539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19764_ datamem.data_ram\[20\]\[25\] _07024_ _06700_ datamem.data_ram\[17\]\[25\]
+ VGND VGND VPWR VPWR _07059_ sky130_fd_sc_hd__o22a_1
XFILLER_0_223_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16976_ net3017 _14459_ _04731_ VGND VGND VPWR VPWR _04740_ sky130_fd_sc_hd__mux2_1
X_18715_ _06055_ _06056_ _06057_ _06067_ VGND VGND VPWR VPWR _06068_ sky130_fd_sc_hd__a31o_1
XFILLER_0_95_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15927_ _14299_ VGND VGND VPWR VPWR _02062_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_223_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19695_ datamem.data_ram\[12\]\[0\] _06955_ _06958_ datamem.data_ram\[9\]\[0\] VGND
+ VGND VPWR VPWR _06991_ sky130_fd_sc_hd__a22o_1
X_31973_ clknet_leaf_129_clk _03395_ VGND VGND VPWR VPWR datamem.data_ram\[54\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18646_ _05866_ _05754_ _06001_ _05720_ VGND VGND VPWR VPWR _06002_ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30924_ clknet_leaf_200_clk _02659_ VGND VGND VPWR VPWR datamem.data_ram\[40\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_15858_ _14261_ VGND VGND VPWR VPWR _02093_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14809_ _13327_ _13339_ _13355_ _13361_ VGND VGND VPWR VPWR _13362_ sky130_fd_sc_hd__a211o_1
X_18577_ _05823_ _05825_ _05675_ VGND VGND VPWR VPWR _05936_ sky130_fd_sc_hd__mux2_1
X_30855_ clknet_leaf_150_clk _02590_ VGND VGND VPWR VPWR datamem.data_ram\[43\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15789_ _14224_ VGND VGND VPWR VPWR _02133_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17528_ _05033_ VGND VGND VPWR VPWR _01279_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_96_Left_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30786_ clknet_leaf_136_clk _02521_ VGND VGND VPWR VPWR datamem.data_ram\[46\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32525_ clknet_leaf_253_clk _03947_ VGND VGND VPWR VPWR datamem.data_ram\[24\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_17459_ _14172_ net3183 _04996_ VGND VGND VPWR VPWR _04997_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20470_ datamem.data_ram\[40\]\[20\] _06778_ _07761_ _06601_ VGND VGND VPWR VPWR
+ _07762_ sky130_fd_sc_hd__o211a_1
X_32456_ clknet_leaf_276_clk _03878_ VGND VGND VPWR VPWR datamem.data_ram\[27\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_229_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19129_ _06447_ net4424 _06419_ VGND VGND VPWR VPWR _06448_ sky130_fd_sc_hd__mux2_1
X_31407_ clknet_leaf_32_clk _03110_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCE\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_1099 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32387_ clknet_leaf_240_clk _03809_ VGND VGND VPWR VPWR datamem.data_ram\[29\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22140_ _09339_ VGND VGND VPWR VPWR _01090_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31338_ clknet_leaf_17_clk _03041_ VGND VGND VPWR VPWR rvcpu.dp.plde.Rs2E\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_796 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23611__230 clknet_1_0__leaf__10179_ VGND VGND VPWR VPWR net356 sky130_fd_sc_hd__inv_2
XFILLER_0_140_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_199_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22071_ rvcpu.dp.plem.WriteDataM\[6\] _09264_ _09265_ rvcpu.dp.plem.WriteDataM\[14\]
+ VGND VGND VPWR VPWR _09287_ sky130_fd_sc_hd__a22o_4
X_23218__868 clknet_1_1__leaf__10124_ VGND VGND VPWR VPWR net994 sky130_fd_sc_hd__inv_2
XFILLER_0_100_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31269_ clknet_leaf_35_clk _02972_ VGND VGND VPWR VPWR rvcpu.dp.plfd.InstrD\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21022_ _06851_ _08302_ _08305_ _08310_ VGND VGND VPWR VPWR _08311_ sky130_fd_sc_hd__a31o_1
XFILLER_0_61_1074 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25830_ rvcpu.dp.plfd.PCPlus4D\[22\] _11215_ _11142_ VGND VGND VPWR VPWR _11216_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_203_5363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_203_5374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25761_ _13823_ _13876_ _13706_ VGND VGND VPWR VPWR _11162_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_198_106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24712_ _10470_ net4251 _10561_ VGND VGND VPWR VPWR _10564_ sky130_fd_sc_hd__mux2_1
X_27500_ _12181_ VGND VGND VPWR VPWR _03608_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_195_5164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28480_ _12722_ VGND VGND VPWR VPWR _12723_ sky130_fd_sc_hd__buf_2
X_21924_ _08541_ _09157_ VGND VGND VPWR VPWR _09158_ sky130_fd_sc_hd__and2_1
X_25692_ _11047_ _11113_ VGND VGND VPWR VPWR _11118_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_195_5175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_195_5186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27431_ _12139_ VGND VGND VPWR VPWR _03581_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_182_Right_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24643_ _10525_ VGND VGND VPWR VPWR _02407_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_171_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21855_ rvcpu.dp.rf.reg_file_arr\[16\]\[25\] rvcpu.dp.rf.reg_file_arr\[17\]\[25\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[25\] rvcpu.dp.rf.reg_file_arr\[19\]\[25\] _08631_
+ _08632_ VGND VGND VPWR VPWR _09092_ sky130_fd_sc_hd__mux4_1
XFILLER_0_78_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27362_ _12099_ VGND VGND VPWR VPWR _03552_ sky130_fd_sc_hd__clkbuf_1
X_20806_ datamem.data_ram\[42\]\[30\] datamem.data_ram\[43\]\[30\] _07835_ VGND VGND
+ VPWR VPWR _08096_ sky130_fd_sc_hd__mux2_1
X_24574_ _10487_ VGND VGND VPWR VPWR _02376_ sky130_fd_sc_hd__clkbuf_1
X_21786_ rvcpu.dp.rf.reg_file_arr\[24\]\[21\] rvcpu.dp.rf.reg_file_arr\[25\]\[21\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[21\] rvcpu.dp.rf.reg_file_arr\[27\]\[21\] _08536_
+ _08693_ VGND VGND VPWR VPWR _09027_ sky130_fd_sc_hd__mux4_1
XFILLER_0_136_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26313_ _11489_ VGND VGND VPWR VPWR _03113_ sky130_fd_sc_hd__clkbuf_1
X_29101_ _13065_ VGND VGND VPWR VPWR _04325_ sky130_fd_sc_hd__clkbuf_1
X_27293_ _12036_ net1475 _12053_ _12059_ VGND VGND VPWR VPWR _03523_ sky130_fd_sc_hd__a31o_1
X_20737_ _08025_ _08026_ _07840_ VGND VGND VPWR VPWR _08027_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_154_4182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_4193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29032_ _12749_ net2253 _13020_ VGND VGND VPWR VPWR _13028_ sky130_fd_sc_hd__mux2_1
X_26244_ _11438_ _11458_ _11459_ _09478_ VGND VGND VPWR VPWR _03074_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_135_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_190_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20668_ datamem.data_ram\[48\]\[29\] _06811_ _06655_ datamem.data_ram\[49\]\[29\]
+ _07958_ VGND VGND VPWR VPWR _07959_ sky130_fd_sc_hd__o221a_1
XFILLER_0_135_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22407_ rvcpu.dp.rf.reg_file_arr\[0\]\[5\] rvcpu.dp.rf.reg_file_arr\[1\]\[5\] rvcpu.dp.rf.reg_file_arr\[2\]\[5\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[5\] _09463_ _09466_ VGND VGND VPWR VPWR _09568_ sky130_fd_sc_hd__mux4_1
X_26175_ _11424_ VGND VGND VPWR VPWR _03040_ sky130_fd_sc_hd__clkbuf_1
X_23387_ _10144_ VGND VGND VPWR VPWR _01532_ sky130_fd_sc_hd__clkbuf_1
X_20599_ datamem.data_ram\[5\]\[13\] _07037_ _06687_ datamem.data_ram\[4\]\[13\] VGND
+ VGND VPWR VPWR _07890_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_167_4510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25126_ _10468_ net3336 net87 VGND VGND VPWR VPWR _10795_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22338_ rvcpu.dp.rf.reg_file_arr\[4\]\[2\] rvcpu.dp.rf.reg_file_arr\[5\]\[2\] rvcpu.dp.rf.reg_file_arr\[6\]\[2\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[2\] _09464_ _09467_ VGND VGND VPWR VPWR _09502_ sky130_fd_sc_hd__mux4_1
XFILLER_0_108_1240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_638 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_163_4407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25057_ _10756_ net2831 _10752_ VGND VGND VPWR VPWR _10757_ sky130_fd_sc_hd__mux2_1
X_29934_ net304 _01669_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[16\]\[25\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_163_4418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22269_ rvcpu.dp.rf.reg_file_arr\[12\]\[0\] rvcpu.dp.rf.reg_file_arr\[13\]\[0\] rvcpu.dp.rf.reg_file_arr\[14\]\[0\]
+ rvcpu.dp.rf.reg_file_arr\[15\]\[0\] _09434_ _09382_ VGND VGND VPWR VPWR _09435_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_218_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29865_ net243 _01600_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[18\]\[28\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24197__36 clknet_1_0__leaf__10267_ VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__inv_2
X_16830_ net1924 _14449_ _04659_ VGND VGND VPWR VPWR _04663_ sky130_fd_sc_hd__mux2_1
X_28816_ _12910_ VGND VGND VPWR VPWR _04195_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_228_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29796_ net1142 _01531_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[20\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_16761_ _04626_ VGND VGND VPWR VPWR _01663_ sky130_fd_sc_hd__clkbuf_1
X_28747_ _12873_ VGND VGND VPWR VPWR _04163_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_219_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25959_ _11143_ VGND VGND VPWR VPWR _11302_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_122_3414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_3425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_139 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18500_ _05398_ _05688_ _05684_ VGND VGND VPWR VPWR _05862_ sky130_fd_sc_hd__and3_1
X_15712_ _13253_ VGND VGND VPWR VPWR _14179_ sky130_fd_sc_hd__buf_4
XFILLER_0_88_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19480_ _06679_ VGND VGND VPWR VPWR _06776_ sky130_fd_sc_hd__buf_8
X_16692_ _14156_ net3492 _04587_ VGND VGND VPWR VPWR _04590_ sky130_fd_sc_hd__mux2_1
XFILLER_0_220_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28678_ _12760_ net3378 _12832_ VGND VGND VPWR VPWR _12837_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_87_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18431_ _05747_ _05794_ VGND VGND VPWR VPWR _05795_ sky130_fd_sc_hd__or2_1
X_15643_ _14132_ VGND VGND VPWR VPWR _02187_ sky130_fd_sc_hd__clkbuf_1
X_27629_ _12249_ VGND VGND VPWR VPWR _03669_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18362_ _05726_ VGND VGND VPWR VPWR _05727_ sky130_fd_sc_hd__clkbuf_4
X_30640_ clknet_leaf_149_clk _02375_ VGND VGND VPWR VPWR datamem.data_ram\[51\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15574_ _14094_ VGND VGND VPWR VPWR _02218_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_83_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26500__53 clknet_1_0__leaf__11601_ VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__inv_2
XFILLER_0_51_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_201_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_189_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23323__963 clknet_1_0__leaf__10134_ VGND VGND VPWR VPWR net1089 sky130_fd_sc_hd__inv_2
XFILLER_0_7_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17313_ _04919_ VGND VGND VPWR VPWR _01388_ sky130_fd_sc_hd__clkbuf_1
X_30571_ clknet_leaf_138_clk _02306_ VGND VGND VPWR VPWR datamem.data_ram\[54\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18293_ _05363_ VGND VGND VPWR VPWR _05658_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_166_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_96_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32310_ clknet_leaf_271_clk _03732_ VGND VGND VPWR VPWR datamem.data_ram\[32\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17244_ _04882_ VGND VGND VPWR VPWR _01420_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_1080 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_226_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17175_ _14162_ net3856 _04840_ VGND VGND VPWR VPWR _04846_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32241_ clknet_leaf_227_clk _03663_ VGND VGND VPWR VPWR datamem.data_ram\[34\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_42_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16126_ _14405_ VGND VGND VPWR VPWR _01961_ sky130_fd_sc_hd__clkbuf_1
X_23102__781 clknet_1_1__leaf__10103_ VGND VGND VPWR VPWR net907 sky130_fd_sc_hd__inv_2
XFILLER_0_106_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32172_ clknet_leaf_226_clk _03594_ VGND VGND VPWR VPWR datamem.data_ram\[37\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_498 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31123_ clknet_leaf_110_clk _02858_ VGND VGND VPWR VPWR datamem.data_ram\[35\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_55_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16057_ net3257 _13238_ _14360_ VGND VGND VPWR VPWR _14369_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3109 rvcpu.dp.rf.reg_file_arr\[13\]\[24\] VGND VGND VPWR VPWR net4259 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15008_ _13344_ _13420_ _13410_ VGND VGND VPWR VPWR _13556_ sky130_fd_sc_hd__a21oi_1
X_31054_ clknet_leaf_114_clk _02789_ VGND VGND VPWR VPWR datamem.data_ram\[38\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2408 datamem.data_ram\[24\]\[27\] VGND VGND VPWR VPWR net3558 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2419 datamem.data_ram\[51\]\[18\] VGND VGND VPWR VPWR net3569 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30005_ clknet_leaf_267_clk _01740_ VGND VGND VPWR VPWR datamem.data_ram\[59\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_19816_ datamem.data_ram\[19\]\[9\] _06636_ _07110_ _06777_ VGND VGND VPWR VPWR _07111_
+ sky130_fd_sc_hd__o211a_1
Xhold1707 datamem.data_ram\[59\]\[21\] VGND VGND VPWR VPWR net2857 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1718 rvcpu.dp.rf.reg_file_arr\[6\]\[1\] VGND VGND VPWR VPWR net2868 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1729 datamem.data_ram\[37\]\[19\] VGND VGND VPWR VPWR net2879 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19747_ datamem.data_ram\[46\]\[25\] _06719_ _06657_ datamem.data_ram\[41\]\[25\]
+ VGND VGND VPWR VPWR _07042_ sky130_fd_sc_hd__o22a_1
X_16959_ _04719_ VGND VGND VPWR VPWR _04731_ sky130_fd_sc_hd__buf_4
XFILLER_0_56_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31956_ clknet_leaf_121_clk _03378_ VGND VGND VPWR VPWR datamem.data_ram\[55\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_19678_ datamem.data_ram\[48\]\[0\] _06973_ _06955_ datamem.data_ram\[52\]\[0\] VGND
+ VGND VPWR VPWR _06974_ sky130_fd_sc_hd__a22o_1
XFILLER_0_189_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18629_ _05900_ _05904_ _05675_ VGND VGND VPWR VPWR _05986_ sky130_fd_sc_hd__mux2_1
X_30907_ clknet_leaf_192_clk _02642_ VGND VGND VPWR VPWR datamem.data_ram\[41\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_31887_ clknet_leaf_114_clk _03341_ VGND VGND VPWR VPWR datamem.data_ram\[36\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_177_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_176_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_190_5050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21640_ _08531_ _08886_ _08888_ _08806_ VGND VGND VPWR VPWR _08889_ sky130_fd_sc_hd__o211a_1
X_30838_ clknet_leaf_280_clk _02573_ VGND VGND VPWR VPWR datamem.data_ram\[44\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_190_5061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_191_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_191_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21571_ _08823_ VGND VGND VPWR VPWR _01037_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_16_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30769_ clknet_leaf_261_clk _02504_ VGND VGND VPWR VPWR datamem.data_ram\[47\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_11 _06603_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23298__940 clknet_1_0__leaf__10132_ VGND VGND VPWR VPWR net1066 sky130_fd_sc_hd__inv_2
XANTENNA_22 _06620_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20522_ datamem.data_ram\[27\]\[21\] _07077_ _07809_ _07812_ VGND VGND VPWR VPWR
+ _07813_ sky130_fd_sc_hd__o211a_1
X_32508_ clknet_leaf_232_clk _03930_ VGND VGND VPWR VPWR datamem.data_ram\[24\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_33 _06654_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_170_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24290_ _10318_ VGND VGND VPWR VPWR _02261_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_44 _06678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_55 _06703_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_66 _06764_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_77 _06777_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_88 _06790_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20453_ datamem.data_ram\[10\]\[20\] _06728_ _06778_ datamem.data_ram\[8\]\[20\]
+ _07744_ VGND VGND VPWR VPWR _07745_ sky130_fd_sc_hd__o221a_1
XFILLER_0_15_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32439_ clknet_leaf_184_clk _03861_ VGND VGND VPWR VPWR datamem.data_ram\[27\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_99 _06862_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_1137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20384_ datamem.data_ram\[51\]\[28\] _06729_ _06668_ datamem.data_ram\[55\]\[28\]
+ _06676_ VGND VGND VPWR VPWR _07676_ sky130_fd_sc_hd__o221a_1
XFILLER_0_113_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22123_ _09329_ VGND VGND VPWR VPWR _09330_ sky130_fd_sc_hd__clkbuf_2
X_27980_ _09266_ VGND VGND VPWR VPWR _12447_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_101_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_205_5414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_205_5425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26931_ _11831_ net1586 _11841_ _11845_ VGND VGND VPWR VPWR _03375_ sky130_fd_sc_hd__a31o_1
X_22054_ _09274_ VGND VGND VPWR VPWR _01069_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_227_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2920 rvcpu.dp.rf.reg_file_arr\[2\]\[9\] VGND VGND VPWR VPWR net4070 sky130_fd_sc_hd__dlygate4sd3_1
X_21005_ datamem.data_ram\[22\]\[15\] _06624_ rvcpu.dp.plem.ALUResultM\[5\] VGND VGND
+ VPWR VPWR _08294_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_195_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2931 datamem.data_ram\[36\]\[27\] VGND VGND VPWR VPWR net4081 sky130_fd_sc_hd__dlygate4sd3_1
X_29650_ net996 _01385_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[24\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_26862_ _11681_ _11798_ VGND VGND VPWR VPWR _11801_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_197_5215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_197_5226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2942 rvcpu.dp.rf.reg_file_arr\[26\]\[9\] VGND VGND VPWR VPWR net4092 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2953 datamem.data_ram\[57\]\[22\] VGND VGND VPWR VPWR net4103 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2964 rvcpu.dp.rf.reg_file_arr\[13\]\[21\] VGND VGND VPWR VPWR net4114 sky130_fd_sc_hd__dlygate4sd3_1
X_28601_ _10777_ _12602_ _12795_ VGND VGND VPWR VPWR _12796_ sky130_fd_sc_hd__a21oi_4
X_25813_ _11200_ _11201_ _11149_ VGND VGND VPWR VPWR _11202_ sky130_fd_sc_hd__o21ai_1
Xhold2975 rvcpu.dp.rf.reg_file_arr\[28\]\[31\] VGND VGND VPWR VPWR net4125 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_214_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26793_ _11672_ _11749_ VGND VGND VPWR VPWR _11759_ sky130_fd_sc_hd__and2_1
Xhold2986 datamem.data_ram\[57\]\[16\] VGND VGND VPWR VPWR net4136 sky130_fd_sc_hd__dlygate4sd3_1
X_29581_ net935 _01316_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[26\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_203_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2997 datamem.data_ram\[4\]\[16\] VGND VGND VPWR VPWR net4147 sky130_fd_sc_hd__dlygate4sd3_1
X_25744_ _08598_ VGND VGND VPWR VPWR _11149_ sky130_fd_sc_hd__buf_2
X_28532_ _12756_ net2369 _12752_ VGND VGND VPWR VPWR _12757_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23804__388 clknet_1_1__leaf__10206_ VGND VGND VPWR VPWR net514 sky130_fd_sc_hd__inv_2
Xmax_cap35 _10995_ VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_2
Xmax_cap46 _12564_ VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_4
XFILLER_0_98_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_223_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_214_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap57 _10829_ VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__buf_4
X_21907_ _08817_ _09139_ _09141_ _08700_ VGND VGND VPWR VPWR _09142_ sky130_fd_sc_hd__a211o_1
X_25675_ _11091_ _11098_ VGND VGND VPWR VPWR _11107_ sky130_fd_sc_hd__and2_1
X_28463_ _12447_ net2651 _12713_ VGND VGND VPWR VPWR _12714_ sky130_fd_sc_hd__mux2_1
X_22887_ _10022_ VGND VGND VPWR VPWR _01154_ sky130_fd_sc_hd__clkbuf_1
Xmax_cap79 _12261_ VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__buf_4
XFILLER_0_211_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_1249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_4233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_4244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27414_ _09235_ VGND VGND VPWR VPWR _12128_ sky130_fd_sc_hd__clkbuf_2
X_24626_ _10448_ net3666 _10511_ VGND VGND VPWR VPWR _10516_ sky130_fd_sc_hd__mux2_1
X_28394_ _12673_ VGND VGND VPWR VPWR _04010_ sky130_fd_sc_hd__clkbuf_1
X_21838_ rvcpu.dp.rf.reg_file_arr\[20\]\[24\] rvcpu.dp.rf.reg_file_arr\[21\]\[24\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[24\] rvcpu.dp.rf.reg_file_arr\[23\]\[24\] _08525_
+ _08528_ VGND VGND VPWR VPWR _09076_ sky130_fd_sc_hd__mux4_1
XFILLER_0_214_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_210_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23919__475 clknet_1_1__leaf__10226_ VGND VGND VPWR VPWR net601 sky130_fd_sc_hd__inv_2
XFILLER_0_214_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27345_ _12088_ VGND VGND VPWR VPWR _03546_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_183_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24557_ _10477_ VGND VGND VPWR VPWR _02369_ sky130_fd_sc_hd__clkbuf_1
X_21769_ _08798_ _09008_ _09010_ _08512_ VGND VGND VPWR VPWR _09011_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_50_clk clknet_5_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_50_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_194_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23508_ _10142_ _09229_ _09361_ VGND VGND VPWR VPWR _10162_ sky130_fd_sc_hd__a21oi_4
X_23618__236 clknet_1_0__leaf__10180_ VGND VGND VPWR VPWR net362 sky130_fd_sc_hd__inv_2
X_15290_ _13706_ _13825_ _13826_ _13827_ _13429_ VGND VGND VPWR VPWR _13828_ sky130_fd_sc_hd__a32o_1
X_27276_ _12049_ VGND VGND VPWR VPWR _03516_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_184_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24488_ _10434_ VGND VGND VPWR VPWR _02343_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29015_ _10075_ _13010_ VGND VGND VPWR VPWR _13019_ sky130_fd_sc_hd__and2_1
XFILLER_0_191_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26227_ _11378_ VGND VGND VPWR VPWR _11452_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_3251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_3262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26158_ rvcpu.dp.plfd.InstrD\[7\] _11408_ VGND VGND VPWR VPWR _11416_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_186_4952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_186_4963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_111_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25109_ _10727_ net4039 _10784_ VGND VGND VPWR VPWR _10786_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_111_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26089_ _06567_ _11367_ _11375_ _11379_ _11372_ VGND VGND VPWR VPWR _02998_ sky130_fd_sc_hd__o41a_1
X_18980_ _05303_ _05785_ _06108_ _05302_ VGND VGND VPWR VPWR _06316_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_221_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17931_ _05302_ _05303_ VGND VGND VPWR VPWR _05304_ sky130_fd_sc_hd__or2_1
X_29917_ net287 _01652_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[16\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17862_ rvcpu.dp.plde.ALUControlE\[3\] rvcpu.dp.plde.ALUControlE\[2\] VGND VGND VPWR
+ VPWR _05236_ sky130_fd_sc_hd__or2_1
X_29848_ net226 _01583_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[18\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_89_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_89_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19601_ _06751_ _06891_ _06896_ VGND VGND VPWR VPWR _06897_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_145_3970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16813_ net4080 _14432_ _04648_ VGND VGND VPWR VPWR _04654_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_145_3981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17793_ _05179_ _05180_ rvcpu.dp.plde.RD2E\[3\] VGND VGND VPWR VPWR _05188_ sky130_fd_sc_hd__a21boi_1
X_29779_ net1125 _01514_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[20\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_85_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31810_ clknet_leaf_109_clk _03264_ VGND VGND VPWR VPWR datamem.data_ram\[17\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_19532_ _06812_ VGND VGND VPWR VPWR _06828_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_85_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16744_ _04617_ VGND VGND VPWR VPWR _01671_ sky130_fd_sc_hd__clkbuf_1
X_32790_ clknet_leaf_283_clk _04212_ VGND VGND VPWR VPWR datamem.data_ram\[14\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_141_3878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_141_3889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19463_ datamem.data_ram\[59\]\[16\] _06739_ _06755_ _06758_ VGND VGND VPWR VPWR
+ _06759_ sky130_fd_sc_hd__o211a_1
X_23779__365 clknet_1_1__leaf__10204_ VGND VGND VPWR VPWR net491 sky130_fd_sc_hd__inv_2
X_31741_ net190 _03199_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[9\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16675_ _14139_ net2829 _04576_ VGND VGND VPWR VPWR _04581_ sky130_fd_sc_hd__mux2_1
X_18414_ _05408_ _05606_ net102 _05604_ _05684_ _05689_ VGND VGND VPWR VPWR _05778_
+ sky130_fd_sc_hd__mux4_1
X_15626_ _14121_ VGND VGND VPWR VPWR _02193_ sky130_fd_sc_hd__clkbuf_1
X_31672_ clknet_leaf_69_clk net1276 VGND VGND VPWR VPWR rvcpu.dp.plmw.ALUResultW\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_19394_ _06689_ VGND VGND VPWR VPWR _06690_ sky130_fd_sc_hd__buf_6
XFILLER_0_75_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_185_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18345_ _05709_ VGND VGND VPWR VPWR _05710_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30623_ clknet_leaf_178_clk _02358_ VGND VGND VPWR VPWR datamem.data_ram\[52\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_15557_ _13496_ _14079_ _14080_ VGND VGND VPWR VPWR _14081_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_44_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_41_clk clknet_5_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_41_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_12_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_204_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15488_ _13358_ _13424_ _13689_ VGND VGND VPWR VPWR _14017_ sky130_fd_sc_hd__or3b_1
X_18276_ _05630_ _05631_ _05640_ VGND VGND VPWR VPWR _05641_ sky130_fd_sc_hd__a21o_1
XFILLER_0_127_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30554_ clknet_leaf_178_clk _02289_ VGND VGND VPWR VPWR datamem.data_ram\[55\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17227_ _04873_ VGND VGND VPWR VPWR _01428_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30485_ clknet_leaf_206_clk _02220_ VGND VGND VPWR VPWR datamem.data_ram\[57\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32224_ clknet_leaf_201_clk _03646_ VGND VGND VPWR VPWR datamem.data_ram\[35\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold804 datamem.data_ram\[12\]\[23\] VGND VGND VPWR VPWR net1954 sky130_fd_sc_hd__dlygate4sd3_1
X_17158_ _14145_ net3273 _04829_ VGND VGND VPWR VPWR _04837_ sky130_fd_sc_hd__mux2_1
Xhold815 rvcpu.dp.rf.reg_file_arr\[10\]\[28\] VGND VGND VPWR VPWR net1965 sky130_fd_sc_hd__dlygate4sd3_1
Xhold826 rvcpu.dp.rf.reg_file_arr\[30\]\[23\] VGND VGND VPWR VPWR net1976 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold837 datamem.data_ram\[12\]\[31\] VGND VGND VPWR VPWR net1987 sky130_fd_sc_hd__dlygate4sd3_1
X_16109_ net1950 _13213_ _14396_ VGND VGND VPWR VPWR _14397_ sky130_fd_sc_hd__mux2_1
Xhold848 datamem.data_ram\[5\]\[30\] VGND VGND VPWR VPWR net1998 sky130_fd_sc_hd__dlygate4sd3_1
X_32155_ clknet_leaf_167_clk _03577_ VGND VGND VPWR VPWR datamem.data_ram\[38\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_17089_ _04800_ VGND VGND VPWR VPWR _01493_ sky130_fd_sc_hd__clkbuf_1
Xhold859 datamem.data_ram\[27\]\[23\] VGND VGND VPWR VPWR net2009 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1023 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31106_ clknet_leaf_108_clk _02841_ VGND VGND VPWR VPWR datamem.data_ram\[19\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_196_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32086_ clknet_leaf_57_clk _03508_ VGND VGND VPWR VPWR datamem.data_ram\[47\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2205 rvcpu.dp.rf.reg_file_arr\[13\]\[5\] VGND VGND VPWR VPWR net3355 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2216 datamem.data_ram\[57\]\[27\] VGND VGND VPWR VPWR net3366 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31037_ clknet_leaf_60_clk _02772_ VGND VGND VPWR VPWR datamem.data_ram\[41\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2227 datamem.data_ram\[19\]\[25\] VGND VGND VPWR VPWR net3377 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2238 datamem.data_ram\[25\]\[17\] VGND VGND VPWR VPWR net3388 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_200_5300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1504 datamem.data_ram\[15\]\[19\] VGND VGND VPWR VPWR net2654 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2249 rvcpu.dp.rf.reg_file_arr\[8\]\[16\] VGND VGND VPWR VPWR net3399 sky130_fd_sc_hd__dlygate4sd3_1
X_24176__17 clknet_1_1__leaf__10265_ VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__inv_2
Xhold1515 rvcpu.dp.rf.reg_file_arr\[6\]\[5\] VGND VGND VPWR VPWR net2665 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_596 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1526 datamem.data_ram\[25\]\[30\] VGND VGND VPWR VPWR net2676 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1537 datamem.data_ram\[58\]\[29\] VGND VGND VPWR VPWR net2687 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1548 datamem.data_ram\[12\]\[30\] VGND VGND VPWR VPWR net2698 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1559 datamem.data_ram\[61\]\[14\] VGND VGND VPWR VPWR net2709 sky130_fd_sc_hd__dlygate4sd3_1
X_22810_ rvcpu.dp.rf.reg_file_arr\[8\]\[26\] rvcpu.dp.rf.reg_file_arr\[10\]\[26\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[26\] rvcpu.dp.rf.reg_file_arr\[11\]\[26\] _09424_
+ _09485_ VGND VGND VPWR VPWR _09950_ sky130_fd_sc_hd__mux4_1
XFILLER_0_28_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_192_5101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_192_5112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32988_ clknet_leaf_206_clk _04410_ VGND VGND VPWR VPWR datamem.data_ram\[62\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22741_ rvcpu.dp.rf.reg_file_arr\[16\]\[23\] rvcpu.dp.rf.reg_file_arr\[17\]\[23\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[23\] rvcpu.dp.rf.reg_file_arr\[19\]\[23\] _09517_
+ _09513_ VGND VGND VPWR VPWR _09884_ sky130_fd_sc_hd__mux4_1
X_31939_ clknet_leaf_120_clk _03361_ VGND VGND VPWR VPWR datamem.data_ram\[59\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25460_ _10405_ _10985_ VGND VGND VPWR VPWR _10986_ sky130_fd_sc_hd__and2_1
X_22672_ _09391_ _09818_ VGND VGND VPWR VPWR _09819_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_176_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24411_ _09266_ VGND VGND VPWR VPWR _10385_ sky130_fd_sc_hd__buf_2
X_21623_ rvcpu.dp.rf.reg_file_arr\[8\]\[12\] rvcpu.dp.rf.reg_file_arr\[10\]\[12\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[12\] rvcpu.dp.rf.reg_file_arr\[11\]\[12\] _08534_
+ _08537_ VGND VGND VPWR VPWR _08873_ sky130_fd_sc_hd__mux4_2
X_25391_ _10948_ VGND VGND VPWR VPWR _10949_ sky130_fd_sc_hd__clkbuf_2
X_23109__787 clknet_1_0__leaf__10104_ VGND VGND VPWR VPWR net913 sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_32_clk clknet_5_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_32_clk sky130_fd_sc_hd__clkbuf_8
X_27130_ _10047_ VGND VGND VPWR VPWR _11965_ sky130_fd_sc_hd__buf_2
XFILLER_0_90_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_151_4130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24342_ _10325_ _10347_ _10269_ VGND VGND VPWR VPWR _10348_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_30_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21554_ _08531_ _08803_ _08805_ _08806_ VGND VGND VPWR VPWR _08807_ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_209_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27061_ _07077_ _11109_ _11839_ VGND VGND VPWR VPWR _11922_ sky130_fd_sc_hd__or3_1
X_20505_ datamem.data_ram\[45\]\[21\] _07019_ _07792_ _07795_ VGND VGND VPWR VPWR
+ _07796_ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24273_ _10309_ VGND VGND VPWR VPWR _02253_ sky130_fd_sc_hd__clkbuf_1
X_21485_ rvcpu.dp.rf.reg_file_arr\[20\]\[6\] rvcpu.dp.rf.reg_file_arr\[21\]\[6\] rvcpu.dp.rf.reg_file_arr\[22\]\[6\]
+ rvcpu.dp.rf.reg_file_arr\[23\]\[6\] _08631_ _08632_ VGND VGND VPWR VPWR _08741_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_200_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26012_ net1296 _11329_ _11325_ _11331_ VGND VGND VPWR VPWR _02970_ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20436_ datamem.data_ram\[22\]\[12\] _07085_ _07726_ _07727_ VGND VGND VPWR VPWR
+ _07728_ sky130_fd_sc_hd__o211a_1
XFILLER_0_209_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__11601_ clknet_0__11601_ VGND VGND VPWR VPWR clknet_1_1__leaf__11601_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_228_5970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20367_ datamem.data_ram\[39\]\[28\] _06668_ _06654_ datamem.data_ram\[33\]\[28\]
+ VGND VGND VPWR VPWR _07659_ sky130_fd_sc_hd__o22a_1
Xclkload280 clknet_1_1__leaf__10260_ VGND VGND VPWR VPWR clkload280/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload291 clknet_1_1__leaf__10227_ VGND VGND VPWR VPWR clkload291/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_149_4070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_4081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22106_ rvcpu.dp.plem.WriteDataM\[4\] _08488_ _09293_ _09295_ rvcpu.dp.plem.WriteDataM\[12\]
+ VGND VGND VPWR VPWR _09316_ sky130_fd_sc_hd__a32o_1
XFILLER_0_219_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27963_ _12435_ net4204 _12431_ VGND VGND VPWR VPWR _12436_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_224_5867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20298_ datamem.data_ram\[5\]\[19\] _06768_ _06699_ datamem.data_ram\[1\]\[19\] VGND
+ VGND VPWR VPWR _07591_ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_99_clk clknet_5_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_99_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_224_5878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29702_ net1048 _01437_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[22\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_26914_ _11833_ _11823_ VGND VGND VPWR VPWR _11834_ sky130_fd_sc_hd__and2_1
X_22037_ _09259_ VGND VGND VPWR VPWR _09260_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_8_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27894_ _11972_ _12394_ VGND VGND VPWR VPWR _12398_ sky130_fd_sc_hd__and2_1
XFILLER_0_215_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2750 rvcpu.dp.rf.reg_file_arr\[30\]\[30\] VGND VGND VPWR VPWR net3900 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29633_ clknet_leaf_147_clk _01368_ VGND VGND VPWR VPWR datamem.data_ram\[5\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26845_ _11781_ net1788 _11785_ _11790_ VGND VGND VPWR VPWR _03344_ sky130_fd_sc_hd__a31o_1
Xhold2761 datamem.data_ram\[53\]\[25\] VGND VGND VPWR VPWR net3911 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2772 datamem.data_ram\[29\]\[8\] VGND VGND VPWR VPWR net3922 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2783 datamem.data_ram\[44\]\[28\] VGND VGND VPWR VPWR net3933 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2794 datamem.data_ram\[17\]\[31\] VGND VGND VPWR VPWR net3944 sky130_fd_sc_hd__dlygate4sd3_1
X_14790_ _13342_ VGND VGND VPWR VPWR _13343_ sky130_fd_sc_hd__buf_2
X_29564_ net918 _01299_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[27\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_26776_ _10325_ _08066_ _11609_ VGND VGND VPWR VPWR _11749_ sky130_fd_sc_hd__and3_2
XFILLER_0_98_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_216_1238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28515_ _09284_ VGND VGND VPWR VPWR _12745_ sky130_fd_sc_hd__clkbuf_2
X_22939_ _10056_ net1429 _10046_ _10068_ VGND VGND VPWR VPWR _01160_ sky130_fd_sc_hd__a31o_1
XFILLER_0_35_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25727_ _11137_ VGND VGND VPWR VPWR _02879_ sky130_fd_sc_hd__clkbuf_1
X_29495_ net857 _01230_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[28\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_80_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28446_ _12430_ net3006 _12704_ VGND VGND VPWR VPWR _12705_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16460_ _04464_ _04465_ VGND VGND VPWR VPWR _04466_ sky130_fd_sc_hd__and2_2
X_25658_ _07077_ _10918_ _10897_ VGND VGND VPWR VPWR _11096_ sky130_fd_sc_hd__or3_1
XFILLER_0_210_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_175_4686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15411_ _13298_ _13681_ _13507_ VGND VGND VPWR VPWR _13943_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_175_4697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23852__415 clknet_1_1__leaf__10219_ VGND VGND VPWR VPWR net541 sky130_fd_sc_hd__inv_2
X_16391_ _14560_ VGND VGND VPWR VPWR _14561_ sky130_fd_sc_hd__buf_4
X_24609_ _10474_ net3354 _10502_ VGND VGND VPWR VPWR _10507_ sky130_fd_sc_hd__mux2_1
X_25589_ _10408_ _11055_ VGND VGND VPWR VPWR _11058_ sky130_fd_sc_hd__and2_1
XFILLER_0_149_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_3302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28377_ _12365_ net3654 _12659_ VGND VGND VPWR VPWR _12664_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_23_clk clknet_5_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_23_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_117_3313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15342_ _13608_ _13528_ _13539_ VGND VGND VPWR VPWR _13878_ sky130_fd_sc_hd__a21o_1
X_18130_ _05494_ _05495_ VGND VGND VPWR VPWR _05496_ sky130_fd_sc_hd__and2_1
X_27328_ _10064_ _12078_ _12079_ net1287 VGND VGND VPWR VPWR _03538_ sky130_fd_sc_hd__o22a_1
XFILLER_0_170_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15273_ _13307_ _13689_ _13811_ VGND VGND VPWR VPWR _13812_ sky130_fd_sc_hd__a21o_1
XFILLER_0_163_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18061_ rvcpu.dp.plde.RD1E\[9\] _05267_ _05271_ _13250_ _05428_ VGND VGND VPWR VPWR
+ _05429_ sky130_fd_sc_hd__a221oi_2
X_27259_ _10064_ net52 _12042_ net1302 VGND VGND VPWR VPWR _03506_ sky130_fd_sc_hd__a22o_1
XFILLER_0_184_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_227_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17012_ net2969 _14426_ _04757_ VGND VGND VPWR VPWR _04760_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_78_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30270_ net624 _02005_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[6\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18963_ _05543_ _05728_ _06108_ _05542_ VGND VGND VPWR VPWR _06300_ sky130_fd_sc_hd__a22o_1
X_17914_ rvcpu.dp.plde.ImmExtE\[30\] rvcpu.dp.SrcBFW_Mux.y\[30\] _05279_ VGND VGND
+ VPWR VPWR _05287_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18894_ _05467_ _05728_ _06179_ _06234_ _06235_ VGND VGND VPWR VPWR _06236_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_119_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_143_3918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32911_ clknet_leaf_278_clk _04333_ VGND VGND VPWR VPWR datamem.data_ram\[7\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_17845_ _05224_ VGND VGND VPWR VPWR rvcpu.dp.SrcBFW_Mux.y\[15\] sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_20_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_201_Left_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32842_ clknet_leaf_96_clk _04264_ VGND VGND VPWR VPWR datamem.data_ram\[7\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_17776_ _05158_ _05164_ _05167_ _05170_ VGND VGND VPWR VPWR _05174_ sky130_fd_sc_hd__or4b_2
X_14988_ _13393_ _13484_ VGND VGND VPWR VPWR _13536_ sky130_fd_sc_hd__nor2_1
XFILLER_0_191_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_178_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19515_ _06644_ VGND VGND VPWR VPWR _06811_ sky130_fd_sc_hd__buf_4
X_16727_ _14191_ net4187 _04598_ VGND VGND VPWR VPWR _04608_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_18_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32773_ clknet_leaf_236_clk _04195_ VGND VGND VPWR VPWR datamem.data_ram\[14\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_46_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19446_ _06741_ VGND VGND VPWR VPWR _06742_ sky130_fd_sc_hd__buf_8
X_31724_ net173 _03182_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[9\]\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_102_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16658_ _04571_ VGND VGND VPWR VPWR _01711_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_102_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23028__730 clknet_1_1__leaf__10088_ VGND VGND VPWR VPWR net856 sky130_fd_sc_hd__inv_2
XFILLER_0_9_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15609_ _14112_ VGND VGND VPWR VPWR _02201_ sky130_fd_sc_hd__clkbuf_1
X_31655_ clknet_leaf_63_clk net4272 VGND VGND VPWR VPWR rvcpu.dp.plmw.ALUResultW\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_19377_ datamem.data_ram\[13\]\[16\] _06665_ _06672_ datamem.data_ram\[15\]\[16\]
+ VGND VGND VPWR VPWR _06673_ sky130_fd_sc_hd__o22a_1
X_16589_ _04534_ VGND VGND VPWR VPWR _01751_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_174_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_14_clk clknet_5_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_8_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18328_ _05692_ VGND VGND VPWR VPWR _05693_ sky130_fd_sc_hd__buf_2
X_30606_ clknet_leaf_207_clk _02341_ VGND VGND VPWR VPWR datamem.data_ram\[52\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_210_Left_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31586_ clknet_leaf_64_clk net1167 VGND VGND VPWR VPWR rvcpu.dp.plmw.PCPlus4W\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18259_ _05621_ _05470_ _05623_ VGND VGND VPWR VPWR _05624_ sky130_fd_sc_hd__o21a_1
X_30537_ clknet_leaf_218_clk _02272_ VGND VGND VPWR VPWR datamem.data_ram\[55\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_839 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21270_ _08531_ VGND VGND VPWR VPWR _08532_ sky130_fd_sc_hd__clkbuf_4
Xhold601 datamem.data_ram\[37\]\[5\] VGND VGND VPWR VPWR net1751 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30468_ net146 _02203_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[19\]\[15\] sky130_fd_sc_hd__dfxtp_1
Xhold612 rvcpu.dp.plfd.InstrD\[10\] VGND VGND VPWR VPWR net1762 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20221_ datamem.data_ram\[19\]\[3\] _06961_ _06948_ datamem.data_ram\[17\]\[3\] VGND
+ VGND VPWR VPWR _07514_ sky130_fd_sc_hd__a22o_1
Xhold623 datamem.data_ram\[54\]\[3\] VGND VGND VPWR VPWR net1773 sky130_fd_sc_hd__dlygate4sd3_1
X_32207_ clknet_leaf_88_clk _03629_ VGND VGND VPWR VPWR datamem.data_ram\[36\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold634 datamem.data_ram\[26\]\[1\] VGND VGND VPWR VPWR net1784 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold645 rvcpu.dp.pcreg.q\[31\] VGND VGND VPWR VPWR net1795 sky130_fd_sc_hd__dlygate4sd3_1
Xhold656 datamem.data_ram\[15\]\[0\] VGND VGND VPWR VPWR net1806 sky130_fd_sc_hd__dlygate4sd3_1
X_30399_ net737 _02134_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[31\]\[10\] sky130_fd_sc_hd__dfxtp_1
Xhold667 datamem.data_ram\[8\]\[2\] VGND VGND VPWR VPWR net1817 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_204_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold678 datamem.data_ram\[24\]\[7\] VGND VGND VPWR VPWR net1828 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20152_ datamem.data_ram\[50\]\[27\] _06609_ _06632_ datamem.data_ram\[51\]\[27\]
+ _06677_ VGND VGND VPWR VPWR _07445_ sky130_fd_sc_hd__o221a_1
X_32138_ clknet_leaf_273_clk _03560_ VGND VGND VPWR VPWR datamem.data_ram\[39\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold689 datamem.data_ram\[16\]\[4\] VGND VGND VPWR VPWR net1839 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2002 datamem.data_ram\[19\]\[19\] VGND VGND VPWR VPWR net3152 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24960_ _10699_ VGND VGND VPWR VPWR _02550_ sky130_fd_sc_hd__clkbuf_1
Xhold2013 rvcpu.dp.rf.reg_file_arr\[28\]\[8\] VGND VGND VPWR VPWR net3163 sky130_fd_sc_hd__dlygate4sd3_1
X_32069_ clknet_leaf_122_clk _03491_ VGND VGND VPWR VPWR datamem.data_ram\[29\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2024 rvcpu.dp.rf.reg_file_arr\[16\]\[6\] VGND VGND VPWR VPWR net3174 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20083_ _06679_ _07374_ _07376_ VGND VGND VPWR VPWR _07377_ sky130_fd_sc_hd__and3_1
Xhold2035 datamem.data_ram\[0\]\[20\] VGND VGND VPWR VPWR net3185 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_209_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1301 rvcpu.dp.rf.reg_file_arr\[20\]\[22\] VGND VGND VPWR VPWR net2451 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2046 datamem.data_ram\[38\]\[10\] VGND VGND VPWR VPWR net3196 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1312 rvcpu.dp.rf.reg_file_arr\[11\]\[2\] VGND VGND VPWR VPWR net2462 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2057 datamem.data_ram\[50\]\[11\] VGND VGND VPWR VPWR net3207 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1323 datamem.data_ram\[3\]\[19\] VGND VGND VPWR VPWR net2473 sky130_fd_sc_hd__dlygate4sd3_1
X_24891_ _10662_ VGND VGND VPWR VPWR _02518_ sky130_fd_sc_hd__clkbuf_1
Xhold2068 rvcpu.dp.rf.reg_file_arr\[23\]\[28\] VGND VGND VPWR VPWR net3218 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1334 rvcpu.dp.rf.reg_file_arr\[13\]\[19\] VGND VGND VPWR VPWR net2484 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2079 datamem.data_ram\[51\]\[8\] VGND VGND VPWR VPWR net3229 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1345 datamem.data_ram\[4\]\[28\] VGND VGND VPWR VPWR net2495 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26630_ _10073_ _11659_ _11660_ net1309 VGND VGND VPWR VPWR _03259_ sky130_fd_sc_hd__a22o_1
X_23842_ _10217_ VGND VGND VPWR VPWR _01914_ sky130_fd_sc_hd__clkbuf_1
Xhold1356 datamem.data_ram\[32\]\[12\] VGND VGND VPWR VPWR net2506 sky130_fd_sc_hd__dlygate4sd3_1
X_24092__601 clknet_1_0__leaf__10248_ VGND VGND VPWR VPWR net727 sky130_fd_sc_hd__inv_2
XFILLER_0_174_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1367 rvcpu.dp.rf.reg_file_arr\[10\]\[30\] VGND VGND VPWR VPWR net2517 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1378 datamem.data_ram\[11\]\[16\] VGND VGND VPWR VPWR net2528 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_192_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1389 datamem.data_ram\[10\]\[14\] VGND VGND VPWR VPWR net2539 sky130_fd_sc_hd__dlygate4sd3_1
X_23263__909 clknet_1_1__leaf__10128_ VGND VGND VPWR VPWR net1035 sky130_fd_sc_hd__inv_2
XANTENNA_507 _13212_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_1_1__f__10130_ clknet_0__10130_ VGND VGND VPWR VPWR clknet_1_1__leaf__10130_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_196_226 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_518 _13228_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26561_ _11625_ VGND VGND VPWR VPWR _03225_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_529 _13423_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20985_ _06928_ _08273_ VGND VGND VPWR VPWR _08274_ sky130_fd_sc_hd__or2_1
XFILLER_0_178_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28300_ _12601_ _12622_ _12573_ VGND VGND VPWR VPWR _12623_ sky130_fd_sc_hd__a21oi_1
X_25512_ _10991_ net1461 _11009_ _11012_ VGND VGND VPWR VPWR _02789_ sky130_fd_sc_hd__a31o_1
X_22724_ rvcpu.dp.rf.reg_file_arr\[20\]\[22\] rvcpu.dp.rf.reg_file_arr\[21\]\[22\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[22\] rvcpu.dp.rf.reg_file_arr\[23\]\[22\] _09406_
+ _09395_ VGND VGND VPWR VPWR _09868_ sky130_fd_sc_hd__mux4_1
Xclkbuf_0__10161_ _10161_ VGND VGND VPWR VPWR clknet_0__10161_ sky130_fd_sc_hd__clkbuf_16
X_29280_ _13161_ VGND VGND VPWR VPWR _04408_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28231_ _12433_ net3808 _12583_ VGND VGND VPWR VPWR _12585_ sky130_fd_sc_hd__mux2_1
X_25443_ _10766_ net3414 _10970_ VGND VGND VPWR VPWR _10978_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_217_5693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22655_ rvcpu.dp.rf.reg_file_arr\[28\]\[18\] rvcpu.dp.rf.reg_file_arr\[30\]\[18\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[18\] rvcpu.dp.rf.reg_file_arr\[31\]\[18\] _09400_
+ _09484_ VGND VGND VPWR VPWR _09803_ sky130_fd_sc_hd__mux4_1
XFILLER_0_47_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21606_ rvcpu.dp.rf.reg_file_arr\[4\]\[11\] rvcpu.dp.rf.reg_file_arr\[5\]\[11\] rvcpu.dp.rf.reg_file_arr\[6\]\[11\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[11\] _08687_ _08856_ VGND VGND VPWR VPWR _08857_
+ sky130_fd_sc_hd__mux4_1
X_25374_ _10408_ _10936_ VGND VGND VPWR VPWR _10939_ sky130_fd_sc_hd__and2_1
X_28162_ _12359_ net2738 _12546_ VGND VGND VPWR VPWR _12548_ sky130_fd_sc_hd__mux2_1
X_22586_ _09461_ _09735_ _09737_ _09489_ VGND VGND VPWR VPWR _09738_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_170_4572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27113_ _11825_ _11953_ VGND VGND VPWR VPWR _11955_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_170_4583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24325_ _09224_ net4372 _10338_ VGND VGND VPWR VPWR _10339_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28093_ _12511_ VGND VGND VPWR VPWR _03871_ sky130_fd_sc_hd__clkbuf_1
X_21537_ rvcpu.dp.rf.reg_file_arr\[12\]\[8\] rvcpu.dp.rf.reg_file_arr\[13\]\[8\] rvcpu.dp.rf.reg_file_arr\[14\]\[8\]
+ rvcpu.dp.rf.reg_file_arr\[15\]\[8\] _08567_ _08570_ VGND VGND VPWR VPWR _08791_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_8_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27044_ _11904_ net1837 _11910_ _11912_ VGND VGND VPWR VPWR _03421_ sky130_fd_sc_hd__a31o_1
XFILLER_0_44_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24256_ _10300_ VGND VGND VPWR VPWR _02245_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21468_ _08531_ VGND VGND VPWR VPWR _08725_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_181_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_226_5918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_587 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_226_5929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20419_ datamem.data_ram\[51\]\[12\] _06633_ _07710_ _06678_ VGND VGND VPWR VPWR
+ _07711_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_147_4018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_4029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21399_ rvcpu.dp.rf.reg_file_arr\[24\]\[2\] rvcpu.dp.rf.reg_file_arr\[25\]\[2\] rvcpu.dp.rf.reg_file_arr\[26\]\[2\]
+ rvcpu.dp.rf.reg_file_arr\[27\]\[2\] _08517_ _08519_ VGND VGND VPWR VPWR _08659_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_31_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_73_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28995_ _12702_ net4144 _12999_ VGND VGND VPWR VPWR _13007_ sky130_fd_sc_hd__mux2_1
XFILLER_0_219_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_222_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27946_ _12425_ VGND VGND VPWR VPWR _03810_ sky130_fd_sc_hd__clkbuf_1
X_23069_ _10096_ VGND VGND VPWR VPWR _01262_ sky130_fd_sc_hd__clkbuf_1
X_15960_ net2559 _13198_ _14311_ VGND VGND VPWR VPWR _14317_ sky130_fd_sc_hd__mux2_1
Xhold3270 rvcpu.dp.rf.reg_file_arr\[24\]\[28\] VGND VGND VPWR VPWR net4420 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_842 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14911_ _13458_ _13360_ _13327_ _13460_ VGND VGND VPWR VPWR _13461_ sky130_fd_sc_hd__a2bb2o_1
Xhold3281 datamem.data_ram\[52\]\[18\] VGND VGND VPWR VPWR net4431 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3292 datamem.data_ram\[2\]\[17\] VGND VGND VPWR VPWR net4442 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27877_ _12387_ VGND VGND VPWR VPWR _03779_ sky130_fd_sc_hd__clkbuf_1
X_15891_ _14280_ VGND VGND VPWR VPWR _02079_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_106_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2580 datamem.data_ram\[4\]\[27\] VGND VGND VPWR VPWR net3730 sky130_fd_sc_hd__dlygate4sd3_1
X_17630_ _05087_ VGND VGND VPWR VPWR _01223_ sky130_fd_sc_hd__clkbuf_1
X_29616_ net970 _01351_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[25\]\[19\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_106_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26828_ _11687_ _11774_ VGND VGND VPWR VPWR _11780_ sky130_fd_sc_hd__and2_1
X_14842_ _13332_ _13392_ _13394_ _13304_ _13314_ VGND VGND VPWR VPWR _13395_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_192_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2591 rvcpu.dp.rf.reg_file_arr\[28\]\[26\] VGND VGND VPWR VPWR net3741 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_37_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_177_4737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1890 datamem.data_ram\[12\]\[24\] VGND VGND VPWR VPWR net3040 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_177_4748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17561_ _13195_ net4254 _05046_ VGND VGND VPWR VPWR _05051_ sky130_fd_sc_hd__mux2_1
X_29547_ net901 _01282_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[27\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_26759_ _11735_ net1706 _11737_ _11739_ VGND VGND VPWR VPWR _03309_ sky130_fd_sc_hd__a31o_1
X_14773_ _13312_ _13314_ VGND VGND VPWR VPWR _13326_ sky130_fd_sc_hd__nor2_2
X_19300_ _06595_ VGND VGND VPWR VPWR _06596_ sky130_fd_sc_hd__clkbuf_16
X_16512_ net2994 _14472_ _04489_ VGND VGND VPWR VPWR _04494_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29478_ net840 _01213_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[2\]\[17\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__10259_ clknet_0__10259_ VGND VGND VPWR VPWR clknet_1_1__leaf__10259_
+ sky130_fd_sc_hd__clkbuf_16
X_17492_ _05014_ VGND VGND VPWR VPWR _01296_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_112_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19231_ _06535_ _06536_ VGND VGND VPWR VPWR _06537_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_195_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16443_ _04456_ VGND VGND VPWR VPWR _01819_ sky130_fd_sc_hd__clkbuf_1
X_28429_ _12693_ VGND VGND VPWR VPWR _04025_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19162_ _06475_ _06471_ net38 VGND VGND VPWR VPWR _06477_ sky130_fd_sc_hd__or3_1
X_31440_ clknet_leaf_28_clk net1289 VGND VGND VPWR VPWR rvcpu.dp.plem.ResultSrcM\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_16374_ net2343 _14472_ _14547_ VGND VGND VPWR VPWR _14552_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_136_3755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_136_3766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18113_ _05475_ _05478_ VGND VGND VPWR VPWR _05480_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15325_ _13517_ _13563_ VGND VGND VPWR VPWR _13862_ sky130_fd_sc_hd__nand2_1
X_19093_ _06400_ _06403_ _06406_ _06409_ VGND VGND VPWR VPWR _06416_ sky130_fd_sc_hd__a211oi_2
X_31371_ clknet_leaf_18_clk _03074_ VGND VGND VPWR VPWR rvcpu.dp.plde.ImmExtE\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_23359__995 clknet_1_1__leaf__10138_ VGND VGND VPWR VPWR net1121 sky130_fd_sc_hd__inv_2
X_18044_ rvcpu.dp.plem.ALUResultM\[10\] _05413_ _05176_ VGND VGND VPWR VPWR _05414_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30322_ net668 _02057_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[4\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_15256_ _13284_ _13425_ VGND VGND VPWR VPWR _13796_ sky130_fd_sc_hd__nand2_2
XFILLER_0_48_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15187_ _13389_ _13353_ _13729_ _13412_ VGND VGND VPWR VPWR _13730_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_39_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30253_ net607 _01988_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[6\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__10081_ clknet_0__10081_ VGND VGND VPWR VPWR clknet_1_0__leaf__10081_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30184_ net538 _01919_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[8\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_19995_ datamem.data_ram\[18\]\[2\] _06930_ _06924_ datamem.data_ram\[23\]\[2\] VGND
+ VGND VPWR VPWR _07289_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18946_ _06174_ _06283_ _05698_ VGND VGND VPWR VPWR _06284_ sky130_fd_sc_hd__mux2_1
XFILLER_0_225_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_3_clk clknet_5_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_225_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18877_ _05520_ _05730_ _06108_ _05472_ VGND VGND VPWR VPWR _06220_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17828_ _13206_ rvcpu.dp.plde.RD2E\[23\] _05195_ VGND VGND VPWR VPWR _05213_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32825_ clknet_leaf_159_clk _04247_ VGND VGND VPWR VPWR datamem.data_ram\[12\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_222_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17759_ rvcpu.dp.plde.Rs2E\[1\] rvcpu.dp.plde.Rs2E\[0\] rvcpu.dp.plde.Rs2E\[2\] rvcpu.dp.plde.Rs2E\[4\]
+ VGND VGND VPWR VPWR _05157_ sky130_fd_sc_hd__or4_1
XFILLER_0_89_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20770_ datamem.data_ram\[60\]\[6\] datamem.data_ram\[61\]\[6\] _07829_ VGND VGND
+ VPWR VPWR _08060_ sky130_fd_sc_hd__mux2_1
X_32756_ clknet_leaf_162_clk _04178_ VGND VGND VPWR VPWR datamem.data_ram\[15\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_187_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31707_ clknet_leaf_31_clk _03165_ VGND VGND VPWR VPWR rvcpu.dp.pcreg.q\[25\] sky130_fd_sc_hd__dfxtp_1
X_19429_ _06668_ VGND VGND VPWR VPWR _06725_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_159_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32687_ clknet_leaf_86_clk _04109_ VGND VGND VPWR VPWR datamem.data_ram\[18\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22440_ rvcpu.dp.rf.reg_file_arr\[16\]\[7\] rvcpu.dp.rf.reg_file_arr\[17\]\[7\] rvcpu.dp.rf.reg_file_arr\[18\]\[7\]
+ rvcpu.dp.rf.reg_file_arr\[19\]\[7\] _09406_ _09408_ VGND VGND VPWR VPWR _09599_
+ sky130_fd_sc_hd__mux4_1
X_31638_ clknet_leaf_68_clk net1184 VGND VGND VPWR VPWR rvcpu.dp.plmw.lAuiPCW\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22371_ _09421_ VGND VGND VPWR VPWR _09534_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_31_1296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_212_5590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31569_ clknet_leaf_62_clk datamem.rd_data_mem\[19\] VGND VGND VPWR VPWR rvcpu.dp.plmw.ReadDataW\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21322_ _08580_ rvcpu.dp.plde.RdE\[0\] rvcpu.dp.plde.RdE\[1\] _08581_ _08583_ VGND
+ VGND VPWR VPWR _08584_ sky130_fd_sc_hd__a221o_1
X_25090_ _10776_ VGND VGND VPWR VPWR _02603_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_107_Left_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_384 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold420 datamem.data_ram\[30\]\[7\] VGND VGND VPWR VPWR net1570 sky130_fd_sc_hd__dlygate4sd3_1
X_21253_ _08514_ VGND VGND VPWR VPWR _08515_ sky130_fd_sc_hd__buf_2
Xhold431 rvcpu.dp.plem.ALUResultM\[1\] VGND VGND VPWR VPWR net1581 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold442 datamem.data_ram\[42\]\[6\] VGND VGND VPWR VPWR net1592 sky130_fd_sc_hd__dlygate4sd3_1
Xhold453 datamem.data_ram\[18\]\[5\] VGND VGND VPWR VPWR net1603 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_596 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20204_ datamem.data_ram\[63\]\[11\] _06761_ _07493_ _07496_ VGND VGND VPWR VPWR
+ _07497_ sky130_fd_sc_hd__o211a_1
XFILLER_0_229_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold464 datamem.data_ram\[31\]\[4\] VGND VGND VPWR VPWR net1614 sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 datamem.data_ram\[63\]\[5\] VGND VGND VPWR VPWR net1625 sky130_fd_sc_hd__dlygate4sd3_1
X_21184_ net118 _08470_ _08466_ VGND VGND VPWR VPWR _08471_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_25_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold486 datamem.data_ram\[10\]\[4\] VGND VGND VPWR VPWR net1636 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_221_5804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold497 datamem.data_ram\[26\]\[6\] VGND VGND VPWR VPWR net1647 sky130_fd_sc_hd__dlygate4sd3_1
X_27800_ _12136_ net4203 _12336_ VGND VGND VPWR VPWR _12342_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_229_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20135_ datamem.data_ram\[38\]\[27\] _06626_ _06820_ datamem.data_ram\[32\]\[27\]
+ VGND VGND VPWR VPWR _07428_ sky130_fd_sc_hd__o22a_1
X_28780_ _12891_ VGND VGND VPWR VPWR _04178_ sky130_fd_sc_hd__clkbuf_1
X_25992_ _08570_ _11315_ _11312_ _11320_ VGND VGND VPWR VPWR _02961_ sky130_fd_sc_hd__o211a_1
XFILLER_0_176_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27731_ _12304_ VGND VGND VPWR VPWR _03716_ sky130_fd_sc_hd__clkbuf_1
X_24943_ _10690_ VGND VGND VPWR VPWR _02542_ sky130_fd_sc_hd__clkbuf_1
X_20066_ datamem.data_ram\[50\]\[26\] _06608_ _06660_ datamem.data_ram\[53\]\[26\]
+ VGND VGND VPWR VPWR _07360_ sky130_fd_sc_hd__o22a_1
X_23580__202 clknet_1_0__leaf__10176_ VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__inv_2
Xhold1120 rvcpu.dp.rf.reg_file_arr\[25\]\[26\] VGND VGND VPWR VPWR net2270 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_137_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1131 datamem.data_ram\[25\]\[27\] VGND VGND VPWR VPWR net2281 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1142 datamem.data_ram\[45\]\[23\] VGND VGND VPWR VPWR net2292 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1153 datamem.data_ram\[47\]\[11\] VGND VGND VPWR VPWR net2303 sky130_fd_sc_hd__dlygate4sd3_1
X_27662_ _12267_ VGND VGND VPWR VPWR _03684_ sky130_fd_sc_hd__clkbuf_1
Xhold1164 rvcpu.dp.rf.reg_file_arr\[2\]\[11\] VGND VGND VPWR VPWR net2314 sky130_fd_sc_hd__dlygate4sd3_1
X_24874_ _10653_ VGND VGND VPWR VPWR _02510_ sky130_fd_sc_hd__clkbuf_1
Xhold1175 datamem.data_ram\[37\]\[22\] VGND VGND VPWR VPWR net2325 sky130_fd_sc_hd__dlygate4sd3_1
X_29401_ clknet_leaf_1_clk _01136_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD2E\[12\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_116_Left_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_79_Right_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26613_ _11654_ VGND VGND VPWR VPWR _03248_ sky130_fd_sc_hd__clkbuf_1
Xhold1186 rvcpu.dp.rf.reg_file_arr\[4\]\[20\] VGND VGND VPWR VPWR net2336 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_304 _14145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1197 rvcpu.dp.rf.reg_file_arr\[5\]\[25\] VGND VGND VPWR VPWR net2347 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_219_5744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27593_ _12230_ VGND VGND VPWR VPWR _03652_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_315 _14177_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_219_5755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_326 _14453_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29332_ clknet_leaf_145_clk _01067_ VGND VGND VPWR VPWR datamem.data_ram\[62\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_337 _14463_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26544_ _11089_ _11610_ VGND VGND VPWR VPWR _11616_ sky130_fd_sc_hd__and2_1
XANTENNA_348 datamem.data_ram\[52\]\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_359 rvcpu.dp.SrcBFW_Mux.y\[21\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20968_ _08255_ _08256_ _06606_ VGND VGND VPWR VPWR _08257_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_172_4612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_4623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22707_ _09850_ _09851_ _09449_ VGND VGND VPWR VPWR _09852_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_4634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29263_ _13152_ VGND VGND VPWR VPWR _04400_ sky130_fd_sc_hd__clkbuf_1
X_26475_ _11535_ rvcpu.ALUResultE\[30\] _11157_ VGND VGND VPWR VPWR _11595_ sky130_fd_sc_hd__a21o_1
XFILLER_0_166_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20899_ datamem.data_ram\[1\]\[22\] _06659_ _08188_ _07845_ VGND VGND VPWR VPWR _08189_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_82_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22985__692 clknet_1_1__leaf__10083_ VGND VGND VPWR VPWR net818 sky130_fd_sc_hd__inv_2
XFILLER_0_166_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28214_ _12359_ net3855 net45 VGND VGND VPWR VPWR _12576_ sky130_fd_sc_hd__mux2_1
XFILLER_0_192_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25426_ _10766_ net4069 _10961_ VGND VGND VPWR VPWR _10969_ sky130_fd_sc_hd__mux2_1
X_22638_ rvcpu.dp.rf.reg_file_arr\[0\]\[17\] rvcpu.dp.rf.reg_file_arr\[1\]\[17\] rvcpu.dp.rf.reg_file_arr\[2\]\[17\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[17\] _09714_ _09585_ VGND VGND VPWR VPWR _09787_
+ sky130_fd_sc_hd__mux4_1
X_29194_ _09309_ net4076 _13112_ VGND VGND VPWR VPWR _13115_ sky130_fd_sc_hd__mux2_1
X_25357_ _10876_ net1480 _10920_ _10927_ VGND VGND VPWR VPWR _02719_ sky130_fd_sc_hd__a31o_1
X_28145_ _12450_ net2815 net73 VGND VGND VPWR VPWR _12539_ sky130_fd_sc_hd__mux2_1
X_22569_ rvcpu.dp.rf.reg_file_arr\[12\]\[13\] rvcpu.dp.rf.reg_file_arr\[13\]\[13\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[13\] rvcpu.dp.rf.reg_file_arr\[15\]\[13\] _09552_
+ _09721_ VGND VGND VPWR VPWR _09722_ sky130_fd_sc_hd__mux4_1
XFILLER_0_51_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_125_Left_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15110_ _13298_ _13463_ _13654_ _13368_ VGND VGND VPWR VPWR _13655_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_75_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_88_Right_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24308_ _10329_ VGND VGND VPWR VPWR _02268_ sky130_fd_sc_hd__clkbuf_1
X_16090_ net1947 _13184_ _14385_ VGND VGND VPWR VPWR _14387_ sky130_fd_sc_hd__mux2_1
X_28076_ _12502_ VGND VGND VPWR VPWR _03863_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_146_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_3630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25288_ _10886_ VGND VGND VPWR VPWR _02691_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_224_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_3641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15041_ _13338_ _13585_ _13587_ _13385_ VGND VGND VPWR VPWR _13588_ sky130_fd_sc_hd__a31o_1
XFILLER_0_106_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27027_ _11827_ _11899_ VGND VGND VPWR VPWR _11902_ sky130_fd_sc_hd__and2_1
XFILLER_0_160_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24239_ _09276_ net3577 _10288_ VGND VGND VPWR VPWR _10291_ sky130_fd_sc_hd__mux2_1
XFILLER_0_224_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24099__607 clknet_1_1__leaf__10258_ VGND VGND VPWR VPWR net733 sky130_fd_sc_hd__inv_2
X_18800_ _06144_ _06145_ _06147_ VGND VGND VPWR VPWR _06148_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19780_ datamem.data_ram\[37\]\[9\] _06865_ _07073_ _07074_ VGND VGND VPWR VPWR _07075_
+ sky130_fd_sc_hd__o211a_1
X_28978_ _10075_ _12989_ VGND VGND VPWR VPWR _12998_ sky130_fd_sc_hd__and2_1
X_16992_ _04748_ VGND VGND VPWR VPWR _01546_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_196_Right_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_207_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18731_ _06081_ _06082_ VGND VGND VPWR VPWR _06083_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_129_3581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27929_ _12416_ VGND VGND VPWR VPWR _03802_ sky130_fd_sc_hd__clkbuf_1
X_15943_ _14307_ VGND VGND VPWR VPWR _02054_ sky130_fd_sc_hd__clkbuf_1
X_23743__334 clknet_1_1__leaf__10199_ VGND VGND VPWR VPWR net460 sky130_fd_sc_hd__inv_2
XFILLER_0_223_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_129_3592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26507__59 clknet_1_0__leaf__11602_ VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_134_Left_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_97_Right_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_222_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_216_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18662_ _05604_ _05424_ VGND VGND VPWR VPWR _06017_ sky130_fd_sc_hd__nor2_1
X_30940_ clknet_leaf_3_clk _02675_ VGND VGND VPWR VPWR datamem.data_ram\[40\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_69_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15874_ _14269_ VGND VGND VPWR VPWR _02085_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_203_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_125_3489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17613_ _13272_ net4109 _05068_ VGND VGND VPWR VPWR _05078_ sky130_fd_sc_hd__mux2_1
X_14825_ _13377_ VGND VGND VPWR VPWR _13378_ sky130_fd_sc_hd__buf_2
XFILLER_0_188_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30871_ clknet_leaf_62_clk _02606_ VGND VGND VPWR VPWR datamem.data_ram\[42\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_18593_ _05750_ _05937_ _05946_ _05951_ VGND VGND VPWR VPWR _05952_ sky130_fd_sc_hd__o211a_1
XFILLER_0_8_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23858__421 clknet_1_0__leaf__10219_ VGND VGND VPWR VPWR net547 sky130_fd_sc_hd__inv_2
XFILLER_0_59_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32610_ clknet_leaf_81_clk _04032_ VGND VGND VPWR VPWR datamem.data_ram\[20\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_17544_ _05041_ VGND VGND VPWR VPWR _01271_ sky130_fd_sc_hd__clkbuf_1
X_14756_ _13304_ _13308_ VGND VGND VPWR VPWR _13309_ sky130_fd_sc_hd__nor2_2
XFILLER_0_25_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32541_ clknet_leaf_78_clk _03963_ VGND VGND VPWR VPWR datamem.data_ram\[23\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17475_ _14189_ net4166 _04996_ VGND VGND VPWR VPWR _05005_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14687_ rvcpu.dp.plmw.ALUResultW\[9\] rvcpu.dp.plmw.ReadDataW\[9\] rvcpu.dp.plmw.PCPlus4W\[9\]
+ rvcpu.dp.plmw.lAuiPCW\[9\] _13168_ _13170_ VGND VGND VPWR VPWR _13250_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_28_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19214_ rvcpu.dp.plde.ImmExtE\[25\] rvcpu.dp.plde.PCE\[25\] VGND VGND VPWR VPWR _06522_
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_28_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16426_ _14579_ VGND VGND VPWR VPWR _01827_ sky130_fd_sc_hd__clkbuf_1
X_32472_ clknet_leaf_4_clk _03894_ VGND VGND VPWR VPWR datamem.data_ram\[26\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_60_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_143_Left_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19145_ _06461_ rvcpu.dp.plde.ImmExtE\[16\] _06419_ VGND VGND VPWR VPWR _06462_ sky130_fd_sc_hd__mux2_1
X_31423_ clknet_leaf_59_clk _03126_ VGND VGND VPWR VPWR datamem.data_ram\[44\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16357_ net2518 _14455_ _14536_ VGND VGND VPWR VPWR _14543_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15308_ _13499_ _13830_ _13835_ _13845_ _13638_ VGND VGND VPWR VPWR _13846_ sky130_fd_sc_hd__o32a_1
XFILLER_0_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19076_ rvcpu.dp.plde.ImmExtE\[8\] rvcpu.dp.plde.PCE\[8\] VGND VGND VPWR VPWR _06401_
+ sky130_fd_sc_hd__nand2_1
X_31354_ clknet_leaf_17_clk _03057_ VGND VGND VPWR VPWR rvcpu.dp.plde.ImmExtE\[3\]
+ sky130_fd_sc_hd__dfxtp_2
Xclkbuf_1_0__f__10202_ clknet_0__10202_ VGND VGND VPWR VPWR clknet_1_0__leaf__10202_
+ sky130_fd_sc_hd__clkbuf_16
X_16288_ _14506_ VGND VGND VPWR VPWR _01892_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_1094 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18027_ _05389_ _05395_ _05396_ VGND VGND VPWR VPWR _05397_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30305_ net651 _02040_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[5\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_15239_ _13419_ _13323_ _13750_ VGND VGND VPWR VPWR _13779_ sky130_fd_sc_hd__or3_1
XFILLER_0_140_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31285_ clknet_leaf_110_clk _02988_ VGND VGND VPWR VPWR datamem.data_ram\[34\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__10133_ clknet_0__10133_ VGND VGND VPWR VPWR clknet_1_0__leaf__10133_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_140_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_199_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30236_ net590 _01971_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[7\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_1270 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_58_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19978_ datamem.data_ram\[19\]\[18\] _06634_ _07271_ _06679_ VGND VGND VPWR VPWR
+ _07272_ sky130_fd_sc_hd__o211a_1
X_30167_ net529 _01902_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[0\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_152_Left_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_163_Right_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18929_ _05531_ _05537_ _06251_ VGND VGND VPWR VPWR _06268_ sky130_fd_sc_hd__or3_1
XFILLER_0_226_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30098_ net460 _01833_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[11\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_21940_ _08682_ _09170_ _09172_ _08575_ VGND VGND VPWR VPWR _09173_ sky130_fd_sc_hd__o211a_1
X_21871_ _08547_ _09105_ _09107_ _08576_ VGND VGND VPWR VPWR _09108_ sky130_fd_sc_hd__o211a_1
XFILLER_0_171_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32808_ clknet_leaf_190_clk _04230_ VGND VGND VPWR VPWR datamem.data_ram\[13\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_20822_ datamem.data_ram\[30\]\[30\] _07860_ _07863_ datamem.data_ram\[28\]\[30\]
+ VGND VGND VPWR VPWR _08112_ sky130_fd_sc_hd__o22a_1
XFILLER_0_210_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24590_ _10394_ net3869 _10491_ VGND VGND VPWR VPWR _10496_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20753_ datamem.data_ram\[15\]\[6\] _07833_ _08042_ _06623_ VGND VGND VPWR VPWR _08043_
+ sky130_fd_sc_hd__o211a_1
X_32739_ clknet_leaf_252_clk _04161_ VGND VGND VPWR VPWR datamem.data_ram\[16\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_214_5630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_214_5641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_611 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26260_ net1371 _11432_ VGND VGND VPWR VPWR _11462_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_161_Left_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20684_ datamem.data_ram\[34\]\[5\] _07136_ _07971_ _07974_ VGND VGND VPWR VPWR _07975_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_119_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_210_5527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25211_ _10844_ VGND VGND VPWR VPWR _02656_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_210_5538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22423_ _09451_ _09580_ _09582_ _09523_ VGND VGND VPWR VPWR _09583_ sky130_fd_sc_hd__o211a_1
X_26191_ rvcpu.ALUControl\[1\] _11432_ VGND VGND VPWR VPWR _11433_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25142_ _10803_ VGND VGND VPWR VPWR _02628_ sky130_fd_sc_hd__clkbuf_1
X_23690__285 clknet_1_1__leaf__10195_ VGND VGND VPWR VPWR net411 sky130_fd_sc_hd__inv_2
X_22354_ _08592_ VGND VGND VPWR VPWR _09517_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_143_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21305_ _08566_ VGND VGND VPWR VPWR _08567_ sky130_fd_sc_hd__buf_8
X_25073_ _10767_ VGND VGND VPWR VPWR _02595_ sky130_fd_sc_hd__clkbuf_1
X_29950_ net320 _01685_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[15\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22285_ _09444_ _09448_ _09449_ VGND VGND VPWR VPWR _09450_ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28901_ _12955_ VGND VGND VPWR VPWR _04235_ sky130_fd_sc_hd__clkbuf_1
Xhold250 datamem.data_ram\[57\]\[6\] VGND VGND VPWR VPWR net1400 sky130_fd_sc_hd__dlygate4sd3_1
X_21236_ datamem.data_ram\[52\]\[12\] datamem.data_ram\[53\]\[12\] VGND VGND VPWR
+ VPWR _08499_ sky130_fd_sc_hd__nand2_2
Xhold261 datamem.data_ram\[39\]\[5\] VGND VGND VPWR VPWR net1411 sky130_fd_sc_hd__dlygate4sd3_1
X_29881_ net259 _01616_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[17\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_208_5478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold272 datamem.data_ram\[28\]\[0\] VGND VGND VPWR VPWR net1422 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_208_5489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold283 datamem.data_ram\[20\]\[1\] VGND VGND VPWR VPWR net1433 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_165_4460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold294 datamem.data_ram\[20\]\[7\] VGND VGND VPWR VPWR net1444 sky130_fd_sc_hd__dlygate4sd3_1
X_28832_ _12760_ net2282 _12914_ VGND VGND VPWR VPWR _12919_ sky130_fd_sc_hd__mux2_1
X_21167_ _08454_ _08455_ _07819_ VGND VGND VPWR VPWR _08456_ sky130_fd_sc_hd__mux2_1
XFILLER_0_217_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20118_ _06715_ _07395_ _07400_ _06860_ _07411_ VGND VGND VPWR VPWR _07412_ sky130_fd_sc_hd__o311a_1
XFILLER_0_176_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_161_4357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_130_Right_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28763_ _12696_ net2980 _12877_ VGND VGND VPWR VPWR _12882_ sky130_fd_sc_hd__mux2_1
X_21098_ datamem.data_ram\[12\]\[7\] datamem.data_ram\[13\]\[7\] _07874_ VGND VGND
+ VPWR VPWR _08387_ sky130_fd_sc_hd__mux2_1
X_25975_ net1785 _11302_ _11300_ _11310_ VGND VGND VPWR VPWR _02954_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_161_4368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27714_ _12295_ VGND VGND VPWR VPWR _03708_ sky130_fd_sc_hd__clkbuf_1
X_20049_ datamem.data_ram\[15\]\[26\] _06760_ _07339_ _07342_ VGND VGND VPWR VPWR
+ _07343_ sky130_fd_sc_hd__o211a_1
X_24926_ _10681_ VGND VGND VPWR VPWR _02534_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_176_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28694_ _12845_ VGND VGND VPWR VPWR _04138_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_176_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_198_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27645_ _12138_ net2737 _12251_ VGND VGND VPWR VPWR _12258_ sky130_fd_sc_hd__mux2_1
XFILLER_0_213_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24857_ _10644_ VGND VGND VPWR VPWR _02502_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_101 _06917_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_112 _07077_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_198_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_123 _07367_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14610_ _13191_ VGND VGND VPWR VPWR _03200_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_64_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_134 _07831_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27576_ _12221_ VGND VGND VPWR VPWR _03644_ sky130_fd_sc_hd__clkbuf_1
X_15590_ _14102_ VGND VGND VPWR VPWR _02210_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_120_3364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24788_ _10606_ VGND VGND VPWR VPWR _02471_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_145 _07840_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_156 _08408_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_3386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29315_ clknet_leaf_290_clk _01050_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD1E\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_167 _08693_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26527_ _10783_ _11604_ _11605_ net1552 VGND VGND VPWR VPWR _03211_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_178 _08937_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_189 _09226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0__10127_ _10127_ VGND VGND VPWR VPWR clknet_0__10127_ sky130_fd_sc_hd__clkbuf_16
X_29246_ _13143_ VGND VGND VPWR VPWR _04392_ sky130_fd_sc_hd__clkbuf_1
X_17260_ _14179_ net4209 _04887_ VGND VGND VPWR VPWR _04891_ sky130_fd_sc_hd__mux2_1
X_26458_ _11576_ _11223_ _11540_ _06518_ _11583_ VGND VGND VPWR VPWR _11584_ sky130_fd_sc_hd__a221o_1
XFILLER_0_3_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23241__889 clknet_1_0__leaf__10126_ VGND VGND VPWR VPWR net1015 sky130_fd_sc_hd__inv_2
X_16211_ _13237_ VGND VGND VPWR VPWR _14459_ sky130_fd_sc_hd__buf_4
X_25409_ _10954_ net1560 _10949_ _10959_ VGND VGND VPWR VPWR _02739_ sky130_fd_sc_hd__a31o_1
XFILLER_0_153_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29177_ _09239_ net2702 net63 VGND VGND VPWR VPWR _13106_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_23_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17191_ _04854_ VGND VGND VPWR VPWR _01445_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26389_ _13387_ _11329_ _11532_ _11534_ VGND VGND VPWR VPWR _03144_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_23_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload109 clknet_leaf_59_clk VGND VGND VPWR VPWR clkload109/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_148_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28128_ _12433_ net3156 _12528_ VGND VGND VPWR VPWR _12530_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16142_ net2289 _13263_ _14407_ VGND VGND VPWR VPWR _14414_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28059_ _12493_ VGND VGND VPWR VPWR _03855_ sky130_fd_sc_hd__clkbuf_1
X_16073_ _14377_ VGND VGND VPWR VPWR _01986_ sky130_fd_sc_hd__clkbuf_1
X_23587__208 clknet_1_0__leaf__10177_ VGND VGND VPWR VPWR net334 sky130_fd_sc_hd__inv_2
X_15024_ _13535_ _13540_ _13544_ _13571_ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__o31a_1
X_19901_ datamem.data_ram\[0\]\[17\] _07191_ _07192_ _07195_ VGND VGND VPWR VPWR _07196_
+ sky130_fd_sc_hd__o211a_1
X_31070_ clknet_leaf_158_clk _02805_ VGND VGND VPWR VPWR datamem.data_ram\[9\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_19832_ _06952_ VGND VGND VPWR VPWR _07127_ sky130_fd_sc_hd__buf_4
X_30021_ net383 _01756_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[13\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_53_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19763_ _06752_ _07052_ _07057_ VGND VGND VPWR VPWR _07058_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_53_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16975_ _04739_ VGND VGND VPWR VPWR _01554_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_208_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18714_ _05702_ _06059_ _06066_ VGND VGND VPWR VPWR _06067_ sky130_fd_sc_hd__a21o_1
X_15926_ net2103 _13248_ _14297_ VGND VGND VPWR VPWR _14299_ sky130_fd_sc_hd__mux2_1
X_19694_ _06937_ VGND VGND VPWR VPWR _06990_ sky130_fd_sc_hd__clkbuf_8
X_31972_ clknet_leaf_130_clk _03394_ VGND VGND VPWR VPWR datamem.data_ram\[54\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_204_631 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18645_ _05692_ _05764_ VGND VGND VPWR VPWR _06001_ sky130_fd_sc_hd__or2_1
X_30923_ clknet_leaf_192_clk _02658_ VGND VGND VPWR VPWR datamem.data_ram\[40\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_15857_ net2887 _13251_ _14258_ VGND VGND VPWR VPWR _14261_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_203_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_204_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14808_ _13357_ _13360_ VGND VGND VPWR VPWR _13361_ sky130_fd_sc_hd__nor2_1
X_30854_ clknet_leaf_155_clk _02589_ VGND VGND VPWR VPWR datamem.data_ram\[43\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_18576_ _05676_ _05828_ VGND VGND VPWR VPWR _05935_ sky130_fd_sc_hd__or2_1
X_15788_ _14177_ net3191 _14221_ VGND VGND VPWR VPWR _14224_ sky130_fd_sc_hd__mux2_1
X_24153__656 clknet_1_0__leaf__10263_ VGND VGND VPWR VPWR net782 sky130_fd_sc_hd__inv_2
X_17527_ _13244_ net2447 _05032_ VGND VGND VPWR VPWR _05033_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14739_ _13291_ VGND VGND VPWR VPWR _13292_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_15_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30785_ clknet_leaf_191_clk _02520_ VGND VGND VPWR VPWR datamem.data_ram\[46\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32524_ clknet_leaf_253_clk _03946_ VGND VGND VPWR VPWR datamem.data_ram\[24\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17458_ _04973_ VGND VGND VPWR VPWR _04996_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_15_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16409_ _14570_ VGND VGND VPWR VPWR _01835_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32455_ clknet_leaf_274_clk _03877_ VGND VGND VPWR VPWR datamem.data_ram\[27\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_23300__942 clknet_1_1__leaf__10132_ VGND VGND VPWR VPWR net1068 sky130_fd_sc_hd__inv_2
X_17389_ _04959_ VGND VGND VPWR VPWR _01344_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_1346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19128_ _06445_ _06446_ VGND VGND VPWR VPWR _06447_ sky130_fd_sc_hd__and2_1
X_31406_ clknet_leaf_30_clk _03109_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCE\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32386_ clknet_leaf_238_clk _03808_ VGND VGND VPWR VPWR datamem.data_ram\[29\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19059_ rvcpu.dp.plde.ImmExtE\[6\] rvcpu.dp.plde.PCE\[6\] VGND VGND VPWR VPWR _06386_
+ sky130_fd_sc_hd__nand2_1
X_31337_ clknet_leaf_14_clk _03040_ VGND VGND VPWR VPWR rvcpu.dp.plde.Rs2E\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22070_ _09286_ VGND VGND VPWR VPWR _01073_ sky130_fd_sc_hd__clkbuf_1
X_31268_ clknet_leaf_35_clk _02971_ VGND VGND VPWR VPWR rvcpu.dp.plfd.InstrD\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21021_ datamem.data_ram\[54\]\[31\] _06626_ _06685_ datamem.data_ram\[52\]\[31\]
+ _08309_ VGND VGND VPWR VPWR _08310_ sky130_fd_sc_hd__o221a_1
X_30219_ net573 _01954_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[7\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31199_ clknet_leaf_43_clk _02902_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCPlus4D\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_227_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_226_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_203_5364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_203_5375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_226_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25760_ net1623 _11144_ _11147_ _11161_ VGND VGND VPWR VPWR _02888_ sky130_fd_sc_hd__o211a_1
XFILLER_0_198_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_491 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24711_ _10563_ VGND VGND VPWR VPWR _02437_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_223_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21923_ rvcpu.dp.rf.reg_file_arr\[12\]\[28\] rvcpu.dp.rf.reg_file_arr\[13\]\[28\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[28\] rvcpu.dp.rf.reg_file_arr\[15\]\[28\] _08549_
+ _08553_ VGND VGND VPWR VPWR _09157_ sky130_fd_sc_hd__mux4_1
X_25691_ _11105_ net1744 _11111_ _11117_ VGND VGND VPWR VPWR _02863_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_195_5165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_195_5176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_210_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_195_5187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27430_ _12138_ net1958 _12126_ VGND VGND VPWR VPWR _12139_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21854_ _09083_ _09087_ _09091_ _08624_ VGND VGND VPWR VPWR _01052_ sky130_fd_sc_hd__o31a_1
X_24642_ _10392_ net3207 _10521_ VGND VGND VPWR VPWR _10525_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_210_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20805_ _08084_ _08088_ _06681_ _08094_ VGND VGND VPWR VPWR _08095_ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_195_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_194_335 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27361_ _12083_ net4098 _12097_ VGND VGND VPWR VPWR _12099_ sky130_fd_sc_hd__mux2_1
X_24573_ _10448_ net3391 _10482_ VGND VGND VPWR VPWR _10487_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21785_ _08725_ _09025_ VGND VGND VPWR VPWR _09026_ sky130_fd_sc_hd__nor2_1
XFILLER_0_203_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29100_ _09325_ net2680 _13058_ VGND VGND VPWR VPWR _13065_ sky130_fd_sc_hd__mux2_1
X_26312_ net1819 _11436_ VGND VGND VPWR VPWR _11489_ sky130_fd_sc_hd__and2_1
Xclkbuf_5_20__f_clk clknet_2_2_0_clk VGND VGND VPWR VPWR clknet_5_20__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_20736_ datamem.data_ram\[36\]\[6\] datamem.data_ram\[37\]\[6\] _07828_ VGND VGND
+ VPWR VPWR _08026_ sky130_fd_sc_hd__mux2_1
X_23524_ _10170_ VGND VGND VPWR VPWR _01643_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27292_ _11946_ _12054_ VGND VGND VPWR VPWR _12059_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_154_4183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23772__360 clknet_1_0__leaf__10202_ VGND VGND VPWR VPWR net486 sky130_fd_sc_hd__inv_2
X_29031_ _13027_ VGND VGND VPWR VPWR _04293_ sky130_fd_sc_hd__clkbuf_1
X_26243_ _11439_ VGND VGND VPWR VPWR _11459_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_154_4194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23455_ clknet_1_0__leaf__10152_ VGND VGND VPWR VPWR _10157_ sky130_fd_sc_hd__buf_1
X_20667_ datamem.data_ram\[51\]\[29\] _06729_ _06684_ datamem.data_ram\[52\]\[29\]
+ VGND VGND VPWR VPWR _07958_ sky130_fd_sc_hd__o22a_1
XFILLER_0_92_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22406_ rvcpu.dp.rf.reg_file_arr\[4\]\[5\] rvcpu.dp.rf.reg_file_arr\[5\]\[5\] rvcpu.dp.rf.reg_file_arr\[6\]\[5\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[5\] _09464_ _09467_ VGND VGND VPWR VPWR _09567_ sky130_fd_sc_hd__mux4_1
XFILLER_0_190_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26174_ _09457_ _11362_ VGND VGND VPWR VPWR _11424_ sky130_fd_sc_hd__and2_1
X_23386_ _09298_ net3725 _10143_ VGND VGND VPWR VPWR _10144_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20598_ _07839_ _07886_ _07888_ _07868_ VGND VGND VPWR VPWR _07889_ sky130_fd_sc_hd__a211o_1
XFILLER_0_116_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_167_4500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_285_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_285_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_167_4511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25125_ _10794_ VGND VGND VPWR VPWR _02620_ sky130_fd_sc_hd__clkbuf_1
X_22337_ _09441_ _09500_ VGND VGND VPWR VPWR _09501_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25056_ _09239_ VGND VGND VPWR VPWR _10756_ sky130_fd_sc_hd__buf_2
X_29933_ net303 _01668_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[16\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_22268_ _09392_ VGND VGND VPWR VPWR _09434_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_163_4408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_4419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21219_ _08487_ _08464_ _08490_ VGND VGND VPWR VPWR _04430_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_104_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29864_ net242 _01599_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[18\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22199_ _09372_ VGND VGND VPWR VPWR _01116_ sky130_fd_sc_hd__clkbuf_1
X_28815_ _12696_ net3779 _12905_ VGND VGND VPWR VPWR _12910_ sky130_fd_sc_hd__mux2_1
XFILLER_0_218_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29795_ net1141 _01530_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[20\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16760_ net3413 _14447_ _04623_ VGND VGND VPWR VPWR _04626_ sky130_fd_sc_hd__mux2_1
X_28746_ _12743_ net3822 net41 VGND VGND VPWR VPWR _12873_ sky130_fd_sc_hd__mux2_1
X_25958_ net13 _11290_ _11300_ _11301_ VGND VGND VPWR VPWR _02946_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_122_3415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_3426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15711_ _14178_ VGND VGND VPWR VPWR _02165_ sky130_fd_sc_hd__clkbuf_1
X_24909_ _10672_ VGND VGND VPWR VPWR _02526_ sky130_fd_sc_hd__clkbuf_1
X_28677_ _12836_ VGND VGND VPWR VPWR _04130_ sky130_fd_sc_hd__clkbuf_1
X_16691_ _04589_ VGND VGND VPWR VPWR _01696_ sky130_fd_sc_hd__clkbuf_1
X_25889_ net1284 _11143_ VGND VGND VPWR VPWR _11262_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_87_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18430_ _05750_ _05765_ _05777_ _05793_ VGND VGND VPWR VPWR _05794_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_158_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15642_ _14127_ net4340 _14131_ VGND VGND VPWR VPWR _14132_ sky130_fd_sc_hd__mux2_1
X_27628_ _12093_ net1899 _12242_ VGND VGND VPWR VPWR _12249_ sky130_fd_sc_hd__mux2_1
X_26497__50 clknet_1_0__leaf__11601_ VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__inv_2
XFILLER_0_158_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_83_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18361_ _05725_ VGND VGND VPWR VPWR _05726_ sky130_fd_sc_hd__buf_2
XFILLER_0_69_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_83_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15573_ net1886 _13184_ _14092_ VGND VGND VPWR VPWR _14094_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_83_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27559_ _12212_ VGND VGND VPWR VPWR _03636_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17312_ net4335 _13228_ _04913_ VGND VGND VPWR VPWR _04919_ sky130_fd_sc_hd__mux2_1
XFILLER_0_189_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30570_ clknet_leaf_138_clk _02305_ VGND VGND VPWR VPWR datamem.data_ram\[54\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_18292_ _05284_ _05290_ _05647_ _05655_ _05656_ VGND VGND VPWR VPWR _05657_ sky130_fd_sc_hd__a311o_1
X_17243_ _14162_ net3734 _04876_ VGND VGND VPWR VPWR _04882_ sky130_fd_sc_hd__mux2_1
X_29229_ _13134_ VGND VGND VPWR VPWR _04384_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_96_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32240_ clknet_leaf_278_clk _03662_ VGND VGND VPWR VPWR datamem.data_ram\[35\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_17174_ _04845_ VGND VGND VPWR VPWR _01453_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_226_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16125_ net2105 _13238_ _14396_ VGND VGND VPWR VPWR _14405_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_276_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_276_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32171_ clknet_leaf_210_clk _03593_ VGND VGND VPWR VPWR datamem.data_ram\[37\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31122_ clknet_leaf_110_clk _02857_ VGND VGND VPWR VPWR datamem.data_ram\[35\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_55_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16056_ _14368_ VGND VGND VPWR VPWR _01994_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_55_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15007_ _13333_ _13326_ _13337_ _13554_ rvcpu.dp.pcreg.q\[9\] VGND VGND VPWR VPWR
+ _13555_ sky130_fd_sc_hd__a311o_1
XFILLER_0_161_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31053_ clknet_leaf_114_clk _02788_ VGND VGND VPWR VPWR datamem.data_ram\[38\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_196_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2409 rvcpu.dp.rf.reg_file_arr\[9\]\[17\] VGND VGND VPWR VPWR net3559 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30004_ net374 _01739_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[14\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_19815_ datamem.data_ram\[16\]\[9\] _06697_ _06700_ datamem.data_ram\[17\]\[9\] _07109_
+ VGND VGND VPWR VPWR _07110_ sky130_fd_sc_hd__o221a_1
XFILLER_0_47_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1708 datamem.data_ram\[56\]\[8\] VGND VGND VPWR VPWR net2858 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1719 rvcpu.dp.rf.reg_file_arr\[3\]\[3\] VGND VGND VPWR VPWR net2869 sky130_fd_sc_hd__dlygate4sd3_1
X_23942__496 clknet_1_0__leaf__10228_ VGND VGND VPWR VPWR net622 sky130_fd_sc_hd__inv_2
X_19746_ datamem.data_ram\[34\]\[25\] _07023_ _07036_ _07040_ VGND VGND VPWR VPWR
+ _07041_ sky130_fd_sc_hd__o211a_1
X_16958_ _04730_ VGND VGND VPWR VPWR _01562_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_224_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_205_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15909_ net2145 _13223_ _14286_ VGND VGND VPWR VPWR _14290_ sky130_fd_sc_hd__mux2_1
X_19677_ _06936_ VGND VGND VPWR VPWR _06973_ sky130_fd_sc_hd__buf_6
X_31955_ clknet_leaf_118_clk _03377_ VGND VGND VPWR VPWR datamem.data_ram\[55\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16889_ net2146 _14440_ _04684_ VGND VGND VPWR VPWR _04694_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_200_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_200_clk
+ sky130_fd_sc_hd__clkbuf_8
X_18628_ _05706_ _05897_ _05984_ _05720_ VGND VGND VPWR VPWR _05985_ sky130_fd_sc_hd__a211o_1
X_30906_ clknet_leaf_216_clk _02641_ VGND VGND VPWR VPWR datamem.data_ram\[41\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31886_ clknet_leaf_112_clk _03340_ VGND VGND VPWR VPWR datamem.data_ram\[57\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23183__854 clknet_1_1__leaf__10111_ VGND VGND VPWR VPWR net980 sky130_fd_sc_hd__inv_2
XFILLER_0_63_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18559_ _05368_ _05726_ _05821_ _05918_ VGND VGND VPWR VPWR _05919_ sky130_fd_sc_hd__a211oi_1
X_30837_ clknet_leaf_263_clk _02572_ VGND VGND VPWR VPWR datamem.data_ram\[44\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_190_5051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_190_5062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21570_ _08672_ _08809_ _08816_ _08822_ VGND VGND VPWR VPWR _08823_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_16_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30768_ clknet_leaf_259_clk _02503_ VGND VGND VPWR VPWR datamem.data_ram\[47\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_12 _06608_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20521_ datamem.data_ram\[26\]\[21\] _07203_ _06604_ _07811_ VGND VGND VPWR VPWR
+ _07812_ sky130_fd_sc_hd__o211a_1
XANTENNA_23 _06620_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32507_ clknet_leaf_240_clk _03929_ VGND VGND VPWR VPWR datamem.data_ram\[24\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_34 _06661_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30699_ clknet_leaf_139_clk _02434_ VGND VGND VPWR VPWR datamem.data_ram\[4\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_45 _06678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_56 _06704_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_67 _06766_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20452_ datamem.data_ram\[14\]\[20\] _06744_ _06765_ datamem.data_ram\[12\]\[20\]
+ VGND VGND VPWR VPWR _07744_ sky130_fd_sc_hd__o22a_1
XANTENNA_78 _06777_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32438_ clknet_leaf_245_clk _03860_ VGND VGND VPWR VPWR datamem.data_ram\[27\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_89 _06797_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23984__519 clknet_1_0__leaf__10239_ VGND VGND VPWR VPWR net645 sky130_fd_sc_hd__inv_2
XFILLER_0_162_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23535__162 clknet_1_0__leaf__10171_ VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_267_clk clknet_5_19__leaf_clk VGND VGND VPWR VPWR clknet_leaf_267_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_127_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32369_ clknet_leaf_263_clk _03791_ VGND VGND VPWR VPWR datamem.data_ram\[2\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_20383_ datamem.data_ram\[53\]\[28\] _06721_ _07242_ datamem.data_ram\[49\]\[28\]
+ VGND VGND VPWR VPWR _07675_ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22122_ rvcpu.dp.plem.WriteDataM\[31\] _09221_ _09295_ rvcpu.dp.plem.WriteDataM\[15\]
+ _09328_ VGND VGND VPWR VPWR _09329_ sky130_fd_sc_hd__a221o_4
XFILLER_0_203_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_1268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_205_5404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_205_5415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_205_5426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26930_ _11827_ _11842_ VGND VGND VPWR VPWR _11845_ sky130_fd_sc_hd__and2_1
X_22053_ _09273_ net2585 _09270_ VGND VGND VPWR VPWR _09274_ sky130_fd_sc_hd__mux2_1
XFILLER_0_203_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_195_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21004_ datamem.data_ram\[19\]\[15\] _07911_ _08292_ _06928_ VGND VGND VPWR VPWR
+ _08293_ sky130_fd_sc_hd__a211o_1
Xhold2910 datamem.data_ram\[14\]\[22\] VGND VGND VPWR VPWR net4060 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26861_ _11795_ net1481 _11797_ _11800_ VGND VGND VPWR VPWR _03350_ sky130_fd_sc_hd__a31o_1
Xhold2921 rvcpu.dp.rf.reg_file_arr\[14\]\[30\] VGND VGND VPWR VPWR net4071 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2932 rvcpu.dp.rf.reg_file_arr\[0\]\[30\] VGND VGND VPWR VPWR net4082 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_197_5216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2943 datamem.data_ram\[7\]\[24\] VGND VGND VPWR VPWR net4093 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_197_5227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2954 datamem.data_ram\[8\]\[21\] VGND VGND VPWR VPWR net4104 sky130_fd_sc_hd__dlygate4sd3_1
X_28600_ _06591_ VGND VGND VPWR VPWR _12795_ sky130_fd_sc_hd__buf_8
X_25812_ rvcpu.dp.pcreg.q\[19\] _11197_ VGND VGND VPWR VPWR _11201_ sky130_fd_sc_hd__nor2_1
X_24021__553 clknet_1_0__leaf__10242_ VGND VGND VPWR VPWR net679 sky130_fd_sc_hd__inv_2
XFILLER_0_227_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2965 datamem.data_ram\[39\]\[10\] VGND VGND VPWR VPWR net4115 sky130_fd_sc_hd__dlygate4sd3_1
X_29580_ net934 _01315_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[26\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_26792_ _11753_ net1613 _11748_ _11758_ VGND VGND VPWR VPWR _03323_ sky130_fd_sc_hd__a31o_1
Xhold2976 datamem.data_ram\[12\]\[27\] VGND VGND VPWR VPWR net4126 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2987 rvcpu.dp.rf.reg_file_arr\[31\]\[24\] VGND VGND VPWR VPWR net4137 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2998 datamem.data_ram\[63\]\[12\] VGND VGND VPWR VPWR net4148 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28531_ _09239_ VGND VGND VPWR VPWR _12756_ sky130_fd_sc_hd__buf_2
X_25743_ net1597 _11144_ _11147_ _11148_ VGND VGND VPWR VPWR _02884_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_3_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22955_ clknet_1_0__leaf__10080_ VGND VGND VPWR VPWR _10081_ sky130_fd_sc_hd__buf_1
XFILLER_0_138_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_179_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21906_ _08541_ _09140_ VGND VGND VPWR VPWR _09141_ sky130_fd_sc_hd__and2_1
X_28462_ _09350_ _12622_ _12668_ VGND VGND VPWR VPWR _12713_ sky130_fd_sc_hd__a21oi_4
X_25674_ _11105_ net3985 _11097_ _11106_ VGND VGND VPWR VPWR _02857_ sky130_fd_sc_hd__a31o_1
Xmax_cap69 _12923_ VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__buf_4
X_22886_ _09388_ _10013_ _10017_ _10021_ VGND VGND VPWR VPWR _10022_ sky130_fd_sc_hd__and4_1
XFILLER_0_214_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_195_633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23307__948 clknet_1_0__leaf__10133_ VGND VGND VPWR VPWR net1074 sky130_fd_sc_hd__inv_2
XFILLER_0_167_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_4234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27413_ _12127_ VGND VGND VPWR VPWR _03575_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_214_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24625_ _10515_ VGND VGND VPWR VPWR _02399_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_214_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_156_4245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28393_ _12437_ net3075 _12669_ VGND VGND VPWR VPWR _12673_ sky130_fd_sc_hd__mux2_1
X_21837_ _08515_ _09074_ VGND VGND VPWR VPWR _09075_ sky130_fd_sc_hd__nor2_1
XFILLER_0_195_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_183_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27344_ _12087_ net3201 _12081_ VGND VGND VPWR VPWR _12088_ sky130_fd_sc_hd__mux2_1
X_23696__291 clknet_1_0__leaf__10195_ VGND VGND VPWR VPWR net417 sky130_fd_sc_hd__inv_2
X_24556_ _10476_ net3640 net60 VGND VGND VPWR VPWR _10477_ sky130_fd_sc_hd__mux2_1
X_21768_ _08742_ _09009_ VGND VGND VPWR VPWR _09010_ sky130_fd_sc_hd__or2_1
XFILLER_0_194_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20719_ _06988_ _07998_ _08009_ VGND VGND VPWR VPWR _08010_ sky130_fd_sc_hd__and3_1
XFILLER_0_53_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27275_ _10822_ net3268 _12043_ VGND VGND VPWR VPWR _12049_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21699_ rvcpu.dp.rf.reg_file_arr\[8\]\[16\] rvcpu.dp.rf.reg_file_arr\[10\]\[16\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[16\] rvcpu.dp.rf.reg_file_arr\[11\]\[16\] _08560_
+ _08561_ VGND VGND VPWR VPWR _08945_ sky130_fd_sc_hd__mux4_1
X_24487_ _09314_ datamem.data_ram\[52\]\[27\] _10430_ VGND VGND VPWR VPWR _10434_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29014_ _06587_ VGND VGND VPWR VPWR _13018_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_184_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_190_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26226_ net4349 _11361_ VGND VGND VPWR VPWR _11451_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_115_3252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_258_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_258_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_34_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_180_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26157_ _11415_ VGND VGND VPWR VPWR _03031_ sky130_fd_sc_hd__clkbuf_1
X_23369_ clknet_1_1__leaf__10130_ VGND VGND VPWR VPWR _10139_ sky130_fd_sc_hd__buf_1
XFILLER_0_1_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_186_4953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_186_4964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25108_ _10785_ VGND VGND VPWR VPWR _02612_ sky130_fd_sc_hd__clkbuf_1
X_26088_ _11378_ VGND VGND VPWR VPWR _11379_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_81_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17930_ _05300_ _05301_ VGND VGND VPWR VPWR _05303_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29916_ net286 _01651_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[16\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_25039_ _10472_ net2382 net90 VGND VGND VPWR VPWR _10746_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_992 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17861_ rvcpu.dp.plem.ALUResultM\[5\] _05176_ _05234_ _05235_ VGND VGND VPWR VPWR
+ rvcpu.dp.SrcBFW_Mux.y\[5\] sky130_fd_sc_hd__o22a_1
X_29847_ net225 _01582_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[18\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_89_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16812_ _04653_ VGND VGND VPWR VPWR _01631_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_89_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19600_ datamem.data_ram\[51\]\[8\] _06634_ _06892_ _06895_ VGND VGND VPWR VPWR _06896_
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_145_3971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17792_ _05187_ VGND VGND VPWR VPWR rvcpu.dp.SrcBFW_Mux.y\[2\] sky130_fd_sc_hd__buf_1
X_29778_ net1124 _01513_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[20\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_145_3982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19531_ datamem.data_ram\[41\]\[24\] _06790_ _06822_ _06826_ VGND VGND VPWR VPWR
+ _06827_ sky130_fd_sc_hd__o211a_1
X_28729_ _12760_ net3534 _12859_ VGND VGND VPWR VPWR _12864_ sky130_fd_sc_hd__mux2_1
X_16743_ net3181 _14430_ _04612_ VGND VGND VPWR VPWR _04617_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_85_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_3868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_141_3879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19462_ datamem.data_ram\[62\]\[16\] _06719_ _06742_ _06757_ VGND VGND VPWR VPWR
+ _06758_ sky130_fd_sc_hd__o211a_1
X_31740_ net189 _03198_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[9\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16674_ _04580_ VGND VGND VPWR VPWR _01704_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_201_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18413_ _05677_ _05767_ _05774_ _05776_ VGND VGND VPWR VPWR _05777_ sky130_fd_sc_hd__a211o_1
XFILLER_0_115_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15625_ net3976 _13263_ _14114_ VGND VGND VPWR VPWR _14121_ sky130_fd_sc_hd__mux2_1
XFILLER_0_202_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31671_ clknet_leaf_68_clk net1290 VGND VGND VPWR VPWR rvcpu.dp.plmw.ALUResultW\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_19393_ _06608_ VGND VGND VPWR VPWR _06689_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_201_475 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18344_ _05688_ _05663_ VGND VGND VPWR VPWR _05709_ sky130_fd_sc_hd__nand2_2
X_30622_ clknet_leaf_191_clk _02357_ VGND VGND VPWR VPWR datamem.data_ram\[52\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15556_ _13363_ _13575_ _13483_ VGND VGND VPWR VPWR _14080_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_185_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18275_ _05543_ _05549_ _05635_ _05639_ VGND VGND VPWR VPWR _05640_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_72_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30553_ clknet_leaf_180_clk _02288_ VGND VGND VPWR VPWR datamem.data_ram\[55\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_15487_ _13682_ _13399_ _13429_ _14015_ VGND VGND VPWR VPWR _14016_ sky130_fd_sc_hd__a31o_1
XFILLER_0_115_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17226_ _14145_ net4408 _04865_ VGND VGND VPWR VPWR _04873_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_1305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30484_ net162 _02219_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[19\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_249_clk clknet_5_17__leaf_clk VGND VGND VPWR VPWR clknet_leaf_249_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_40_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32223_ clknet_leaf_193_clk _03645_ VGND VGND VPWR VPWR datamem.data_ram\[35\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_17157_ _04836_ VGND VGND VPWR VPWR _01461_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold805 rvcpu.dp.rf.reg_file_arr\[16\]\[12\] VGND VGND VPWR VPWR net1955 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold816 rvcpu.dp.rf.reg_file_arr\[19\]\[2\] VGND VGND VPWR VPWR net1966 sky130_fd_sc_hd__dlygate4sd3_1
Xhold827 rvcpu.dp.rf.reg_file_arr\[3\]\[14\] VGND VGND VPWR VPWR net1977 sky130_fd_sc_hd__dlygate4sd3_1
X_16108_ _14384_ VGND VGND VPWR VPWR _14396_ sky130_fd_sc_hd__buf_4
X_32154_ clknet_leaf_160_clk _03576_ VGND VGND VPWR VPWR datamem.data_ram\[38\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold838 rvcpu.dp.rf.reg_file_arr\[1\]\[0\] VGND VGND VPWR VPWR net1988 sky130_fd_sc_hd__dlygate4sd3_1
X_17088_ _14143_ net2557 _04793_ VGND VGND VPWR VPWR _04800_ sky130_fd_sc_hd__mux2_1
Xhold849 datamem.data_ram\[42\]\[31\] VGND VGND VPWR VPWR net1999 sky130_fd_sc_hd__dlygate4sd3_1
X_31105_ clknet_leaf_108_clk _02840_ VGND VGND VPWR VPWR datamem.data_ram\[19\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16039_ _14359_ VGND VGND VPWR VPWR _02002_ sky130_fd_sc_hd__clkbuf_1
X_32085_ clknet_leaf_64_clk _03507_ VGND VGND VPWR VPWR datamem.data_ram\[47\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2206 rvcpu.dp.rf.reg_file_arr\[16\]\[24\] VGND VGND VPWR VPWR net3356 sky130_fd_sc_hd__dlygate4sd3_1
X_31036_ clknet_leaf_102_clk _02771_ VGND VGND VPWR VPWR datamem.data_ram\[12\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2217 datamem.data_ram\[47\]\[13\] VGND VGND VPWR VPWR net3367 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2228 datamem.data_ram\[17\]\[20\] VGND VGND VPWR VPWR net3378 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_224_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2239 datamem.data_ram\[55\]\[10\] VGND VGND VPWR VPWR net3389 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_200_5301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1505 datamem.data_ram\[12\]\[19\] VGND VGND VPWR VPWR net2655 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1516 datamem.data_ram\[3\]\[23\] VGND VGND VPWR VPWR net2666 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1527 rvcpu.dp.rf.reg_file_arr\[2\]\[5\] VGND VGND VPWR VPWR net2677 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1538 rvcpu.dp.rf.reg_file_arr\[7\]\[28\] VGND VGND VPWR VPWR net2688 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1549 rvcpu.dp.rf.reg_file_arr\[25\]\[0\] VGND VGND VPWR VPWR net2699 sky130_fd_sc_hd__dlygate4sd3_1
X_24159__662 clknet_1_1__leaf__10263_ VGND VGND VPWR VPWR net788 sky130_fd_sc_hd__inv_2
X_23565__188 clknet_1_1__leaf__10175_ VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__inv_2
X_19729_ _06766_ VGND VGND VPWR VPWR _07024_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_0_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32987_ clknet_leaf_199_clk _04409_ VGND VGND VPWR VPWR datamem.data_ram\[62\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_192_5102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_192_5113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22740_ _09875_ _09879_ _09883_ _09491_ VGND VGND VPWR VPWR _01146_ sky130_fd_sc_hd__o31a_1
X_31938_ clknet_leaf_111_clk _03360_ VGND VGND VPWR VPWR datamem.data_ram\[59\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22671_ rvcpu.dp.rf.reg_file_arr\[24\]\[19\] rvcpu.dp.rf.reg_file_arr\[25\]\[19\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[19\] rvcpu.dp.rf.reg_file_arr\[27\]\[19\] _09393_
+ _09465_ VGND VGND VPWR VPWR _09818_ sky130_fd_sc_hd__mux4_1
XFILLER_0_88_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31869_ clknet_leaf_123_clk _03323_ VGND VGND VPWR VPWR datamem.data_ram\[63\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_21622_ _08626_ _08867_ _08869_ _08871_ _08808_ VGND VGND VPWR VPWR _08872_ sky130_fd_sc_hd__a221o_1
XFILLER_0_87_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24410_ _10384_ VGND VGND VPWR VPWR _02315_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25390_ _10946_ _10947_ VGND VGND VPWR VPWR _10948_ sky130_fd_sc_hd__or2_1
XFILLER_0_168_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24051__579 clknet_1_1__leaf__10246_ VGND VGND VPWR VPWR net705 sky130_fd_sc_hd__inv_2
XFILLER_0_192_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_4120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24341_ _10326_ net112 VGND VGND VPWR VPWR _10347_ sky130_fd_sc_hd__nor2_8
XFILLER_0_114_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21553_ rvcpu.dp.plfd.InstrD\[18\] VGND VGND VPWR VPWR _08806_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_151_4131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20504_ datamem.data_ram\[42\]\[21\] _07203_ _07793_ _07794_ VGND VGND VPWR VPWR
+ _07795_ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27060_ _11919_ net4119 _11910_ _11921_ VGND VGND VPWR VPWR _03428_ sky130_fd_sc_hd__a31o_1
X_24272_ _09236_ net4157 _10307_ VGND VGND VPWR VPWR _10309_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21484_ rvcpu.dp.rf.reg_file_arr\[16\]\[6\] rvcpu.dp.rf.reg_file_arr\[17\]\[6\] rvcpu.dp.rf.reg_file_arr\[18\]\[6\]
+ rvcpu.dp.rf.reg_file_arr\[19\]\[6\] _08703_ _08721_ VGND VGND VPWR VPWR _08740_
+ sky130_fd_sc_hd__mux4_1
X_26011_ net19 _11152_ VGND VGND VPWR VPWR _11331_ sky130_fd_sc_hd__or2_1
XFILLER_0_200_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20435_ datamem.data_ram\[19\]\[12\] _06632_ _06780_ datamem.data_ram\[17\]\[12\]
+ _06677_ VGND VGND VPWR VPWR _07727_ sky130_fd_sc_hd__o221a_1
XFILLER_0_99_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_228_5960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload270 clknet_leaf_135_clk VGND VGND VPWR VPWR clkload270/Y sky130_fd_sc_hd__clkinv_4
X_20366_ datamem.data_ram\[38\]\[28\] _06717_ _06685_ datamem.data_ram\[36\]\[28\]
+ VGND VGND VPWR VPWR _07658_ sky130_fd_sc_hd__o22a_1
XFILLER_0_101_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_228_5971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload281 clknet_1_0__leaf__10258_ VGND VGND VPWR VPWR clkload281/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_149_4060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload292 clknet_1_0__leaf__10225_ VGND VGND VPWR VPWR clkload292/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_219_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_4071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22105_ _09315_ VGND VGND VPWR VPWR _01079_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_149_4082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27962_ _09239_ VGND VGND VPWR VPWR _12435_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_101_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20297_ datamem.data_ram\[6\]\[19\] _06764_ _07024_ datamem.data_ram\[4\]\[19\] VGND
+ VGND VPWR VPWR _07590_ sky130_fd_sc_hd__o22a_1
XFILLER_0_105_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_224_5868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29701_ net1047 _01436_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[22\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_224_5879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_181_4850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26913_ _10069_ VGND VGND VPWR VPWR _11833_ sky130_fd_sc_hd__clkbuf_4
X_22036_ rvcpu.dp.plem.WriteDataM\[7\] _09215_ _09219_ _09258_ VGND VGND VPWR VPWR
+ _09259_ sky130_fd_sc_hd__a31o_4
XFILLER_0_228_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27893_ _12391_ net1791 _12393_ _12397_ VGND VGND VPWR VPWR _03785_ sky130_fd_sc_hd__a31o_1
XFILLER_0_41_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29632_ clknet_leaf_148_clk _01367_ VGND VGND VPWR VPWR datamem.data_ram\[5\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2740 datamem.data_ram\[35\]\[27\] VGND VGND VPWR VPWR net3890 sky130_fd_sc_hd__dlygate4sd3_1
X_26844_ _11684_ _11786_ VGND VGND VPWR VPWR _11790_ sky130_fd_sc_hd__and2_1
XFILLER_0_76_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2751 datamem.data_ram\[41\]\[13\] VGND VGND VPWR VPWR net3901 sky130_fd_sc_hd__dlygate4sd3_1
X_24163__5 clknet_1_1__leaf__10264_ VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__inv_2
XFILLER_0_76_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2762 rvcpu.dp.rf.reg_file_arr\[26\]\[16\] VGND VGND VPWR VPWR net3912 sky130_fd_sc_hd__dlygate4sd3_1
X_23051__751 clknet_1_1__leaf__10090_ VGND VGND VPWR VPWR net877 sky130_fd_sc_hd__inv_2
Xhold2773 datamem.data_ram\[43\]\[10\] VGND VGND VPWR VPWR net3923 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2784 datamem.data_ram\[30\]\[29\] VGND VGND VPWR VPWR net3934 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2795 datamem.data_ram\[0\]\[22\] VGND VGND VPWR VPWR net3945 sky130_fd_sc_hd__dlygate4sd3_1
X_29563_ net917 _01298_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[27\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_26775_ _11747_ VGND VGND VPWR VPWR _11748_ sky130_fd_sc_hd__buf_2
XFILLER_0_203_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28514_ _12744_ VGND VGND VPWR VPWR _04059_ sky130_fd_sc_hd__clkbuf_1
X_25726_ _10818_ net3091 _11133_ VGND VGND VPWR VPWR _11137_ sky130_fd_sc_hd__mux2_1
XFILLER_0_225_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22938_ _10067_ _10053_ VGND VGND VPWR VPWR _10068_ sky130_fd_sc_hd__and2_1
X_29494_ net856 _01229_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[28\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_179_4790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28445_ _09350_ _12612_ _12668_ VGND VGND VPWR VPWR _12704_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_80_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25657_ _10783_ _11094_ _11095_ net1322 VGND VGND VPWR VPWR _02851_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_80_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22869_ rvcpu.dp.rf.reg_file_arr\[16\]\[30\] rvcpu.dp.rf.reg_file_arr\[17\]\[30\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[30\] rvcpu.dp.rf.reg_file_arr\[19\]\[30\] _09517_
+ _09513_ VGND VGND VPWR VPWR _10005_ sky130_fd_sc_hd__mux4_1
X_15410_ _13682_ _13378_ _13941_ VGND VGND VPWR VPWR _13942_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_151_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_175_4687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24608_ _10506_ VGND VGND VPWR VPWR _02391_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_175_4698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28376_ _12663_ VGND VGND VPWR VPWR _04002_ sky130_fd_sc_hd__clkbuf_1
X_16390_ _13177_ _14090_ VGND VGND VPWR VPWR _14560_ sky130_fd_sc_hd__nor2_2
X_25588_ _10055_ VGND VGND VPWR VPWR _11057_ sky130_fd_sc_hd__buf_2
XFILLER_0_182_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_3303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_3314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15341_ _13368_ _13646_ _13876_ VGND VGND VPWR VPWR _13877_ sky130_fd_sc_hd__and3_1
X_27327_ _10061_ _12078_ _12079_ net1292 VGND VGND VPWR VPWR _03537_ sky130_fd_sc_hd__o22a_1
XFILLER_0_26_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24539_ _09297_ VGND VGND VPWR VPWR _10465_ sky130_fd_sc_hd__buf_2
XFILLER_0_109_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_227_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18060_ rvcpu.dp.plem.ALUResultM\[9\] _05272_ VGND VGND VPWR VPWR _05428_ sky130_fd_sc_hd__and2_1
X_15272_ _13332_ _13363_ VGND VGND VPWR VPWR _13811_ sky130_fd_sc_hd__nand2_1
X_27258_ _10061_ net52 _12042_ net1360 VGND VGND VPWR VPWR _03505_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17011_ _04759_ VGND VGND VPWR VPWR _01530_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_78_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26209_ net1652 _11442_ _03038_ _11443_ VGND VGND VPWR VPWR _03055_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27189_ _11991_ net1410 _11995_ _12002_ VGND VGND VPWR VPWR _03476_ sky130_fd_sc_hd__a31o_1
XFILLER_0_123_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24028__559 clknet_1_0__leaf__10243_ VGND VGND VPWR VPWR net685 sky130_fd_sc_hd__inv_2
XFILLER_0_225_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18962_ _05694_ _06297_ _06298_ _05703_ VGND VGND VPWR VPWR _06299_ sky130_fd_sc_hd__o211a_1
XFILLER_0_192_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17913_ rvcpu.dp.plde.RD1E\[30\] _05265_ _05269_ _13183_ _05285_ VGND VGND VPWR VPWR
+ _05286_ sky130_fd_sc_hd__a221o_2
XFILLER_0_28_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18893_ _05465_ _05785_ _06108_ _05466_ VGND VGND VPWR VPWR _06235_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_28_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17844_ rvcpu.dp.plem.ALUResultM\[15\] _05223_ _05175_ VGND VGND VPWR VPWR _05224_
+ sky130_fd_sc_hd__mux2_1
X_23484__131 clknet_1_1__leaf__10159_ VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__inv_2
X_32910_ clknet_leaf_174_clk _04332_ VGND VGND VPWR VPWR datamem.data_ram\[7\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_32841_ clknet_leaf_96_clk _04263_ VGND VGND VPWR VPWR datamem.data_ram\[7\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_17775_ _05154_ _05161_ rvcpu.dp.plde.RD2E\[0\] VGND VGND VPWR VPWR _05173_ sky130_fd_sc_hd__a21bo_1
X_14987_ _13479_ _13530_ _13534_ _13439_ VGND VGND VPWR VPWR _13535_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_178_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19514_ _06741_ VGND VGND VPWR VPWR _06810_ sky130_fd_sc_hd__buf_8
X_16726_ _04607_ VGND VGND VPWR VPWR _01679_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32772_ clknet_leaf_233_clk _04194_ VGND VGND VPWR VPWR datamem.data_ram\[14\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_18_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19445_ _06599_ VGND VGND VPWR VPWR _06741_ sky130_fd_sc_hd__buf_8
X_31723_ net172 _03181_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[9\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_187_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16657_ _14189_ net2979 _04562_ VGND VGND VPWR VPWR _04571_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_102_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15608_ net1901 _13238_ _14103_ VGND VGND VPWR VPWR _14112_ sky130_fd_sc_hd__mux2_1
X_31654_ clknet_leaf_66_clk net1742 VGND VGND VPWR VPWR rvcpu.dp.plmw.ALUResultW\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19376_ _06671_ VGND VGND VPWR VPWR _06672_ sky130_fd_sc_hd__clkbuf_8
X_16588_ _14189_ net2863 _04525_ VGND VGND VPWR VPWR _04534_ sky130_fd_sc_hd__mux2_1
XFILLER_0_173_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18327_ _05370_ VGND VGND VPWR VPWR _05692_ sky130_fd_sc_hd__buf_2
X_30605_ clknet_leaf_207_clk _02340_ VGND VGND VPWR VPWR datamem.data_ram\[52\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_15539_ _13665_ _13294_ _13559_ _13689_ _13483_ VGND VGND VPWR VPWR _14065_ sky130_fd_sc_hd__a221o_1
X_31585_ clknet_leaf_52_clk net1241 VGND VGND VPWR VPWR rvcpu.dp.plmw.PCPlus4W\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18258_ _05473_ _05622_ _05478_ VGND VGND VPWR VPWR _05623_ sky130_fd_sc_hd__or3_1
XFILLER_0_155_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30536_ clknet_leaf_218_clk _02271_ VGND VGND VPWR VPWR datamem.data_ram\[55\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17209_ _04863_ VGND VGND VPWR VPWR _01436_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_555 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18189_ _05539_ _05540_ VGND VGND VPWR VPWR _05554_ sky130_fd_sc_hd__or2_1
X_30467_ net145 _02202_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[19\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold602 datamem.data_ram\[61\]\[3\] VGND VGND VPWR VPWR net1752 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold613 datamem.data_ram\[8\]\[3\] VGND VGND VPWR VPWR net1763 sky130_fd_sc_hd__dlygate4sd3_1
X_20220_ datamem.data_ram\[22\]\[3\] _07127_ _06976_ datamem.data_ram\[20\]\[3\] VGND
+ VGND VPWR VPWR _07513_ sky130_fd_sc_hd__a22o_1
X_32206_ clknet_leaf_88_clk _03628_ VGND VGND VPWR VPWR datamem.data_ram\[36\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold624 datamem.data_ram\[51\]\[7\] VGND VGND VPWR VPWR net1774 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_1110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold635 rvcpu.dp.plfd.InstrD\[9\] VGND VGND VPWR VPWR net1785 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30398_ net736 _02133_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[31\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold646 datamem.data_ram\[26\]\[7\] VGND VGND VPWR VPWR net1796 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold657 rvcpu.dp.plfd.PCD\[7\] VGND VGND VPWR VPWR net1807 sky130_fd_sc_hd__dlygate4sd3_1
Xhold668 datamem.data_ram\[61\]\[6\] VGND VGND VPWR VPWR net1818 sky130_fd_sc_hd__dlygate4sd3_1
X_32137_ clknet_leaf_242_clk _03559_ VGND VGND VPWR VPWR datamem.data_ram\[39\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_20151_ datamem.data_ram\[54\]\[27\] _06626_ _06811_ datamem.data_ram\[48\]\[27\]
+ VGND VGND VPWR VPWR _07444_ sky130_fd_sc_hd__o22a_1
Xhold679 datamem.data_ram\[53\]\[1\] VGND VGND VPWR VPWR net1829 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2003 rvcpu.dp.rf.reg_file_arr\[30\]\[27\] VGND VGND VPWR VPWR net3153 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32068_ clknet_leaf_126_clk _03490_ VGND VGND VPWR VPWR datamem.data_ram\[29\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_20082_ datamem.data_ram\[32\]\[10\] _06821_ _06789_ datamem.data_ram\[33\]\[10\]
+ _07375_ VGND VGND VPWR VPWR _07376_ sky130_fd_sc_hd__o221a_1
XFILLER_0_176_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2014 rvcpu.dp.rf.reg_file_arr\[29\]\[10\] VGND VGND VPWR VPWR net3164 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2025 rvcpu.dp.rf.reg_file_arr\[4\]\[2\] VGND VGND VPWR VPWR net3175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2036 datamem.data_ram\[63\]\[22\] VGND VGND VPWR VPWR net3186 sky130_fd_sc_hd__dlygate4sd3_1
X_31019_ clknet_leaf_156_clk _02754_ VGND VGND VPWR VPWR datamem.data_ram\[42\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1302 rvcpu.dp.rf.reg_file_arr\[17\]\[12\] VGND VGND VPWR VPWR net2452 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2047 datamem.data_ram\[49\]\[29\] VGND VGND VPWR VPWR net3197 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1313 datamem.data_ram\[6\]\[13\] VGND VGND VPWR VPWR net2463 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_176_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24890_ _10444_ net3930 _10659_ VGND VGND VPWR VPWR _10662_ sky130_fd_sc_hd__mux2_1
Xhold2058 datamem.data_ram\[54\]\[31\] VGND VGND VPWR VPWR net3208 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2069 rvcpu.dp.rf.reg_file_arr\[15\]\[9\] VGND VGND VPWR VPWR net3219 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1324 datamem.data_ram\[15\]\[27\] VGND VGND VPWR VPWR net2474 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1335 rvcpu.dp.rf.reg_file_arr\[11\]\[4\] VGND VGND VPWR VPWR net2485 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1346 datamem.data_ram\[13\]\[8\] VGND VGND VPWR VPWR net2496 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1357 datamem.data_ram\[34\]\[16\] VGND VGND VPWR VPWR net2507 sky130_fd_sc_hd__dlygate4sd3_1
X_23841_ _09326_ net2442 _10210_ VGND VGND VPWR VPWR _10217_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1368 rvcpu.dp.rf.reg_file_arr\[10\]\[15\] VGND VGND VPWR VPWR net2518 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_1264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1379 datamem.data_ram\[7\]\[10\] VGND VGND VPWR VPWR net2529 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_508 _13212_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26560_ _10820_ net2826 _11620_ VGND VGND VPWR VPWR _11625_ sky130_fd_sc_hd__mux2_1
X_20984_ datamem.data_ram\[10\]\[15\] datamem.data_ram\[11\]\[15\] _06651_ VGND VGND
+ VPWR VPWR _08273_ sky130_fd_sc_hd__mux2_1
XANTENNA_519 _13251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25511_ _10408_ _11010_ VGND VGND VPWR VPWR _11012_ sky130_fd_sc_hd__and2_1
Xclkbuf_0__10160_ _10160_ VGND VGND VPWR VPWR clknet_0__10160_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_67_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22723_ rvcpu.dp.rf.reg_file_arr\[16\]\[22\] rvcpu.dp.rf.reg_file_arr\[17\]\[22\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[22\] rvcpu.dp.rf.reg_file_arr\[19\]\[22\] _09385_
+ _09637_ VGND VGND VPWR VPWR _09867_ sky130_fd_sc_hd__mux4_1
X_26491_ clknet_1_1__leaf__10079_ VGND VGND VPWR VPWR _11601_ sky130_fd_sc_hd__buf_1
XFILLER_0_220_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28230_ _12584_ VGND VGND VPWR VPWR _03935_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25442_ _10977_ VGND VGND VPWR VPWR _02754_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__10091_ _10091_ VGND VGND VPWR VPWR clknet_0__10091_ sky130_fd_sc_hd__clkbuf_16
X_22654_ _09391_ _09801_ VGND VGND VPWR VPWR _09802_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_217_5694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28161_ _12547_ VGND VGND VPWR VPWR _03903_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21605_ _08533_ VGND VGND VPWR VPWR _08856_ sky130_fd_sc_hd__buf_4
X_25373_ _10055_ VGND VGND VPWR VPWR _10938_ sky130_fd_sc_hd__buf_2
X_22585_ _09636_ _09736_ VGND VGND VPWR VPWR _09737_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_211_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27112_ _11938_ net1778 _11952_ _11954_ VGND VGND VPWR VPWR _03447_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_4573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24324_ _10325_ _10337_ _10269_ VGND VGND VPWR VPWR _10338_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_63_656 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_170_4584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28092_ _12447_ net3826 net75 VGND VGND VPWR VPWR _12511_ sky130_fd_sc_hd__mux2_1
X_21536_ _08663_ _08787_ _08789_ _08575_ VGND VGND VPWR VPWR _08790_ sky130_fd_sc_hd__o211a_1
XFILLER_0_145_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27043_ _11822_ _11911_ VGND VGND VPWR VPWR _11912_ sky130_fd_sc_hd__and2_1
X_21467_ _08722_ _08723_ _08541_ VGND VGND VPWR VPWR _08724_ sky130_fd_sc_hd__mux2_1
X_24255_ _09306_ net2285 _10298_ VGND VGND VPWR VPWR _10300_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_177_Right_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_226_5908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_226_5919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_189_Left_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20418_ datamem.data_ram\[54\]\[12\] _06743_ _06645_ datamem.data_ram\[48\]\[12\]
+ _07709_ VGND VGND VPWR VPWR _07710_ sky130_fd_sc_hd__o221a_1
XFILLER_0_160_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_147_4019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21398_ _08532_ _08657_ VGND VGND VPWR VPWR _08658_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_73_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20349_ datamem.data_ram\[54\]\[4\] _06951_ _06931_ datamem.data_ram\[50\]\[4\] _06601_
+ VGND VGND VPWR VPWR _07641_ sky130_fd_sc_hd__a221o_1
X_23435__86 clknet_1_1__leaf__10155_ VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__inv_2
XFILLER_0_219_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28994_ _13006_ VGND VGND VPWR VPWR _04277_ sky130_fd_sc_hd__clkbuf_1
X_27945_ _12363_ net3968 _12421_ VGND VGND VPWR VPWR _12425_ sky130_fd_sc_hd__mux2_1
X_23068_ _09276_ net4398 _10093_ VGND VGND VPWR VPWR _10096_ sky130_fd_sc_hd__mux2_1
X_24101__609 clknet_1_1__leaf__10258_ VGND VGND VPWR VPWR net735 sky130_fd_sc_hd__inv_2
XFILLER_0_179_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3260 rvcpu.dp.rf.reg_file_arr\[22\]\[27\] VGND VGND VPWR VPWR net4410 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14910_ _13321_ _13459_ _13337_ VGND VGND VPWR VPWR _13460_ sky130_fd_sc_hd__a21o_1
Xhold3271 datamem.data_ram\[58\]\[16\] VGND VGND VPWR VPWR net4421 sky130_fd_sc_hd__dlygate4sd3_1
X_22019_ _09245_ VGND VGND VPWR VPWR _01063_ sky130_fd_sc_hd__clkbuf_1
Xhold3282 rvcpu.dp.rf.reg_file_arr\[15\]\[11\] VGND VGND VPWR VPWR net4432 sky130_fd_sc_hd__dlygate4sd3_1
X_27876_ _12151_ net3352 net77 VGND VGND VPWR VPWR _12387_ sky130_fd_sc_hd__mux2_1
X_15890_ net2894 _13195_ _14275_ VGND VGND VPWR VPWR _14280_ sky130_fd_sc_hd__mux2_1
XFILLER_0_216_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold3293 rvcpu.dp.rf.reg_file_arr\[24\]\[2\] VGND VGND VPWR VPWR net4443 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_175_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2570 datamem.data_ram\[11\]\[25\] VGND VGND VPWR VPWR net3720 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26827_ _11767_ net1467 _11773_ _11779_ VGND VGND VPWR VPWR _03337_ sky130_fd_sc_hd__a31o_1
X_14841_ _13291_ _13346_ _13393_ VGND VGND VPWR VPWR _13394_ sky130_fd_sc_hd__and3_1
Xhold2581 rvcpu.dp.rf.reg_file_arr\[29\]\[14\] VGND VGND VPWR VPWR net3731 sky130_fd_sc_hd__dlygate4sd3_1
X_29615_ net969 _01350_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[25\]\[18\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_106_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2592 datamem.data_ram\[22\]\[11\] VGND VGND VPWR VPWR net3742 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_198_Left_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1880 rvcpu.dp.rf.reg_file_arr\[14\]\[21\] VGND VGND VPWR VPWR net3030 sky130_fd_sc_hd__dlygate4sd3_1
X_29546_ net900 _01281_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[27\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_17560_ _05050_ VGND VGND VPWR VPWR _01256_ sky130_fd_sc_hd__clkbuf_1
X_26758_ _11676_ _11738_ VGND VGND VPWR VPWR _11739_ sky130_fd_sc_hd__and2_1
X_14772_ _13317_ _13319_ _13324_ rvcpu.dp.pcreg.q\[9\] VGND VGND VPWR VPWR _13325_
+ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_177_4738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1891 datamem.data_ram\[7\]\[19\] VGND VGND VPWR VPWR net3041 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_177_4749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16511_ _04493_ VGND VGND VPWR VPWR _01788_ sky130_fd_sc_hd__clkbuf_1
X_25709_ _10818_ net3730 _11124_ VGND VGND VPWR VPWR _11128_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29477_ net839 _01212_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[2\]\[16\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__10258_ clknet_0__10258_ VGND VGND VPWR VPWR clknet_1_1__leaf__10258_
+ sky130_fd_sc_hd__clkbuf_16
X_17491_ _13190_ net3118 _05010_ VGND VGND VPWR VPWR _05014_ sky130_fd_sc_hd__mux2_1
X_26689_ _11683_ net1714 _11693_ _11698_ VGND VGND VPWR VPWR _03280_ sky130_fd_sc_hd__a31o_1
XFILLER_0_196_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19230_ rvcpu.dp.plde.ImmExtE\[27\] rvcpu.dp.plde.PCE\[27\] VGND VGND VPWR VPWR _06536_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16442_ net2371 _14472_ _04451_ VGND VGND VPWR VPWR _04456_ sky130_fd_sc_hd__mux2_1
X_28428_ _12692_ net2852 _12688_ VGND VGND VPWR VPWR _12693_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19161_ _06471_ net38 _06475_ VGND VGND VPWR VPWR _06476_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_144_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28359_ _12654_ VGND VGND VPWR VPWR _03994_ sky130_fd_sc_hd__clkbuf_1
X_16373_ _14551_ VGND VGND VPWR VPWR _01852_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_136_3756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18112_ _05475_ _05478_ VGND VGND VPWR VPWR _05479_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15324_ _13442_ _13852_ _13854_ _13856_ _13860_ VGND VGND VPWR VPWR _13861_ sky130_fd_sc_hd__o311a_1
XFILLER_0_186_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_3767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19092_ _06413_ _06414_ VGND VGND VPWR VPWR _06415_ sky130_fd_sc_hd__and2b_1
X_31370_ clknet_leaf_17_clk _03073_ VGND VGND VPWR VPWR rvcpu.dp.plde.ImmExtE\[19\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_26_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22962__671 clknet_1_0__leaf__10081_ VGND VGND VPWR VPWR net797 sky130_fd_sc_hd__inv_2
XFILLER_0_48_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_227_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18043_ _13247_ rvcpu.dp.plde.RD2E\[10\] _05195_ VGND VGND VPWR VPWR _05413_ sky130_fd_sc_hd__mux2_1
X_30321_ net667 _02056_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[4\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15255_ _13438_ _13794_ VGND VGND VPWR VPWR _13795_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_1154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_144_Right_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30252_ net606 _01987_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[6\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_15186_ _13451_ _13728_ VGND VGND VPWR VPWR _13729_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_39_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__10080_ clknet_0__10080_ VGND VGND VPWR VPWR clknet_1_0__leaf__10080_
+ sky130_fd_sc_hd__clkbuf_16
X_23058__757 clknet_1_0__leaf__10091_ VGND VGND VPWR VPWR net883 sky130_fd_sc_hd__inv_2
XFILLER_0_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30183_ net537 _01918_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[8\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_19994_ datamem.data_ram\[22\]\[2\] _06951_ _06936_ datamem.data_ram\[16\]\[2\] VGND
+ VGND VPWR VPWR _07288_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18945_ _06230_ _06282_ _05707_ VGND VGND VPWR VPWR _06283_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18876_ _05658_ _06216_ _06218_ _06109_ _06004_ VGND VGND VPWR VPWR _06219_ sky130_fd_sc_hd__o221a_1
XFILLER_0_222_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17827_ _05212_ VGND VGND VPWR VPWR rvcpu.dp.SrcBFW_Mux.y\[24\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_55_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23720__313 clknet_1_1__leaf__10197_ VGND VGND VPWR VPWR net439 sky130_fd_sc_hd__inv_2
X_32824_ clknet_leaf_186_clk _04246_ VGND VGND VPWR VPWR datamem.data_ram\[12\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_17758_ _14346_ rvcpu.dp.plde.Rs2E\[0\] rvcpu.dp.plde.Rs2E\[3\] _13175_ _05155_ VGND
+ VGND VPWR VPWR _05156_ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16709_ _14172_ net4432 _04598_ VGND VGND VPWR VPWR _04599_ sky130_fd_sc_hd__mux2_1
X_32755_ clknet_leaf_166_clk _04177_ VGND VGND VPWR VPWR datamem.data_ram\[15\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_17689_ _13173_ net3938 _05118_ VGND VGND VPWR VPWR _05119_ sky130_fd_sc_hd__mux2_1
Xclkbuf_5_1__f_clk clknet_2_0_0_clk VGND VGND VPWR VPWR clknet_5_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_9_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31706_ clknet_leaf_31_clk _03164_ VGND VGND VPWR VPWR rvcpu.dp.pcreg.q\[24\] sky130_fd_sc_hd__dfxtp_1
X_19428_ _06723_ VGND VGND VPWR VPWR _06724_ sky130_fd_sc_hd__clkbuf_8
X_32686_ clknet_leaf_84_clk _04108_ VGND VGND VPWR VPWR datamem.data_ram\[18\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31637_ clknet_leaf_47_clk net1181 VGND VGND VPWR VPWR rvcpu.dp.plmw.lAuiPCW\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19359_ _06654_ VGND VGND VPWR VPWR _06655_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_174_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22370_ rvcpu.dp.rf.reg_file_arr\[8\]\[3\] rvcpu.dp.rf.reg_file_arr\[10\]\[3\] rvcpu.dp.rf.reg_file_arr\[9\]\[3\]
+ rvcpu.dp.rf.reg_file_arr\[11\]\[3\] _09431_ _09532_ VGND VGND VPWR VPWR _09533_
+ sky130_fd_sc_hd__mux4_1
X_31568_ clknet_leaf_62_clk datamem.rd_data_mem\[18\] VGND VGND VPWR VPWR rvcpu.dp.plmw.ReadDataW\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_212_5580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_212_5591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21321_ rvcpu.dp.plfd.InstrD\[18\] _08582_ rvcpu.dp.plde.RdE\[4\] _08509_ VGND VGND
+ VPWR VPWR _08583_ sky130_fd_sc_hd__a22o_1
XFILLER_0_142_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30519_ clknet_leaf_144_clk _02254_ VGND VGND VPWR VPWR datamem.data_ram\[56\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31499_ clknet_leaf_26_clk rvcpu.dp.lAuiPCE\[25\] VGND VGND VPWR VPWR rvcpu.dp.plem.lAuiPCM\[25\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold410 datamem.data_ram\[22\]\[7\] VGND VGND VPWR VPWR net1560 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_111_Right_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21252_ rvcpu.dp.plfd.InstrD\[17\] VGND VGND VPWR VPWR _08514_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_29_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold421 rvcpu.dp.plfd.PCPlus4D\[7\] VGND VGND VPWR VPWR net1571 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold432 datamem.data_ram\[38\]\[7\] VGND VGND VPWR VPWR net1582 sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 rvcpu.dp.plfd.PCD\[8\] VGND VGND VPWR VPWR net1593 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20203_ datamem.data_ram\[56\]\[11\] _06778_ _07494_ _07495_ VGND VGND VPWR VPWR
+ _07496_ sky130_fd_sc_hd__o211a_1
Xhold454 datamem.data_ram\[37\]\[3\] VGND VGND VPWR VPWR net1604 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21183_ rvcpu.dp.plem.funct3M\[0\] rvcpu.dp.plem.funct3M\[1\] rvcpu.dp.plem.funct3M\[2\]
+ VGND VGND VPWR VPWR _08470_ sky130_fd_sc_hd__nor3_1
XFILLER_0_111_750 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold465 datamem.data_ram\[10\]\[0\] VGND VGND VPWR VPWR net1615 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold476 rvcpu.dp.plem.ALUResultM\[5\] VGND VGND VPWR VPWR net1626 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold487 datamem.data_ram\[36\]\[2\] VGND VGND VPWR VPWR net1637 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_221_5805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold498 datamem.data_ram\[33\]\[3\] VGND VGND VPWR VPWR net1648 sky130_fd_sc_hd__dlygate4sd3_1
X_20134_ datamem.data_ram\[34\]\[27\] _06610_ _06805_ datamem.data_ram\[36\]\[27\]
+ VGND VGND VPWR VPWR _07427_ sky130_fd_sc_hd__o22a_1
X_23881__442 clknet_1_1__leaf__10221_ VGND VGND VPWR VPWR net568 sky130_fd_sc_hd__inv_2
XFILLER_0_217_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25991_ net9 _11317_ VGND VGND VPWR VPWR _11320_ sky130_fd_sc_hd__or2_1
XFILLER_0_229_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27730_ _12091_ net3065 net49 VGND VGND VPWR VPWR _12304_ sky130_fd_sc_hd__mux2_1
XFILLER_0_216_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24942_ _10444_ net3136 _10687_ VGND VGND VPWR VPWR _10690_ sky130_fd_sc_hd__mux2_1
X_20065_ _07354_ _07356_ _07358_ VGND VGND VPWR VPWR _07359_ sky130_fd_sc_hd__and3_1
Xhold1110 rvcpu.dp.rf.reg_file_arr\[23\]\[29\] VGND VGND VPWR VPWR net2260 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1121 datamem.data_ram\[39\]\[30\] VGND VGND VPWR VPWR net2271 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_176_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1132 datamem.data_ram\[14\]\[20\] VGND VGND VPWR VPWR net2282 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27661_ _12153_ net3345 net79 VGND VGND VPWR VPWR _12267_ sky130_fd_sc_hd__mux2_1
XFILLER_0_225_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24873_ _10470_ net3844 net92 VGND VGND VPWR VPWR _10653_ sky130_fd_sc_hd__mux2_1
Xhold1143 rvcpu.dp.rf.reg_file_arr\[1\]\[2\] VGND VGND VPWR VPWR net2293 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1154 rvcpu.dp.rf.reg_file_arr\[16\]\[8\] VGND VGND VPWR VPWR net2304 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1165 datamem.data_ram\[9\]\[16\] VGND VGND VPWR VPWR net2315 sky130_fd_sc_hd__dlygate4sd3_1
X_29400_ clknet_leaf_0_clk _01135_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD2E\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_213_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26612_ _10818_ net3277 _11650_ VGND VGND VPWR VPWR _11654_ sky130_fd_sc_hd__mux2_1
Xhold1176 rvcpu.dp.rf.reg_file_arr\[4\]\[8\] VGND VGND VPWR VPWR net2326 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1187 datamem.data_ram\[29\]\[22\] VGND VGND VPWR VPWR net2337 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27592_ _12136_ net2859 _12224_ VGND VGND VPWR VPWR _12230_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_219_5745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_305 _14151_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1198 rvcpu.dp.rf.reg_file_arr\[25\]\[15\] VGND VGND VPWR VPWR net2348 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_316 _14177_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_219_5756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29331_ clknet_leaf_140_clk _01066_ VGND VGND VPWR VPWR datamem.data_ram\[62\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__10112_ clknet_0__10112_ VGND VGND VPWR VPWR clknet_1_1__leaf__10112_
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_327 _14455_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26543_ _11517_ net1548 _11608_ _11615_ VGND VGND VPWR VPWR _03217_ sky130_fd_sc_hd__a31o_1
XANTENNA_338 _14463_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_212_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23755_ clknet_1_1__leaf__10192_ VGND VGND VPWR VPWR _10201_ sky130_fd_sc_hd__buf_1
XFILLER_0_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20967_ datamem.data_ram\[36\]\[15\] datamem.data_ram\[37\]\[15\] _06651_ VGND VGND
+ VPWR VPWR _08256_ sky130_fd_sc_hd__mux2_1
XANTENNA_349 datamem.data_ram\[53\]\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_172_4613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29262_ _09272_ net3480 _13150_ VGND VGND VPWR VPWR _13152_ sky130_fd_sc_hd__mux2_1
X_22706_ rvcpu.dp.rf.reg_file_arr\[20\]\[21\] rvcpu.dp.rf.reg_file_arr\[21\]\[21\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[21\] rvcpu.dp.rf.reg_file_arr\[23\]\[21\] _09434_
+ _09558_ VGND VGND VPWR VPWR _09851_ sky130_fd_sc_hd__mux4_1
X_26474_ net4452 _11573_ _11594_ _10041_ VGND VGND VPWR VPWR _03169_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_172_4624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_4635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20898_ _08186_ _08187_ _07822_ VGND VGND VPWR VPWR _08188_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28213_ _12575_ VGND VGND VPWR VPWR _03927_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25425_ _10968_ VGND VGND VPWR VPWR _02746_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22637_ _09510_ _09779_ _09781_ _09785_ _09525_ VGND VGND VPWR VPWR _09786_ sky130_fd_sc_hd__a311o_1
X_29193_ _13114_ VGND VGND VPWR VPWR _04368_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28144_ _12538_ VGND VGND VPWR VPWR _03895_ sky130_fd_sc_hd__clkbuf_1
X_25356_ _10413_ _10923_ VGND VGND VPWR VPWR _10927_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22568_ _09381_ VGND VGND VPWR VPWR _09721_ sky130_fd_sc_hd__buf_4
XFILLER_0_134_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24307_ _09298_ net3096 _10328_ VGND VGND VPWR VPWR _10329_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28075_ _12430_ net4207 _12501_ VGND VGND VPWR VPWR _12502_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21519_ rvcpu.dp.rf.reg_file_arr\[8\]\[7\] rvcpu.dp.rf.reg_file_arr\[10\]\[7\] rvcpu.dp.rf.reg_file_arr\[9\]\[7\]
+ rvcpu.dp.rf.reg_file_arr\[11\]\[7\] _08649_ _08537_ VGND VGND VPWR VPWR _08774_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_131_3631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25287_ _10739_ net2307 _10878_ VGND VGND VPWR VPWR _10886_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_131_3642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22499_ _09495_ _09654_ VGND VGND VPWR VPWR _09655_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_20_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27026_ _11889_ net1629 _11897_ _11901_ VGND VGND VPWR VPWR _03414_ sky130_fd_sc_hd__a31o_1
X_15040_ _13398_ _13322_ _13586_ VGND VGND VPWR VPWR _13587_ sky130_fd_sc_hd__or3_1
X_24238_ _10290_ VGND VGND VPWR VPWR _02237_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16991_ net1879 _14474_ _04742_ VGND VGND VPWR VPWR _04748_ sky130_fd_sc_hd__mux2_1
X_28977_ _12995_ net1368 _12988_ _12997_ VGND VGND VPWR VPWR _04269_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_34_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23131__807 clknet_1_0__leaf__10106_ VGND VGND VPWR VPWR net933 sky130_fd_sc_hd__inv_2
XFILLER_0_78_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_990 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18730_ _05406_ _05433_ _05451_ VGND VGND VPWR VPWR _06082_ sky130_fd_sc_hd__a21o_1
XFILLER_0_120_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15942_ net3175 _13272_ _14297_ VGND VGND VPWR VPWR _14307_ sky130_fd_sc_hd__mux2_1
X_27928_ _12132_ net4332 _12412_ VGND VGND VPWR VPWR _12416_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_129_3582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_3593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3090 datamem.data_ram\[11\]\[13\] VGND VGND VPWR VPWR net4240 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_30_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18661_ _06015_ _05431_ VGND VGND VPWR VPWR _06016_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_204_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27859_ _12134_ net2233 _12373_ VGND VGND VPWR VPWR _12378_ sky130_fd_sc_hd__mux2_1
X_15873_ net2883 _13275_ _14235_ VGND VGND VPWR VPWR _14269_ sky130_fd_sc_hd__mux2_1
XFILLER_0_215_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_203_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14824_ _13288_ _13306_ VGND VGND VPWR VPWR _13377_ sky130_fd_sc_hd__or2_1
XFILLER_0_215_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17612_ _05077_ VGND VGND VPWR VPWR _01231_ sky130_fd_sc_hd__clkbuf_1
X_30870_ clknet_leaf_62_clk _02605_ VGND VGND VPWR VPWR datamem.data_ram\[42\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_18592_ _05776_ _05947_ _05948_ _05782_ _05950_ VGND VGND VPWR VPWR _05951_ sky130_fd_sc_hd__o32a_1
XFILLER_0_192_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17543_ _13269_ net2431 _05032_ VGND VGND VPWR VPWR _05041_ sky130_fd_sc_hd__mux2_1
X_14755_ _13305_ _13307_ VGND VGND VPWR VPWR _13308_ sky130_fd_sc_hd__nor2_4
X_29529_ clknet_leaf_264_clk _01264_ VGND VGND VPWR VPWR datamem.data_ram\[5\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32540_ clknet_leaf_80_clk _03962_ VGND VGND VPWR VPWR datamem.data_ram\[23\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_138_3818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17474_ _05004_ VGND VGND VPWR VPWR _01304_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_213_Right_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14686_ _13249_ VGND VGND VPWR VPWR _03182_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_28_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19213_ _06520_ _06517_ _06514_ VGND VGND VPWR VPWR _06521_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_28_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16425_ net3051 _14455_ _14572_ VGND VGND VPWR VPWR _14579_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32471_ clknet_leaf_79_clk _03893_ VGND VGND VPWR VPWR datamem.data_ram\[26\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31422_ clknet_leaf_103_clk _03125_ VGND VGND VPWR VPWR datamem.data_ram\[15\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_19144_ _06457_ _06460_ VGND VGND VPWR VPWR _06461_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_172_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16356_ _14542_ VGND VGND VPWR VPWR _01860_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_99_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15307_ _13466_ _13840_ _13844_ VGND VGND VPWR VPWR _13845_ sky130_fd_sc_hd__a21oi_1
X_19075_ rvcpu.dp.plde.ImmExtE\[8\] rvcpu.dp.plde.PCE\[8\] VGND VGND VPWR VPWR _06400_
+ sky130_fd_sc_hd__or2_1
X_31353_ clknet_leaf_17_clk _03056_ VGND VGND VPWR VPWR rvcpu.dp.plde.ImmExtE\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_26_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__10201_ clknet_0__10201_ VGND VGND VPWR VPWR clknet_1_0__leaf__10201_
+ sky130_fd_sc_hd__clkbuf_16
X_16287_ net4281 _14453_ _14500_ VGND VGND VPWR VPWR _14506_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18026_ _05384_ _05385_ _05388_ VGND VGND VPWR VPWR _05396_ sky130_fd_sc_hd__a21oi_1
X_30304_ net650 _02039_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[5\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_15238_ _13542_ _13525_ _13717_ _13317_ _13438_ VGND VGND VPWR VPWR _13778_ sky130_fd_sc_hd__a221o_1
X_31284_ clknet_leaf_112_clk _02987_ VGND VGND VPWR VPWR datamem.data_ram\[34\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__10132_ clknet_0__10132_ VGND VGND VPWR VPWR clknet_1_0__leaf__10132_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_160_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30235_ net589 _01970_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[7\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_15169_ _13705_ _13712_ _13572_ VGND VGND VPWR VPWR _13713_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_58_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_205_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30166_ net528 _01901_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[0\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_23414__67 clknet_1_1__leaf__10153_ VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__inv_2
X_19977_ datamem.data_ram\[22\]\[18\] _06744_ _06646_ datamem.data_ram\[16\]\[18\]
+ _07270_ VGND VGND VPWR VPWR _07271_ sky130_fd_sc_hd__o221a_1
XFILLER_0_157_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18928_ _06252_ _05630_ _06266_ VGND VGND VPWR VPWR _06267_ sky130_fd_sc_hd__a21o_1
XFILLER_0_66_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30097_ net459 _01832_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[11\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18859_ _06109_ _06202_ VGND VGND VPWR VPWR _06203_ sky130_fd_sc_hd__nor2_1
XFILLER_0_206_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_207_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_206_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21870_ _08842_ _09106_ VGND VGND VPWR VPWR _09107_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32807_ clknet_leaf_156_clk _04229_ VGND VGND VPWR VPWR datamem.data_ram\[13\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_20821_ _08109_ _08110_ _07833_ VGND VGND VPWR VPWR _08111_ sky130_fd_sc_hd__a21o_1
XFILLER_0_221_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30999_ clknet_leaf_102_clk _02734_ VGND VGND VPWR VPWR datamem.data_ram\[22\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_212_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_203_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22969__677 clknet_1_1__leaf__10082_ VGND VGND VPWR VPWR net803 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_214_5620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20752_ datamem.data_ram\[14\]\[6\] _07829_ VGND VGND VPWR VPWR _08042_ sky130_fd_sc_hd__or2_1
XFILLER_0_147_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32738_ clknet_leaf_285_clk _04160_ VGND VGND VPWR VPWR datamem.data_ram\[16\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_212_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_214_5631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_214_5642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24130__635 clknet_1_1__leaf__10261_ VGND VGND VPWR VPWR net761 sky130_fd_sc_hd__inv_2
X_20683_ datamem.data_ram\[32\]\[5\] _07122_ _07972_ _07973_ VGND VGND VPWR VPWR _07974_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_148_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_623 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32669_ clknet_leaf_287_clk _04091_ VGND VGND VPWR VPWR datamem.data_ram\[19\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25210_ _10820_ net3596 net56 VGND VGND VPWR VPWR _10844_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_210_5528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22422_ _09390_ _09581_ VGND VGND VPWR VPWR _09582_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_210_5539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26190_ _11413_ VGND VGND VPWR VPWR _11432_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25141_ _10751_ net3908 _10802_ VGND VGND VPWR VPWR _10803_ sky130_fd_sc_hd__mux2_1
X_22353_ _09398_ VGND VGND VPWR VPWR _09516_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_182_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21304_ _08549_ VGND VGND VPWR VPWR _08566_ sky130_fd_sc_hd__clkbuf_8
X_25072_ _10766_ net3410 _10752_ VGND VGND VPWR VPWR _10767_ sky130_fd_sc_hd__mux2_1
X_22284_ _09421_ VGND VGND VPWR VPWR _09449_ sky130_fd_sc_hd__buf_4
XFILLER_0_206_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28900_ _12743_ net4286 net68 VGND VGND VPWR VPWR _12955_ sky130_fd_sc_hd__mux2_1
X_24023_ clknet_1_0__leaf__10224_ VGND VGND VPWR VPWR _10243_ sky130_fd_sc_hd__buf_1
X_21235_ datamem.data_ram\[53\]\[10\] datamem.data_ram\[53\]\[3\] _08496_ _08497_
+ VGND VGND VPWR VPWR _08498_ sky130_fd_sc_hd__or4_1
Xhold240 datamem.data_ram\[3\]\[4\] VGND VGND VPWR VPWR net1390 sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 datamem.data_ram\[48\]\[3\] VGND VGND VPWR VPWR net1401 sky130_fd_sc_hd__dlygate4sd3_1
X_29880_ net258 _01615_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[17\]\[11\] sky130_fd_sc_hd__dfxtp_1
Xhold262 datamem.data_ram\[59\]\[1\] VGND VGND VPWR VPWR net1412 sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 datamem.data_ram\[20\]\[4\] VGND VGND VPWR VPWR net1423 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_208_5479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_4450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold284 datamem.data_ram\[45\]\[1\] VGND VGND VPWR VPWR net1434 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_165_4461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28831_ _12918_ VGND VGND VPWR VPWR _04202_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21166_ datamem.data_ram\[10\]\[23\] datamem.data_ram\[11\]\[23\] _06933_ VGND VGND
+ VPWR VPWR _08455_ sky130_fd_sc_hd__mux2_1
X_23727__319 clknet_1_0__leaf__10198_ VGND VGND VPWR VPWR net445 sky130_fd_sc_hd__inv_2
Xhold295 datamem.data_ram\[14\]\[2\] VGND VGND VPWR VPWR net1445 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_591 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20117_ _06752_ _07405_ _07410_ VGND VGND VPWR VPWR _07411_ sky130_fd_sc_hd__or3_1
X_28762_ _12881_ VGND VGND VPWR VPWR _04170_ sky130_fd_sc_hd__clkbuf_1
X_25974_ net33 _11289_ VGND VGND VPWR VPWR _11310_ sky130_fd_sc_hd__or2_1
X_21097_ datamem.data_ram\[1\]\[7\] _06946_ _08385_ _07867_ VGND VGND VPWR VPWR _08386_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_161_4358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_4369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27713_ _12153_ net2390 net50 VGND VGND VPWR VPWR _12295_ sky130_fd_sc_hd__mux2_1
X_20048_ datamem.data_ram\[13\]\[26\] _06662_ _07340_ _07341_ VGND VGND VPWR VPWR
+ _07342_ sky130_fd_sc_hd__o211a_1
X_24925_ _10470_ net2865 net91 VGND VGND VPWR VPWR _10681_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28693_ _12741_ net3805 net42 VGND VGND VPWR VPWR _12845_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27644_ _12257_ VGND VGND VPWR VPWR _03676_ sky130_fd_sc_hd__clkbuf_1
X_24856_ _10390_ net3557 net93 VGND VGND VPWR VPWR _10644_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_102 _06917_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_113 _07077_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_124 _07552_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27575_ _12091_ net2640 net82 VGND VGND VPWR VPWR _12221_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_135 _07831_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24787_ _10472_ net2461 net94 VGND VGND VPWR VPWR _10606_ sky130_fd_sc_hd__mux2_1
XANTENNA_146 _07863_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21999_ _09227_ net104 VGND VGND VPWR VPWR _09229_ sky130_fd_sc_hd__nor2_8
XTAP_TAPCELL_ROW_120_3365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_157 _08464_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29314_ clknet_leaf_0_clk _01049_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD1E\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_212_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26526_ _10073_ _11604_ _11605_ net1585 VGND VGND VPWR VPWR _03210_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_120_3387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_168 _08693_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_179 _08966_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__10126_ _10126_ VGND VGND VPWR VPWR clknet_0__10126_ sky130_fd_sc_hd__clkbuf_16
X_29245_ _09235_ net3177 _13141_ VGND VGND VPWR VPWR _13143_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26457_ _11535_ rvcpu.ALUResultE\[24\] _11288_ VGND VGND VPWR VPWR _11583_ sky130_fd_sc_hd__a21o_1
XFILLER_0_193_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16210_ _14458_ VGND VGND VPWR VPWR _01930_ sky130_fd_sc_hd__clkbuf_1
X_25408_ _10076_ _10950_ VGND VGND VPWR VPWR _10959_ sky130_fd_sc_hd__and2_1
XFILLER_0_148_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29176_ _13105_ VGND VGND VPWR VPWR _04360_ sky130_fd_sc_hd__clkbuf_1
X_17190_ _14177_ net2672 _04851_ VGND VGND VPWR VPWR _04854_ sky130_fd_sc_hd__mux2_1
X_26388_ _11533_ VGND VGND VPWR VPWR _11534_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28127_ _12529_ VGND VGND VPWR VPWR _03887_ sky130_fd_sc_hd__clkbuf_1
X_16141_ _14413_ VGND VGND VPWR VPWR _01954_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25339_ _10915_ VGND VGND VPWR VPWR _02713_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_12_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23888__448 clknet_1_1__leaf__10222_ VGND VGND VPWR VPWR net574 sky130_fd_sc_hd__inv_2
XFILLER_0_84_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28058_ _12355_ net3661 _12492_ VGND VGND VPWR VPWR _12493_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_94_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16072_ net2050 _13260_ _14371_ VGND VGND VPWR VPWR _14377_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15023_ _13409_ _13549_ _13557_ _13570_ VGND VGND VPWR VPWR _13571_ sky130_fd_sc_hd__a211o_1
X_27009_ _11829_ _11886_ VGND VGND VPWR VPWR _11891_ sky130_fd_sc_hd__and2_1
X_19900_ datamem.data_ram\[5\]\[17\] _06665_ _07193_ _07194_ VGND VGND VPWR VPWR _07195_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30020_ net382 _01755_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[13\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_19831_ datamem.data_ram\[34\]\[1\] _07000_ _06970_ datamem.data_ram\[37\]\[1\] VGND
+ VGND VPWR VPWR _07126_ sky130_fd_sc_hd__a22o_1
XFILLER_0_208_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19762_ datamem.data_ram\[49\]\[25\] _06658_ _07053_ _07056_ VGND VGND VPWR VPWR
+ _07057_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_53_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16974_ net3824 _14457_ _04731_ VGND VGND VPWR VPWR _04739_ sky130_fd_sc_hd__mux2_1
X_18713_ _06062_ _06065_ VGND VGND VPWR VPWR _06066_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15925_ _14298_ VGND VGND VPWR VPWR _02063_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_223_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19693_ _06931_ VGND VGND VPWR VPWR _06989_ sky130_fd_sc_hd__buf_4
X_31971_ clknet_leaf_130_clk _03393_ VGND VGND VPWR VPWR datamem.data_ram\[54\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_56 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18644_ _05997_ _05406_ VGND VGND VPWR VPWR _06000_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30922_ clknet_leaf_216_clk _02657_ VGND VGND VPWR VPWR datamem.data_ram\[40\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_15856_ _14260_ VGND VGND VPWR VPWR _02094_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_203_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_189_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14807_ _13358_ _13359_ VGND VGND VPWR VPWR _13360_ sky130_fd_sc_hd__nand2_2
XFILLER_0_203_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30853_ clknet_leaf_154_clk _02588_ VGND VGND VPWR VPWR datamem.data_ram\[43\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18575_ _05588_ _05910_ _05591_ _05654_ VGND VGND VPWR VPWR _05934_ sky130_fd_sc_hd__a31o_1
X_15787_ _14223_ VGND VGND VPWR VPWR _02134_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14738_ _13283_ VGND VGND VPWR VPWR _13291_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_146_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17526_ _05009_ VGND VGND VPWR VPWR _05032_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_87_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30784_ clknet_leaf_155_clk _02519_ VGND VGND VPWR VPWR datamem.data_ram\[46\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32523_ clknet_leaf_247_clk _03945_ VGND VGND VPWR VPWR datamem.data_ram\[24\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_17457_ _04995_ VGND VGND VPWR VPWR _01312_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_172_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14669_ _13236_ VGND VGND VPWR VPWR _03186_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_229_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16408_ net1896 _14438_ _14561_ VGND VGND VPWR VPWR _14570_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32454_ clknet_leaf_250_clk _03876_ VGND VGND VPWR VPWR datamem.data_ram\[27\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_17388_ _14170_ net3423 _04949_ VGND VGND VPWR VPWR _04959_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19127_ _06440_ _06444_ _06443_ VGND VGND VPWR VPWR _06446_ sky130_fd_sc_hd__a21o_1
X_31405_ clknet_leaf_44_clk _03108_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCE\[22\] sky130_fd_sc_hd__dfxtp_1
X_16339_ _14533_ VGND VGND VPWR VPWR _01868_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_171_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32385_ clknet_leaf_231_clk _03807_ VGND VGND VPWR VPWR datamem.data_ram\[29\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23947__501 clknet_1_1__leaf__10228_ VGND VGND VPWR VPWR net627 sky130_fd_sc_hd__inv_2
X_19058_ _06385_ VGND VGND VPWR VPWR rvcpu.dp.lAuiPCE\[5\] sky130_fd_sc_hd__clkbuf_1
X_31336_ clknet_leaf_17_clk _03039_ VGND VGND VPWR VPWR rvcpu.dp.plde.Rs2E\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18009_ _05277_ rvcpu.dp.plde.ImmExtE\[2\] VGND VGND VPWR VPWR _05379_ sky130_fd_sc_hd__or2_1
X_31267_ clknet_leaf_35_clk _02970_ VGND VGND VPWR VPWR rvcpu.dp.plfd.InstrD\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21020_ datamem.data_ram\[53\]\[31\] _06721_ _06654_ datamem.data_ram\[49\]\[31\]
+ _08308_ VGND VGND VPWR VPWR _08309_ sky130_fd_sc_hd__o221a_1
XFILLER_0_168_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30218_ net572 _01953_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[7\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_31198_ clknet_leaf_46_clk _02901_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCPlus4D\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_30149_ net511 _01884_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[0\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_919 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_203_5365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_203_5376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_199_5280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24710_ _10468_ net3220 net59 VGND VGND VPWR VPWR _10563_ sky130_fd_sc_hd__mux2_1
X_21922_ rvcpu.dp.rf.reg_file_arr\[8\]\[28\] rvcpu.dp.rf.reg_file_arr\[10\]\[28\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[28\] rvcpu.dp.rf.reg_file_arr\[11\]\[28\] _08534_
+ _08818_ VGND VGND VPWR VPWR _09156_ sky130_fd_sc_hd__mux4_1
X_25690_ _11086_ _11113_ VGND VGND VPWR VPWR _11117_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_195_5166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_195_5177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24641_ _10524_ VGND VGND VPWR VPWR _02406_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_210_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21853_ _08547_ _09088_ _09090_ _08576_ VGND VGND VPWR VPWR _09091_ sky130_fd_sc_hd__o211a_1
XFILLER_0_194_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20804_ _08091_ _08093_ _07872_ VGND VGND VPWR VPWR _08094_ sky130_fd_sc_hd__a21o_1
X_27360_ _12098_ VGND VGND VPWR VPWR _03551_ sky130_fd_sc_hd__clkbuf_1
X_24572_ _10486_ VGND VGND VPWR VPWR _02375_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_194_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21784_ rvcpu.dp.rf.reg_file_arr\[28\]\[21\] rvcpu.dp.rf.reg_file_arr\[30\]\[21\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[21\] rvcpu.dp.rf.reg_file_arr\[31\]\[21\] _08629_
+ _08683_ VGND VGND VPWR VPWR _09025_ sky130_fd_sc_hd__mux4_1
X_26311_ _11488_ VGND VGND VPWR VPWR _03112_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23523_ _09260_ net3977 _10162_ VGND VGND VPWR VPWR _10170_ sky130_fd_sc_hd__mux2_1
X_27291_ _12036_ net1737 _12053_ _12058_ VGND VGND VPWR VPWR _03522_ sky130_fd_sc_hd__a31o_1
XFILLER_0_203_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20735_ datamem.data_ram\[38\]\[6\] datamem.data_ram\[39\]\[6\] _07828_ VGND VGND
+ VPWR VPWR _08025_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23160__833 clknet_1_1__leaf__10109_ VGND VGND VPWR VPWR net959 sky130_fd_sc_hd__inv_2
XFILLER_0_92_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29030_ _12747_ net4210 _13020_ VGND VGND VPWR VPWR _13027_ sky130_fd_sc_hd__mux2_1
X_26242_ _11457_ VGND VGND VPWR VPWR _11458_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_154_4184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_4195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20666_ datamem.data_ram\[54\]\[29\] _06718_ _06670_ datamem.data_ram\[55\]\[29\]
+ VGND VGND VPWR VPWR _07957_ sky130_fd_sc_hd__o22a_1
XFILLER_0_61_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22405_ _09441_ _09565_ VGND VGND VPWR VPWR _09566_ sky130_fd_sc_hd__nor2_1
X_26173_ _11423_ VGND VGND VPWR VPWR _03039_ sky130_fd_sc_hd__clkbuf_1
X_23385_ _10142_ _09301_ _09361_ VGND VGND VPWR VPWR _10143_ sky130_fd_sc_hd__a21oi_4
X_20597_ _07823_ datamem.data_ram\[3\]\[13\] _07821_ _07887_ VGND VGND VPWR VPWR _07888_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_144_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23275__920 clknet_1_0__leaf__10129_ VGND VGND VPWR VPWR net1046 sky130_fd_sc_hd__inv_2
XFILLER_0_6_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_167_4501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25124_ _10465_ net2432 net87 VGND VGND VPWR VPWR _10794_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_167_4512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22336_ _09442_ _09494_ _09497_ _09499_ VGND VGND VPWR VPWR _09500_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_104_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25055_ _10755_ VGND VGND VPWR VPWR _02589_ sky130_fd_sc_hd__clkbuf_1
X_29932_ net302 _01667_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[16\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_22267_ _09421_ VGND VGND VPWR VPWR _09433_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_163_4409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21218_ _08487_ _08240_ _08490_ VGND VGND VPWR VPWR _04429_ sky130_fd_sc_hd__o21ai_1
X_29863_ net241 _01598_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[18\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_22198_ _09267_ net3433 _09371_ VGND VGND VPWR VPWR _09372_ sky130_fd_sc_hd__mux2_1
X_28814_ _12909_ VGND VGND VPWR VPWR _04194_ sky130_fd_sc_hd__clkbuf_1
X_21149_ datamem.data_ram\[22\]\[23\] _06625_ _06645_ datamem.data_ram\[16\]\[23\]
+ VGND VGND VPWR VPWR _08438_ sky130_fd_sc_hd__o22a_1
X_29794_ net1140 _01529_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[20\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_126_3530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25957_ rvcpu.dp.plfd.InstrD\[0\] _11155_ VGND VGND VPWR VPWR _11301_ sky130_fd_sc_hd__or2_1
X_28745_ _12872_ VGND VGND VPWR VPWR _04162_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_122_3416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15710_ _14177_ net2104 _14173_ VGND VGND VPWR VPWR _14178_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_122_3427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24908_ _10390_ net3994 _10669_ VGND VGND VPWR VPWR _10672_ sky130_fd_sc_hd__mux2_1
X_28676_ _12758_ net2663 _12832_ VGND VGND VPWR VPWR _12836_ sky130_fd_sc_hd__mux2_1
X_16690_ _14154_ net4128 _04587_ VGND VGND VPWR VPWR _04589_ sky130_fd_sc_hd__mux2_1
X_25888_ _11148_ _11260_ _11261_ VGND VGND VPWR VPWR _02916_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_87_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15641_ _14130_ VGND VGND VPWR VPWR _14131_ sky130_fd_sc_hd__clkbuf_4
X_24839_ _10634_ VGND VGND VPWR VPWR _02494_ sky130_fd_sc_hd__clkbuf_1
X_27627_ _12248_ VGND VGND VPWR VPWR _03668_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_197_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_185_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18360_ _05722_ _05652_ rvcpu.dp.plde.ALUControlE\[1\] VGND VGND VPWR VPWR _05725_
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_29_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15572_ _14093_ VGND VGND VPWR VPWR _02219_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27558_ _12153_ net2048 _12206_ VGND VGND VPWR VPWR _12212_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17311_ _04918_ VGND VGND VPWR VPWR _01389_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_25_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18291_ _05283_ _05649_ VGND VGND VPWR VPWR _05656_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27489_ _12136_ net2802 _12169_ VGND VGND VPWR VPWR _12175_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__10109_ _10109_ VGND VGND VPWR VPWR clknet_0__10109_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_154_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17242_ _04881_ VGND VGND VPWR VPWR _01421_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29228_ _09305_ net3627 _13132_ VGND VGND VPWR VPWR _13134_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_96_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23673__270 clknet_1_1__leaf__10193_ VGND VGND VPWR VPWR net396 sky130_fd_sc_hd__inv_2
X_29159_ _13096_ VGND VGND VPWR VPWR _04352_ sky130_fd_sc_hd__clkbuf_1
X_17173_ _14160_ net4170 _04840_ VGND VGND VPWR VPWR _04845_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16124_ _14404_ VGND VGND VPWR VPWR _01962_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32170_ clknet_leaf_229_clk _03592_ VGND VGND VPWR VPWR datamem.data_ram\[37\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31121_ clknet_leaf_109_clk _02856_ VGND VGND VPWR VPWR datamem.data_ram\[35\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_23137__813 clknet_1_1__leaf__10106_ VGND VGND VPWR VPWR net939 sky130_fd_sc_hd__inv_2
X_16055_ net3013 _13235_ _14360_ VGND VGND VPWR VPWR _14368_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_55_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15006_ _13552_ _13553_ _13514_ VGND VGND VPWR VPWR _13554_ sky130_fd_sc_hd__o21a_1
X_31052_ clknet_leaf_186_clk _02787_ VGND VGND VPWR VPWR datamem.data_ram\[9\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30003_ net373 _01738_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[14\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_196_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19814_ datamem.data_ram\[21\]\[9\] _06702_ _06619_ datamem.data_ram\[20\]\[9\] VGND
+ VGND VPWR VPWR _07109_ sky130_fd_sc_hd__o22a_1
XFILLER_0_224_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23330__969 clknet_1_0__leaf__10135_ VGND VGND VPWR VPWR net1095 sky130_fd_sc_hd__inv_2
Xhold1709 datamem.data_ram\[35\]\[21\] VGND VGND VPWR VPWR net2859 sky130_fd_sc_hd__dlygate4sd3_1
X_19745_ datamem.data_ram\[37\]\[25\] _07037_ _07038_ _07039_ VGND VGND VPWR VPWR
+ _07040_ sky130_fd_sc_hd__o211a_1
X_16957_ net2081 _14440_ _04720_ VGND VGND VPWR VPWR _04730_ sky130_fd_sc_hd__mux2_1
XFILLER_0_223_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15908_ _14289_ VGND VGND VPWR VPWR _02071_ sky130_fd_sc_hd__clkbuf_1
X_19676_ datamem.data_ram\[50\]\[0\] _06932_ _06971_ VGND VGND VPWR VPWR _06972_ sky130_fd_sc_hd__a21o_1
X_31954_ clknet_leaf_132_clk _03376_ VGND VGND VPWR VPWR datamem.data_ram\[55\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_16888_ _04693_ VGND VGND VPWR VPWR _01595_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_32 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18627_ _05705_ _05890_ VGND VGND VPWR VPWR _05984_ sky130_fd_sc_hd__nor2_1
X_30905_ clknet_leaf_220_clk _02640_ VGND VGND VPWR VPWR datamem.data_ram\[41\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15839_ _14251_ VGND VGND VPWR VPWR _02102_ sky130_fd_sc_hd__clkbuf_1
X_31885_ clknet_leaf_112_clk _03339_ VGND VGND VPWR VPWR datamem.data_ram\[57\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_539 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30836_ clknet_leaf_135_clk _02571_ VGND VGND VPWR VPWR datamem.data_ram\[44\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_18558_ _05367_ _05729_ _05808_ _05366_ VGND VGND VPWR VPWR _05918_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_190_5052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_190_5063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23756__345 clknet_1_0__leaf__10201_ VGND VGND VPWR VPWR net471 sky130_fd_sc_hd__inv_2
X_17509_ _05023_ VGND VGND VPWR VPWR _01288_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18489_ _05587_ _05664_ VGND VGND VPWR VPWR _05851_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_16_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30767_ clknet_leaf_265_clk _02502_ VGND VGND VPWR VPWR datamem.data_ram\[47\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23224__874 clknet_1_0__leaf__10124_ VGND VGND VPWR VPWR net1000 sky130_fd_sc_hd__inv_2
XANTENNA_13 _06608_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20520_ datamem.data_ram\[24\]\[21\] _06649_ _06621_ datamem.data_ram\[28\]\[21\]
+ _07810_ VGND VGND VPWR VPWR _07811_ sky130_fd_sc_hd__o221a_1
X_32506_ clknet_leaf_239_clk _03928_ VGND VGND VPWR VPWR datamem.data_ram\[24\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_24 _06620_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30698_ clknet_leaf_135_clk _02433_ VGND VGND VPWR VPWR datamem.data_ram\[4\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_35 _06670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_46 _06678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_57 _06704_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20451_ datamem.data_ram\[13\]\[20\] _06768_ _06699_ datamem.data_ram\[9\]\[20\]
+ _07742_ VGND VGND VPWR VPWR _07743_ sky130_fd_sc_hd__o221a_1
XANTENNA_68 _06769_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32437_ clknet_leaf_245_clk _03859_ VGND VGND VPWR VPWR datamem.data_ram\[27\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_79 _06778_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20382_ datamem.data_ram\[54\]\[28\] _06717_ _06695_ datamem.data_ram\[48\]\[28\]
+ VGND VGND VPWR VPWR _07674_ sky130_fd_sc_hd__o22a_1
X_32368_ clknet_leaf_90_clk _03790_ VGND VGND VPWR VPWR datamem.data_ram\[2\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_207_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22121_ rvcpu.dp.plem.WriteDataM\[7\] _08488_ _09293_ VGND VGND VPWR VPWR _09328_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_112_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31319_ clknet_leaf_27_clk _03022_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCPlus4E\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_32299_ clknet_leaf_168_clk _03721_ VGND VGND VPWR VPWR datamem.data_ram\[32\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_205_5405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_205_5416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22052_ _09272_ VGND VGND VPWR VPWR _09273_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_205_5427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Left_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2900 datamem.data_ram\[3\]\[9\] VGND VGND VPWR VPWR net4050 sky130_fd_sc_hd__dlygate4sd3_1
X_21003_ datamem.data_ram\[18\]\[15\] _06639_ VGND VGND VPWR VPWR _08292_ sky130_fd_sc_hd__and2_1
X_26860_ _11679_ _11798_ VGND VGND VPWR VPWR _11800_ sky130_fd_sc_hd__and2_1
Xhold2911 datamem.data_ram\[35\]\[8\] VGND VGND VPWR VPWR net4061 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2922 datamem.data_ram\[25\]\[9\] VGND VGND VPWR VPWR net4072 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_197_5217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2933 rvcpu.dp.rf.reg_file_arr\[29\]\[29\] VGND VGND VPWR VPWR net4083 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_197_5228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25811_ rvcpu.dp.pcreg.q\[19\] _11197_ VGND VGND VPWR VPWR _11200_ sky130_fd_sc_hd__and2_1
Xhold2944 datamem.data_ram\[53\]\[6\] VGND VGND VPWR VPWR net4094 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2955 rvcpu.dp.rf.reg_file_arr\[14\]\[5\] VGND VGND VPWR VPWR net4105 sky130_fd_sc_hd__dlygate4sd3_1
X_26791_ _11689_ _11749_ VGND VGND VPWR VPWR _11758_ sky130_fd_sc_hd__and2_1
Xhold2966 datamem.data_ram\[22\]\[10\] VGND VGND VPWR VPWR net4116 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2977 datamem.data_ram\[26\]\[27\] VGND VGND VPWR VPWR net4127 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_173_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28530_ _12755_ VGND VGND VPWR VPWR _04064_ sky130_fd_sc_hd__clkbuf_1
Xhold2988 datamem.data_ram\[28\]\[30\] VGND VGND VPWR VPWR net4138 sky130_fd_sc_hd__dlygate4sd3_1
X_25742_ _13328_ _11142_ VGND VGND VPWR VPWR _11148_ sky130_fd_sc_hd__nand2_1
Xhold2999 datamem.data_ram\[20\]\[18\] VGND VGND VPWR VPWR net4149 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_214_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22954_ clknet_1_0__leaf__10079_ VGND VGND VPWR VPWR _10080_ sky130_fd_sc_hd__buf_1
XFILLER_0_74_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28461_ _12712_ VGND VGND VPWR VPWR _04038_ sky130_fd_sc_hd__clkbuf_1
X_21905_ rvcpu.dp.rf.reg_file_arr\[12\]\[27\] rvcpu.dp.rf.reg_file_arr\[13\]\[27\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[27\] rvcpu.dp.rf.reg_file_arr\[15\]\[27\] _08549_
+ _08553_ VGND VGND VPWR VPWR _09140_ sky130_fd_sc_hd__mux4_1
X_25673_ _11089_ _11098_ VGND VGND VPWR VPWR _11106_ sky130_fd_sc_hd__and2_1
XFILLER_0_179_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24136__641 clknet_1_0__leaf__10261_ VGND VGND VPWR VPWR net767 sky130_fd_sc_hd__inv_2
Xmax_cap48 _12316_ VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__buf_4
Xmax_cap59 _10561_ VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_4
X_23542__167 clknet_1_1__leaf__10173_ VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__inv_2
XFILLER_0_35_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22885_ _09452_ _10018_ _10020_ _09795_ VGND VGND VPWR VPWR _10021_ sky130_fd_sc_hd__a211o_1
X_27412_ _12125_ net3891 _12126_ VGND VGND VPWR VPWR _12127_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24624_ _10446_ net3683 _10511_ VGND VGND VPWR VPWR _10515_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_194_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_4235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28392_ _12672_ VGND VGND VPWR VPWR _04009_ sky130_fd_sc_hd__clkbuf_1
X_21836_ rvcpu.dp.rf.reg_file_arr\[16\]\[24\] rvcpu.dp.rf.reg_file_arr\[17\]\[24\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[24\] rvcpu.dp.rf.reg_file_arr\[19\]\[24\] _08517_
+ _08519_ VGND VGND VPWR VPWR _09074_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_156_4246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_211_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_214_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27343_ _09313_ VGND VGND VPWR VPWR _12087_ sky130_fd_sc_hd__buf_2
X_24555_ _09321_ VGND VGND VPWR VPWR _10476_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_77_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21767_ rvcpu.dp.rf.reg_file_arr\[24\]\[20\] rvcpu.dp.rf.reg_file_arr\[25\]\[20\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[20\] rvcpu.dp.rf.reg_file_arr\[27\]\[20\] _08548_
+ _08526_ VGND VGND VPWR VPWR _09009_ sky130_fd_sc_hd__mux4_1
XFILLER_0_4_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_1132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20718_ _08003_ _08008_ _07177_ VGND VGND VPWR VPWR _08009_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27274_ _12048_ VGND VGND VPWR VPWR _03515_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_184_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24486_ _10433_ VGND VGND VPWR VPWR _02342_ sky130_fd_sc_hd__clkbuf_1
X_21698_ rvcpu.dp.rf.reg_file_arr\[12\]\[16\] rvcpu.dp.rf.reg_file_arr\[13\]\[16\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[16\] rvcpu.dp.rf.reg_file_arr\[15\]\[16\] _08551_
+ _08555_ VGND VGND VPWR VPWR _08944_ sky130_fd_sc_hd__mux4_1
XFILLER_0_80_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29013_ _12995_ net1655 _13009_ _13017_ VGND VGND VPWR VPWR _04285_ sky130_fd_sc_hd__a31o_1
XFILLER_0_110_1165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26225_ _11450_ VGND VGND VPWR VPWR _03064_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20649_ datamem.data_ram\[27\]\[29\] _06863_ _07936_ _07939_ VGND VGND VPWR VPWR
+ _07940_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_115_3253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_3264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26156_ rvcpu.dp.plfd.InstrD\[14\] _11413_ VGND VGND VPWR VPWR _11415_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_186_4954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25107_ _10724_ net3190 net88 VGND VGND VPWR VPWR _10785_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22319_ _09401_ VGND VGND VPWR VPWR _09484_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_186_4965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26087_ _11369_ net116 VGND VGND VPWR VPWR _11378_ sky130_fd_sc_hd__or2_1
X_29915_ net285 _01650_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[16\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_25038_ _10745_ VGND VGND VPWR VPWR _02582_ sky130_fd_sc_hd__clkbuf_1
X_17860_ _13262_ _05179_ _05180_ net114 VGND VGND VPWR VPWR _05235_ sky130_fd_sc_hd__a31o_1
X_29846_ net224 _01581_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[18\]\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_89_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_89_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16811_ net2756 _14430_ _04648_ VGND VGND VPWR VPWR _04653_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_89_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_3972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17791_ _05175_ _05183_ _05184_ _05186_ VGND VGND VPWR VPWR _05187_ sky130_fd_sc_hd__a31o_1
X_29777_ net1123 _01512_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[20\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_26989_ _10758_ net3949 _11875_ VGND VGND VPWR VPWR _11879_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_145_3983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19530_ datamem.data_ram\[45\]\[24\] _06823_ _06824_ _06825_ VGND VGND VPWR VPWR
+ _06826_ sky130_fd_sc_hd__o211a_1
X_28728_ _12863_ VGND VGND VPWR VPWR _04154_ sky130_fd_sc_hd__clkbuf_1
X_16742_ _04616_ VGND VGND VPWR VPWR _01672_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_85_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_141_3869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23167__839 clknet_1_0__leaf__10110_ VGND VGND VPWR VPWR net965 sky130_fd_sc_hd__inv_2
XFILLER_0_191_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19461_ datamem.data_ram\[56\]\[16\] _06696_ _06686_ datamem.data_ram\[60\]\[16\]
+ _06756_ VGND VGND VPWR VPWR _06757_ sky130_fd_sc_hd__o221a_1
X_16673_ _14137_ net2657 _04576_ VGND VGND VPWR VPWR _04580_ sky130_fd_sc_hd__mux2_1
X_23705__299 clknet_1_1__leaf__10196_ VGND VGND VPWR VPWR net425 sky130_fd_sc_hd__inv_2
X_28659_ _12694_ net3563 _12823_ VGND VGND VPWR VPWR _12827_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_194_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_194_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_159_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18412_ _05775_ _05749_ VGND VGND VPWR VPWR _05776_ sky130_fd_sc_hd__nand2_4
XFILLER_0_186_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15624_ _14120_ VGND VGND VPWR VPWR _02194_ sky130_fd_sc_hd__clkbuf_1
X_31670_ clknet_leaf_68_clk net1324 VGND VGND VPWR VPWR rvcpu.dp.plmw.ALUResultW\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_19392_ _06687_ VGND VGND VPWR VPWR _06688_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_48_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_104_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15555_ _13431_ _13559_ _13780_ _13531_ VGND VGND VPWR VPWR _14079_ sky130_fd_sc_hd__a31o_1
XFILLER_0_201_487 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18343_ _05296_ _05300_ _05665_ VGND VGND VPWR VPWR _05708_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30621_ clknet_leaf_178_clk _02356_ VGND VGND VPWR VPWR datamem.data_ram\[52\]\[8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_16_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18274_ _05636_ _05540_ _05543_ _05638_ VGND VGND VPWR VPWR _05639_ sky130_fd_sc_hd__o22a_1
XFILLER_0_12_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30552_ clknet_leaf_179_clk _02287_ VGND VGND VPWR VPWR datamem.data_ram\[55\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_15486_ _13321_ _13421_ _13495_ _14014_ _13385_ VGND VGND VPWR VPWR _14015_ sky130_fd_sc_hd__o311a_1
XFILLER_0_16_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17225_ _04872_ VGND VGND VPWR VPWR _01429_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30483_ net161 _02218_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[19\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32222_ clknet_leaf_230_clk _03644_ VGND VGND VPWR VPWR datamem.data_ram\[35\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17156_ _14143_ net2642 _04829_ VGND VGND VPWR VPWR _04836_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold806 datamem.data_ram\[4\]\[14\] VGND VGND VPWR VPWR net1956 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold817 rvcpu.dp.rf.reg_file_arr\[8\]\[3\] VGND VGND VPWR VPWR net1967 sky130_fd_sc_hd__dlygate4sd3_1
X_16107_ _14395_ VGND VGND VPWR VPWR _01970_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_220_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32153_ clknet_leaf_161_clk _03575_ VGND VGND VPWR VPWR datamem.data_ram\[38\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold828 rvcpu.dp.rf.reg_file_arr\[5\]\[10\] VGND VGND VPWR VPWR net1978 sky130_fd_sc_hd__dlygate4sd3_1
Xhold839 rvcpu.dp.rf.reg_file_arr\[18\]\[14\] VGND VGND VPWR VPWR net1989 sky130_fd_sc_hd__dlygate4sd3_1
X_17087_ _04799_ VGND VGND VPWR VPWR _01494_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_228_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31104_ clknet_leaf_106_clk _02839_ VGND VGND VPWR VPWR datamem.data_ram\[19\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_16038_ net1973 _13210_ _14349_ VGND VGND VPWR VPWR _14359_ sky130_fd_sc_hd__mux2_1
X_32084_ clknet_leaf_57_clk _03506_ VGND VGND VPWR VPWR datamem.data_ram\[47\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31035_ clknet_leaf_102_clk _02770_ VGND VGND VPWR VPWR datamem.data_ram\[12\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_24005__538 clknet_1_0__leaf__10241_ VGND VGND VPWR VPWR net664 sky130_fd_sc_hd__inv_2
Xhold2207 datamem.data_ram\[25\]\[20\] VGND VGND VPWR VPWR net3357 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2218 rvcpu.dp.rf.reg_file_arr\[1\]\[25\] VGND VGND VPWR VPWR net3368 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2229 datamem.data_ram\[57\]\[26\] VGND VGND VPWR VPWR net3379 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_200_5302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1506 datamem.data_ram\[1\]\[13\] VGND VGND VPWR VPWR net2656 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1517 datamem.data_ram\[37\]\[23\] VGND VGND VPWR VPWR net2667 sky130_fd_sc_hd__dlygate4sd3_1
X_17989_ rvcpu.dp.plde.ImmExtE\[5\] rvcpu.dp.SrcBFW_Mux.y\[5\] _05277_ VGND VGND VPWR
+ VPWR _05359_ sky130_fd_sc_hd__mux2_2
Xhold1528 datamem.data_ram\[15\]\[31\] VGND VGND VPWR VPWR net2678 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1539 datamem.data_ram\[35\]\[11\] VGND VGND VPWR VPWR net2689 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19728_ _06754_ VGND VGND VPWR VPWR _07023_ sky130_fd_sc_hd__buf_8
XFILLER_0_212_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32986_ clknet_leaf_207_clk _04408_ VGND VGND VPWR VPWR datamem.data_ram\[62\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_192_5103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23461__110 clknet_1_0__leaf__10157_ VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_192_5114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31937_ clknet_leaf_123_clk _03359_ VGND VGND VPWR VPWR datamem.data_ram\[59\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_211_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19659_ _06954_ VGND VGND VPWR VPWR _06955_ sky130_fd_sc_hd__buf_4
XFILLER_0_189_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_185_clk clknet_5_22__leaf_clk VGND VGND VPWR VPWR clknet_leaf_185_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_204_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22670_ _09815_ _09816_ _09421_ VGND VGND VPWR VPWR _09817_ sky130_fd_sc_hd__mux2_1
X_31868_ clknet_leaf_123_clk _03322_ VGND VGND VPWR VPWR datamem.data_ram\[63\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_21621_ _08531_ _08870_ _08806_ VGND VGND VPWR VPWR _08871_ sky130_fd_sc_hd__o21a_1
X_30819_ clknet_leaf_173_clk _02554_ VGND VGND VPWR VPWR datamem.data_ram\[45\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31799_ clknet_leaf_98_clk _03253_ VGND VGND VPWR VPWR datamem.data_ram\[46\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_158_Right_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_151_4110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24340_ _10346_ VGND VGND VPWR VPWR _02283_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_151_4121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21552_ _08742_ _08804_ VGND VGND VPWR VPWR _08805_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23005__710 clknet_1_0__leaf__10085_ VGND VGND VPWR VPWR net836 sky130_fd_sc_hd__inv_2
XFILLER_0_74_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_191_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20503_ datamem.data_ram\[40\]\[21\] _06698_ _06636_ datamem.data_ram\[43\]\[21\]
+ _07081_ VGND VGND VPWR VPWR _07794_ sky130_fd_sc_hd__o221a_1
XFILLER_0_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24271_ _10308_ VGND VGND VPWR VPWR _02252_ sky130_fd_sc_hd__clkbuf_1
X_21483_ _08731_ _08735_ _08739_ _08625_ VGND VGND VPWR VPWR _01033_ sky130_fd_sc_hd__o31a_1
X_26010_ rvcpu.dp.plfd.InstrD\[24\] _11329_ _11325_ _11330_ VGND VGND VPWR VPWR _02969_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20434_ datamem.data_ram\[21\]\[12\] _06661_ _06704_ datamem.data_ram\[23\]\[12\]
+ VGND VGND VPWR VPWR _07726_ sky130_fd_sc_hd__o22a_1
XFILLER_0_160_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload260 clknet_leaf_147_clk VGND VGND VPWR VPWR clkload260/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_228_5961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20365_ _07647_ _07648_ _07651_ _07656_ VGND VGND VPWR VPWR _07657_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_228_5972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload271 clknet_leaf_136_clk VGND VGND VPWR VPWR clkload271/Y sky130_fd_sc_hd__clkinv_4
Xclkload282 clknet_1_0__leaf__10248_ VGND VGND VPWR VPWR clkload282/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_149_4061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload293 clknet_1_0__leaf__10203_ VGND VGND VPWR VPWR clkload293/X sky130_fd_sc_hd__clkbuf_8
X_23810__394 clknet_1_0__leaf__10206_ VGND VGND VPWR VPWR net520 sky130_fd_sc_hd__inv_2
X_22104_ _09314_ net3775 _09302_ VGND VGND VPWR VPWR _09315_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_149_4072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27961_ _12434_ VGND VGND VPWR VPWR _03816_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_149_4083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20296_ datamem.data_ram\[11\]\[19\] _06739_ _07585_ _07588_ VGND VGND VPWR VPWR
+ _07589_ sky130_fd_sc_hd__o211a_1
X_23084_ clknet_1_1__leaf__10087_ VGND VGND VPWR VPWR _10102_ sky130_fd_sc_hd__buf_1
XFILLER_0_179_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29700_ net1046 _01435_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[23\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_224_5869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26912_ _11831_ net1634 _11821_ _11832_ VGND VGND VPWR VPWR _03369_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_181_4840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22035_ rvcpu.dp.plem.WriteDataM\[23\] _09220_ VGND VGND VPWR VPWR _09258_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_181_4851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27892_ _11970_ _12394_ VGND VGND VPWR VPWR _12397_ sky130_fd_sc_hd__and2_1
XFILLER_0_179_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2730 datamem.data_ram\[4\]\[25\] VGND VGND VPWR VPWR net3880 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2741 datamem.data_ram\[38\]\[16\] VGND VGND VPWR VPWR net3891 sky130_fd_sc_hd__dlygate4sd3_1
X_29631_ clknet_leaf_148_clk _01366_ VGND VGND VPWR VPWR datamem.data_ram\[5\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_23925__481 clknet_1_0__leaf__10226_ VGND VGND VPWR VPWR net607 sky130_fd_sc_hd__inv_2
XFILLER_0_227_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26843_ _11781_ net1637 _11785_ _11789_ VGND VGND VPWR VPWR _03343_ sky130_fd_sc_hd__a31o_1
Xhold2752 rvcpu.dp.rf.reg_file_arr\[26\]\[23\] VGND VGND VPWR VPWR net3902 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2763 datamem.data_ram\[58\]\[20\] VGND VGND VPWR VPWR net3913 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2774 datamem.data_ram\[61\]\[22\] VGND VGND VPWR VPWR net3924 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2785 rvcpu.dp.rf.reg_file_arr\[22\]\[28\] VGND VGND VPWR VPWR net3935 sky130_fd_sc_hd__dlygate4sd3_1
X_26774_ _07791_ _11725_ _11494_ VGND VGND VPWR VPWR _11747_ sky130_fd_sc_hd__or3_1
XFILLER_0_138_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29562_ net916 _01297_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[27\]\[29\] sky130_fd_sc_hd__dfxtp_1
Xhold2796 rvcpu.dp.rf.reg_file_arr\[23\]\[0\] VGND VGND VPWR VPWR net3946 sky130_fd_sc_hd__dlygate4sd3_1
X_23624__242 clknet_1_1__leaf__10180_ VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_108_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28513_ _12743_ net4445 net43 VGND VGND VPWR VPWR _12744_ sky130_fd_sc_hd__mux2_1
X_25725_ _11136_ VGND VGND VPWR VPWR _02878_ sky130_fd_sc_hd__clkbuf_1
X_22937_ _10066_ VGND VGND VPWR VPWR _10067_ sky130_fd_sc_hd__buf_2
XFILLER_0_168_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_176_clk clknet_5_24__leaf_clk VGND VGND VPWR VPWR clknet_leaf_176_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_86_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29493_ net855 _01228_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[28\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_179_4780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_179_4791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25656_ _10073_ _11094_ _11095_ net1357 VGND VGND VPWR VPWR _02850_ sky130_fd_sc_hd__a22o_1
XFILLER_0_168_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28444_ _12703_ VGND VGND VPWR VPWR _04030_ sky130_fd_sc_hd__clkbuf_1
X_22868_ _10004_ VGND VGND VPWR VPWR _01153_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_195_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_80_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24607_ _10472_ net3806 _10502_ VGND VGND VPWR VPWR _10506_ sky130_fd_sc_hd__mux2_1
Xwire90 _10742_ VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__buf_4
XFILLER_0_183_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_175_4688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28375_ _12363_ net4230 _12659_ VGND VGND VPWR VPWR _12663_ sky130_fd_sc_hd__mux2_1
X_21819_ rvcpu.dp.rf.reg_file_arr\[20\]\[23\] rvcpu.dp.rf.reg_file_arr\[21\]\[23\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[23\] rvcpu.dp.rf.reg_file_arr\[23\]\[23\] _08778_
+ _08825_ VGND VGND VPWR VPWR _09058_ sky130_fd_sc_hd__mux4_1
X_25587_ _11018_ net1468 _11053_ _11056_ VGND VGND VPWR VPWR _02820_ sky130_fd_sc_hd__a31o_1
XFILLER_0_13_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_175_4699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22799_ rvcpu.dp.rf.reg_file_arr\[28\]\[26\] rvcpu.dp.rf.reg_file_arr\[30\]\[26\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[26\] rvcpu.dp.rf.reg_file_arr\[31\]\[26\] _09443_
+ _09453_ VGND VGND VPWR VPWR _09939_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_125_Right_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15340_ _13414_ _13336_ VGND VGND VPWR VPWR _13876_ sky130_fd_sc_hd__nor2_2
XFILLER_0_186_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27326_ _11533_ _12078_ VGND VGND VPWR VPWR _12079_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_117_3304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_3315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24538_ _10464_ VGND VGND VPWR VPWR _02363_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_182_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15271_ _13435_ _13809_ _13353_ VGND VGND VPWR VPWR _13810_ sky130_fd_sc_hd__o21a_1
X_27257_ _10058_ net52 _12042_ net1599 VGND VGND VPWR VPWR _03504_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_191_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24469_ _10424_ VGND VGND VPWR VPWR _02334_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_227_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17010_ net2804 _14424_ _04757_ VGND VGND VPWR VPWR _04759_ sky130_fd_sc_hd__mux2_1
X_26208_ _11369_ _11441_ VGND VGND VPWR VPWR _11443_ sky130_fd_sc_hd__or2_1
XFILLER_0_123_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27188_ _11976_ _11996_ VGND VGND VPWR VPWR _12002_ sky130_fd_sc_hd__and2_1
XFILLER_0_22_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26139_ _11405_ VGND VGND VPWR VPWR _03022_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_100_clk clknet_5_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_100_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18961_ _05698_ _06185_ VGND VGND VPWR VPWR _06298_ sky130_fd_sc_hd__or2_1
XFILLER_0_219_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23785__371 clknet_1_0__leaf__10204_ VGND VGND VPWR VPWR net497 sky130_fd_sc_hd__inv_2
X_17912_ rvcpu.dp.plem.ALUResultM\[30\] _05268_ VGND VGND VPWR VPWR _05285_ sky130_fd_sc_hd__and2_1
X_18892_ _06136_ _05963_ VGND VGND VPWR VPWR _06234_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_37_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17843_ _13231_ rvcpu.dp.plde.RD2E\[15\] _05194_ VGND VGND VPWR VPWR _05223_ sky130_fd_sc_hd__mux2_1
X_29829_ net207 _01564_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[1\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_32840_ clknet_leaf_282_clk _04262_ VGND VGND VPWR VPWR datamem.data_ram\[12\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_17774_ _13277_ _05154_ _05161_ net115 VGND VGND VPWR VPWR _05172_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_221_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14986_ _13475_ _13360_ _13532_ _13533_ VGND VGND VPWR VPWR _13534_ sky130_fd_sc_hd__o22a_1
X_19513_ datamem.data_ram\[50\]\[24\] _06804_ _06806_ datamem.data_ram\[52\]\[24\]
+ _06808_ VGND VGND VPWR VPWR _06809_ sky130_fd_sc_hd__o221a_1
XFILLER_0_117_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16725_ _14189_ net2650 _04598_ VGND VGND VPWR VPWR _04607_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_167_clk clknet_5_24__leaf_clk VGND VGND VPWR VPWR clknet_leaf_167_clk
+ sky130_fd_sc_hd__clkbuf_8
X_32771_ clknet_leaf_213_clk _04193_ VGND VGND VPWR VPWR datamem.data_ram\[14\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_18_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24181__22 clknet_1_0__leaf__10265_ VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_18_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19444_ datamem.data_ram\[44\]\[16\] _06687_ _06700_ datamem.data_ram\[41\]\[16\]
+ VGND VGND VPWR VPWR _06740_ sky130_fd_sc_hd__o22a_1
X_31722_ net171 _03180_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[9\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_46_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16656_ _04570_ VGND VGND VPWR VPWR _01712_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_102_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_102_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15607_ _14111_ VGND VGND VPWR VPWR _02202_ sky130_fd_sc_hd__clkbuf_1
X_31653_ clknet_leaf_66_clk net1581 VGND VGND VPWR VPWR rvcpu.dp.plmw.ALUResultW\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_19375_ _06670_ VGND VGND VPWR VPWR _06671_ sky130_fd_sc_hd__buf_8
XFILLER_0_9_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16587_ _04533_ VGND VGND VPWR VPWR _01752_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_146_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_226_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18326_ _05680_ _05690_ _05676_ VGND VGND VPWR VPWR _05691_ sky130_fd_sc_hd__mux2_2
XFILLER_0_45_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30604_ clknet_leaf_198_clk _02339_ VGND VGND VPWR VPWR datamem.data_ram\[53\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_15538_ _13422_ _13531_ _13616_ VGND VGND VPWR VPWR _14064_ sky130_fd_sc_hd__or3_1
XFILLER_0_151_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31584_ clknet_leaf_52_clk net1185 VGND VGND VPWR VPWR rvcpu.dp.plmw.PCPlus4W\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15469_ _13341_ _13668_ _13858_ VGND VGND VPWR VPWR _13999_ sky130_fd_sc_hd__o21ai_1
X_18257_ rvcpu.dp.plde.RD1E\[20\] _05564_ _05474_ VGND VGND VPWR VPWR _05622_ sky130_fd_sc_hd__o21ai_2
X_30535_ clknet_leaf_196_clk _02270_ VGND VGND VPWR VPWR datamem.data_ram\[55\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17208_ _14195_ net3204 _04828_ VGND VGND VPWR VPWR _04863_ sky130_fd_sc_hd__mux2_1
X_30466_ net144 _02201_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[19\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18188_ _05549_ _05552_ _05542_ _05547_ VGND VGND VPWR VPWR _05553_ sky130_fd_sc_hd__a211o_1
XFILLER_0_29_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold603 datamem.data_ram\[61\]\[2\] VGND VGND VPWR VPWR net1753 sky130_fd_sc_hd__dlygate4sd3_1
X_32205_ clknet_leaf_167_clk _03627_ VGND VGND VPWR VPWR datamem.data_ram\[36\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold614 datamem.data_ram\[0\]\[7\] VGND VGND VPWR VPWR net1764 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17139_ _04826_ VGND VGND VPWR VPWR _01469_ sky130_fd_sc_hd__clkbuf_1
Xhold625 rvcpu.dp.plfd.PCPlus4D\[18\] VGND VGND VPWR VPWR net1775 sky130_fd_sc_hd__dlygate4sd3_1
X_30397_ net735 _02132_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[31\]\[8\] sky130_fd_sc_hd__dfxtp_1
Xhold636 datamem.data_ram\[51\]\[3\] VGND VGND VPWR VPWR net1786 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold647 datamem.data_ram\[51\]\[1\] VGND VGND VPWR VPWR net1797 sky130_fd_sc_hd__dlygate4sd3_1
Xhold658 rvcpu.dp.plfd.PCD\[31\] VGND VGND VPWR VPWR net1808 sky130_fd_sc_hd__dlygate4sd3_1
X_20150_ datamem.data_ram\[53\]\[27\] _06815_ _06670_ datamem.data_ram\[55\]\[27\]
+ VGND VGND VPWR VPWR _07443_ sky130_fd_sc_hd__o22a_1
X_32136_ clknet_leaf_188_clk _03558_ VGND VGND VPWR VPWR datamem.data_ram\[10\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold669 rvcpu.dp.plfd.PCD\[27\] VGND VGND VPWR VPWR net1819 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20081_ datamem.data_ram\[37\]\[10\] _06722_ _06669_ datamem.data_ram\[39\]\[10\]
+ VGND VGND VPWR VPWR _07375_ sky130_fd_sc_hd__o22a_1
X_32067_ clknet_leaf_122_clk _03489_ VGND VGND VPWR VPWR datamem.data_ram\[29\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2004 datamem.data_ram\[1\]\[21\] VGND VGND VPWR VPWR net3154 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23035__736 clknet_1_1__leaf__10089_ VGND VGND VPWR VPWR net862 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_5_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2015 datamem.data_ram\[6\]\[10\] VGND VGND VPWR VPWR net3165 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_176_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2026 datamem.data_ram\[18\]\[19\] VGND VGND VPWR VPWR net3176 sky130_fd_sc_hd__dlygate4sd3_1
X_31018_ clknet_leaf_137_clk _02753_ VGND VGND VPWR VPWR datamem.data_ram\[42\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2037 rvcpu.dp.rf.reg_file_arr\[19\]\[17\] VGND VGND VPWR VPWR net3187 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2048 datamem.data_ram\[31\]\[23\] VGND VGND VPWR VPWR net3198 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1303 datamem.data_ram\[63\]\[31\] VGND VGND VPWR VPWR net2453 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1314 rvcpu.dp.rf.reg_file_arr\[25\]\[1\] VGND VGND VPWR VPWR net2464 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2059 rvcpu.dp.rf.reg_file_arr\[23\]\[14\] VGND VGND VPWR VPWR net3209 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1325 rvcpu.dp.rf.reg_file_arr\[20\]\[20\] VGND VGND VPWR VPWR net2475 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1336 datamem.data_ram\[33\]\[19\] VGND VGND VPWR VPWR net2486 sky130_fd_sc_hd__dlygate4sd3_1
X_23115__793 clknet_1_0__leaf__10104_ VGND VGND VPWR VPWR net919 sky130_fd_sc_hd__inv_2
XFILLER_0_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_227_Right_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_225_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23840_ _10216_ VGND VGND VPWR VPWR _01913_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_174_1232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1347 rvcpu.dp.rf.reg_file_arr\[10\]\[21\] VGND VGND VPWR VPWR net2497 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1358 rvcpu.dp.rf.reg_file_arr\[0\]\[19\] VGND VGND VPWR VPWR net2508 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1369 datamem.data_ram\[34\]\[15\] VGND VGND VPWR VPWR net2519 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_174_1276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_158_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_158_clk
+ sky130_fd_sc_hd__clkbuf_8
X_32969_ clknet_leaf_142_clk _04391_ VGND VGND VPWR VPWR datamem.data_ram\[63\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_509 _13216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20983_ _08270_ _08271_ _06640_ VGND VGND VPWR VPWR _08272_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25510_ _10991_ net1419 _11009_ _11011_ VGND VGND VPWR VPWR _02788_ sky130_fd_sc_hd__a31o_1
XFILLER_0_149_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22722_ _09858_ _09862_ _09866_ _09491_ VGND VGND VPWR VPWR _01145_ sky130_fd_sc_hd__o31a_1
XFILLER_0_95_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_189_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_178_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25441_ _10764_ net2340 _10970_ VGND VGND VPWR VPWR _10977_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0__10090_ _10090_ VGND VGND VPWR VPWR clknet_0__10090_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_94_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22653_ rvcpu.dp.rf.reg_file_arr\[24\]\[18\] rvcpu.dp.rf.reg_file_arr\[25\]\[18\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[18\] rvcpu.dp.rf.reg_file_arr\[27\]\[18\] _09393_
+ _09465_ VGND VGND VPWR VPWR _09801_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_217_5695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28160_ _12355_ net2998 _12546_ VGND VGND VPWR VPWR _12547_ sky130_fd_sc_hd__mux2_1
X_21604_ rvcpu.dp.rf.reg_file_arr\[0\]\[11\] rvcpu.dp.rf.reg_file_arr\[1\]\[11\] rvcpu.dp.rf.reg_file_arr\[2\]\[11\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[11\] _08810_ _08811_ VGND VGND VPWR VPWR _08855_
+ sky130_fd_sc_hd__mux4_1
X_25372_ _10876_ net1681 _10934_ _10937_ VGND VGND VPWR VPWR _02724_ sky130_fd_sc_hd__a31o_1
XFILLER_0_36_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22584_ rvcpu.dp.rf.reg_file_arr\[8\]\[14\] rvcpu.dp.rf.reg_file_arr\[10\]\[14\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[14\] rvcpu.dp.rf.reg_file_arr\[11\]\[14\] _09418_
+ _09485_ VGND VGND VPWR VPWR _09736_ sky130_fd_sc_hd__mux4_2
X_27111_ _11822_ _11953_ VGND VGND VPWR VPWR _11954_ sky130_fd_sc_hd__and2_1
XFILLER_0_152_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24323_ _10326_ net104 VGND VGND VPWR VPWR _10337_ sky130_fd_sc_hd__nor2_8
XFILLER_0_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_211_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_170_4574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28091_ _10141_ _12345_ _12482_ VGND VGND VPWR VPWR _12510_ sky130_fd_sc_hd__a21oi_1
X_21535_ _08542_ _08788_ VGND VGND VPWR VPWR _08789_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_170_4585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27042_ _10402_ _11039_ VGND VGND VPWR VPWR _11911_ sky130_fd_sc_hd__nor2_1
XFILLER_0_160_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24254_ _10299_ VGND VGND VPWR VPWR _02244_ sky130_fd_sc_hd__clkbuf_1
X_21466_ rvcpu.dp.rf.reg_file_arr\[20\]\[5\] rvcpu.dp.rf.reg_file_arr\[21\]\[5\] rvcpu.dp.rf.reg_file_arr\[22\]\[5\]
+ rvcpu.dp.rf.reg_file_arr\[23\]\[5\] _08631_ _08632_ VGND VGND VPWR VPWR _08723_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_161_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_226_5909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23205_ _10123_ VGND VGND VPWR VPWR _01371_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20417_ datamem.data_ram\[55\]\[12\] _06667_ _06684_ datamem.data_ram\[52\]\[12\]
+ VGND VGND VPWR VPWR _07709_ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21397_ rvcpu.dp.rf.reg_file_arr\[28\]\[2\] rvcpu.dp.rf.reg_file_arr\[30\]\[2\] rvcpu.dp.rf.reg_file_arr\[29\]\[2\]
+ rvcpu.dp.rf.reg_file_arr\[31\]\[2\] _08635_ _08637_ VGND VGND VPWR VPWR _08657_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_73_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20348_ datamem.data_ram\[51\]\[4\] _06942_ _06958_ datamem.data_ram\[49\]\[4\] VGND
+ VGND VPWR VPWR _07640_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_1031 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28993_ _12700_ net2286 _12999_ VGND VGND VPWR VPWR _13006_ sky130_fd_sc_hd__mux2_1
XFILLER_0_219_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23468__116 clknet_1_0__leaf__10158_ VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__inv_2
X_27944_ _12424_ VGND VGND VPWR VPWR _03809_ sky130_fd_sc_hd__clkbuf_1
X_23067_ _10095_ VGND VGND VPWR VPWR _01261_ sky130_fd_sc_hd__clkbuf_1
X_20279_ datamem.data_ram\[42\]\[19\] _07023_ _07568_ _07571_ VGND VGND VPWR VPWR
+ _07572_ sky130_fd_sc_hd__o211a_1
XFILLER_0_80_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold3250 datamem.data_ram\[60\]\[19\] VGND VGND VPWR VPWR net4400 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3261 datamem.data_ram\[53\]\[3\] VGND VGND VPWR VPWR net4411 sky130_fd_sc_hd__dlygate4sd3_1
X_22018_ _09244_ net4068 _09232_ VGND VGND VPWR VPWR _09245_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_216_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold3272 rvcpu.dp.plfd.InstrD\[14\] VGND VGND VPWR VPWR net4422 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold3283 datamem.data_ram\[31\]\[29\] VGND VGND VPWR VPWR net4433 sky130_fd_sc_hd__dlygate4sd3_1
X_27875_ _12386_ VGND VGND VPWR VPWR _03778_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_227_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3294 rvcpu.dp.rf.reg_file_arr\[24\]\[0\] VGND VGND VPWR VPWR net4444 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2560 rvcpu.dp.rf.reg_file_arr\[5\]\[28\] VGND VGND VPWR VPWR net3710 sky130_fd_sc_hd__dlygate4sd3_1
X_23548__173 clknet_1_1__leaf__10173_ VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__inv_2
X_29614_ net968 _01349_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[25\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_26826_ _11645_ _11774_ VGND VGND VPWR VPWR _11779_ sky130_fd_sc_hd__and2_1
X_14840_ _13281_ _13288_ VGND VGND VPWR VPWR _13393_ sky130_fd_sc_hd__nand2b_4
Xhold2571 datamem.data_ram\[61\]\[12\] VGND VGND VPWR VPWR net3721 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2582 datamem.data_ram\[56\]\[18\] VGND VGND VPWR VPWR net3732 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2593 datamem.data_ram\[49\]\[30\] VGND VGND VPWR VPWR net3743 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1870 datamem.data_ram\[5\]\[25\] VGND VGND VPWR VPWR net3020 sky130_fd_sc_hd__dlygate4sd3_1
X_14771_ _13320_ _13323_ VGND VGND VPWR VPWR _13324_ sky130_fd_sc_hd__nor2_4
XFILLER_0_187_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1881 rvcpu.dp.rf.reg_file_arr\[21\]\[15\] VGND VGND VPWR VPWR net3031 sky130_fd_sc_hd__dlygate4sd3_1
X_29545_ net899 _01280_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[27\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_26757_ _11725_ _10947_ VGND VGND VPWR VPWR _11738_ sky130_fd_sc_hd__nor2_2
XFILLER_0_216_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_177_4739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_149_clk clknet_5_28__leaf_clk VGND VGND VPWR VPWR clknet_leaf_149_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold1892 datamem.data_ram\[49\]\[31\] VGND VGND VPWR VPWR net3042 sky130_fd_sc_hd__dlygate4sd3_1
X_16510_ net3101 _14470_ _04489_ VGND VGND VPWR VPWR _04493_ sky130_fd_sc_hd__mux2_1
X_25708_ _11127_ VGND VGND VPWR VPWR _02870_ sky130_fd_sc_hd__clkbuf_1
X_26688_ _11684_ _11694_ VGND VGND VPWR VPWR _11698_ sky130_fd_sc_hd__and2_1
X_17490_ _05013_ VGND VGND VPWR VPWR _01297_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29476_ net838 _01211_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[2\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16441_ _04455_ VGND VGND VPWR VPWR _01820_ sky130_fd_sc_hd__clkbuf_1
X_28427_ _09309_ VGND VGND VPWR VPWR _12692_ sky130_fd_sc_hd__clkbuf_2
X_25639_ _11085_ net1721 _11077_ _11088_ VGND VGND VPWR VPWR _02840_ sky130_fd_sc_hd__a31o_1
XFILLER_0_183_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19160_ _06473_ _06474_ VGND VGND VPWR VPWR _06475_ sky130_fd_sc_hd__and2_1
X_16372_ net2210 _14470_ _14547_ VGND VGND VPWR VPWR _14551_ sky130_fd_sc_hd__mux2_1
X_28358_ _12454_ net3742 net95 VGND VGND VPWR VPWR _12654_ sky130_fd_sc_hd__mux2_1
X_15323_ _13857_ _13858_ _13859_ _13501_ VGND VGND VPWR VPWR _13860_ sky130_fd_sc_hd__a31o_1
X_18111_ rvcpu.dp.plde.ImmExtE\[20\] rvcpu.dp.SrcBFW_Mux.y\[20\] _05279_ VGND VGND
+ VPWR VPWR _05478_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_136_3757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27309_ _12061_ net1698 _12065_ _12069_ VGND VGND VPWR VPWR _03529_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_136_3768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19091_ rvcpu.dp.plde.ImmExtE\[10\] rvcpu.dp.plde.PCE\[10\] VGND VGND VPWR VPWR _06414_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_170_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28289_ _12437_ net3502 _12613_ VGND VGND VPWR VPWR _12617_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30320_ net666 _02055_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[4\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15254_ _13373_ _13416_ _13793_ VGND VGND VPWR VPWR _13794_ sky130_fd_sc_hd__or3_1
X_18042_ rvcpu.dp.plde.RD1E\[10\] _05267_ _05271_ _13247_ _05411_ VGND VGND VPWR VPWR
+ _05412_ sky130_fd_sc_hd__a221o_2
XFILLER_0_124_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_227_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30251_ net605 _01986_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[6\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_15185_ _13320_ _13523_ VGND VGND VPWR VPWR _13728_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30182_ net536 _01917_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[8\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_19993_ datamem.data_ram\[0\]\[2\] _06973_ _07283_ _07286_ VGND VGND VPWR VPWR _07287_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_10_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18944_ _05456_ _05527_ _05533_ _05545_ _05768_ _05769_ VGND VGND VPWR VPWR _06282_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_24_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18875_ _06156_ _06217_ _05707_ VGND VGND VPWR VPWR _06218_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17826_ rvcpu.dp.plem.ALUResultM\[24\] _05211_ _05178_ VGND VGND VPWR VPWR _05212_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_207_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32823_ clknet_leaf_212_clk _04245_ VGND VGND VPWR VPWR datamem.data_ram\[12\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_17757_ rvcpu.dp.plmw.RdW\[1\] rvcpu.dp.plde.Rs2E\[1\] VGND VGND VPWR VPWR _05155_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_221_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14969_ _13517_ _13337_ VGND VGND VPWR VPWR _13518_ sky130_fd_sc_hd__nand2_1
XFILLER_0_222_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16708_ _04575_ VGND VGND VPWR VPWR _04598_ sky130_fd_sc_hd__clkbuf_4
X_32754_ clknet_leaf_158_clk _04176_ VGND VGND VPWR VPWR datamem.data_ram\[15\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f__11602_ clknet_0__11602_ VGND VGND VPWR VPWR clknet_1_0__leaf__11602_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_77_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17688_ _05117_ VGND VGND VPWR VPWR _05118_ sky130_fd_sc_hd__clkbuf_4
X_31705_ clknet_leaf_30_clk _03163_ VGND VGND VPWR VPWR rvcpu.dp.pcreg.q\[23\] sky130_fd_sc_hd__dfxtp_1
X_19427_ _06722_ VGND VGND VPWR VPWR _06723_ sky130_fd_sc_hd__clkbuf_8
X_16639_ _04561_ VGND VGND VPWR VPWR _01720_ sky130_fd_sc_hd__clkbuf_1
X_32685_ clknet_leaf_80_clk _04107_ VGND VGND VPWR VPWR datamem.data_ram\[18\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31636_ clknet_leaf_47_clk net1227 VGND VGND VPWR VPWR rvcpu.dp.plmw.lAuiPCW\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19358_ _06653_ VGND VGND VPWR VPWR _06654_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_174_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_174_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18309_ _05380_ VGND VGND VPWR VPWR _05674_ sky130_fd_sc_hd__buf_2
XFILLER_0_29_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31567_ clknet_leaf_62_clk datamem.rd_data_mem\[17\] VGND VGND VPWR VPWR rvcpu.dp.plmw.ReadDataW\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19289_ _06584_ VGND VGND VPWR VPWR _06585_ sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_212_5581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_212_5592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21320_ rvcpu.dp.plde.RdE\[3\] VGND VGND VPWR VPWR _08582_ sky130_fd_sc_hd__inv_2
X_30518_ clknet_leaf_144_clk _02253_ VGND VGND VPWR VPWR datamem.data_ram\[56\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31498_ clknet_leaf_27_clk rvcpu.dp.lAuiPCE\[24\] VGND VGND VPWR VPWR rvcpu.dp.plem.lAuiPCM\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold400 datamem.data_ram\[38\]\[4\] VGND VGND VPWR VPWR net1550 sky130_fd_sc_hd__dlygate4sd3_1
X_21251_ _08512_ VGND VGND VPWR VPWR _08513_ sky130_fd_sc_hd__clkbuf_4
Xhold411 datamem.data_ram\[56\]\[7\] VGND VGND VPWR VPWR net1561 sky130_fd_sc_hd__dlygate4sd3_1
X_30449_ net787 _02184_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[29\]\[28\] sky130_fd_sc_hd__dfxtp_1
Xhold422 datamem.data_ram\[48\]\[5\] VGND VGND VPWR VPWR net1572 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold433 datamem.data_ram\[31\]\[0\] VGND VGND VPWR VPWR net1583 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20202_ datamem.data_ram\[58\]\[11\] _06690_ _07243_ datamem.data_ram\[57\]\[11\]
+ _06600_ VGND VGND VPWR VPWR _07495_ sky130_fd_sc_hd__o221a_1
Xhold444 rvcpu.dp.plfd.PCPlus4D\[5\] VGND VGND VPWR VPWR net1594 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold455 datamem.data_ram\[22\]\[2\] VGND VGND VPWR VPWR net1605 sky130_fd_sc_hd__dlygate4sd3_1
X_21182_ rvcpu.dp.plem.funct3M\[0\] rvcpu.dp.plem.funct3M\[2\] rvcpu.dp.plem.funct3M\[1\]
+ VGND VGND VPWR VPWR _00000_ sky130_fd_sc_hd__o21a_1
XFILLER_0_106_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_198_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold466 datamem.data_ram\[42\]\[1\] VGND VGND VPWR VPWR net1616 sky130_fd_sc_hd__dlygate4sd3_1
Xhold477 rvcpu.dp.plfd.PCD\[9\] VGND VGND VPWR VPWR net1627 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold488 datamem.data_ram\[22\]\[4\] VGND VGND VPWR VPWR net1638 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_86 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32119_ clknet_leaf_84_clk _03541_ VGND VGND VPWR VPWR datamem.data_ram\[0\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20133_ _06777_ _07418_ _07420_ _07425_ VGND VGND VPWR VPWR _07426_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_221_5806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold499 datamem.data_ram\[57\]\[2\] VGND VGND VPWR VPWR net1649 sky130_fd_sc_hd__dlygate4sd3_1
X_25990_ _08567_ _11315_ _11312_ _11319_ VGND VGND VPWR VPWR _02960_ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_216_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24941_ _10689_ VGND VGND VPWR VPWR _02541_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20064_ datamem.data_ram\[61\]\[26\] _06721_ _06645_ datamem.data_ram\[56\]\[26\]
+ _07357_ VGND VGND VPWR VPWR _07358_ sky130_fd_sc_hd__o221a_1
Xhold1100 rvcpu.dp.rf.reg_file_arr\[12\]\[15\] VGND VGND VPWR VPWR net2250 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1111 rvcpu.dp.rf.reg_file_arr\[6\]\[9\] VGND VGND VPWR VPWR net2261 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1122 datamem.data_ram\[50\]\[15\] VGND VGND VPWR VPWR net2272 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1133 datamem.data_ram\[11\]\[19\] VGND VGND VPWR VPWR net2283 sky130_fd_sc_hd__dlygate4sd3_1
X_24872_ _10652_ VGND VGND VPWR VPWR _02509_ sky130_fd_sc_hd__clkbuf_1
X_27660_ _12266_ VGND VGND VPWR VPWR _03683_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_213_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23996__530 clknet_1_0__leaf__10240_ VGND VGND VPWR VPWR net656 sky130_fd_sc_hd__inv_2
Xhold1144 datamem.data_ram\[37\]\[11\] VGND VGND VPWR VPWR net2294 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1155 datamem.data_ram\[38\]\[31\] VGND VGND VPWR VPWR net2305 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26611_ _11653_ VGND VGND VPWR VPWR _03247_ sky130_fd_sc_hd__clkbuf_1
Xhold1166 rvcpu.dp.rf.reg_file_arr\[27\]\[22\] VGND VGND VPWR VPWR net2316 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27591_ _12229_ VGND VGND VPWR VPWR _03651_ sky130_fd_sc_hd__clkbuf_1
Xhold1177 datamem.data_ram\[29\]\[25\] VGND VGND VPWR VPWR net2327 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1188 datamem.data_ram\[30\]\[24\] VGND VGND VPWR VPWR net2338 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1199 datamem.data_ram\[14\]\[16\] VGND VGND VPWR VPWR net2349 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_306 _14156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_219_5746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_219_5757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26542_ _11047_ _11610_ VGND VGND VPWR VPWR _11615_ sky130_fd_sc_hd__and2_1
XFILLER_0_197_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29330_ clknet_leaf_138_clk _01065_ VGND VGND VPWR VPWR datamem.data_ram\[62\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__10111_ clknet_0__10111_ VGND VGND VPWR VPWR clknet_1_1__leaf__10111_
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_317 _14177_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_200_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_328 _14457_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_339 _14466_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20966_ datamem.data_ram\[38\]\[15\] datamem.data_ram\[39\]\[15\] _06651_ VGND VGND
+ VPWR VPWR _08255_ sky130_fd_sc_hd__mux2_1
X_22705_ rvcpu.dp.rf.reg_file_arr\[16\]\[21\] rvcpu.dp.rf.reg_file_arr\[17\]\[21\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[21\] rvcpu.dp.rf.reg_file_arr\[19\]\[21\] _09445_
+ _09447_ VGND VGND VPWR VPWR _09850_ sky130_fd_sc_hd__mux4_1
XFILLER_0_193_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26473_ _11576_ _11244_ _11522_ _06551_ _11593_ VGND VGND VPWR VPWR _11594_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_172_4614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29261_ _13151_ VGND VGND VPWR VPWR _04399_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_172_4625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20897_ datamem.data_ram\[6\]\[22\] datamem.data_ram\[7\]\[22\] _07836_ VGND VGND
+ VPWR VPWR _08187_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25424_ _10764_ net3682 _10961_ VGND VGND VPWR VPWR _10968_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28212_ _12355_ net3093 net45 VGND VGND VPWR VPWR _12575_ sky130_fd_sc_hd__mux2_1
XFILLER_0_192_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29192_ _09305_ net3719 _13112_ VGND VGND VPWR VPWR _13114_ sky130_fd_sc_hd__mux2_1
X_22636_ _09451_ _09782_ _09784_ _09523_ VGND VGND VPWR VPWR _09785_ sky130_fd_sc_hd__o211a_1
XFILLER_0_119_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_192_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25355_ _10876_ net1713 _10920_ _10926_ VGND VGND VPWR VPWR _02718_ sky130_fd_sc_hd__a31o_1
XFILLER_0_165_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28143_ _12447_ net3756 net73 VGND VGND VPWR VPWR _12538_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22567_ rvcpu.dp.rf.reg_file_arr\[8\]\[13\] rvcpu.dp.rf.reg_file_arr\[10\]\[13\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[13\] rvcpu.dp.rf.reg_file_arr\[11\]\[13\] _09608_
+ _09532_ VGND VGND VPWR VPWR _09720_ sky130_fd_sc_hd__mux4_1
XFILLER_0_64_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_1090 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24306_ _10325_ _10327_ _10269_ VGND VGND VPWR VPWR _10328_ sky130_fd_sc_hd__a21oi_4
X_28074_ _10141_ _12335_ _12482_ VGND VGND VPWR VPWR _12501_ sky130_fd_sc_hd__a21oi_4
X_21518_ rvcpu.dp.rf.reg_file_arr\[12\]\[7\] rvcpu.dp.rf.reg_file_arr\[13\]\[7\] rvcpu.dp.rf.reg_file_arr\[14\]\[7\]
+ rvcpu.dp.rf.reg_file_arr\[15\]\[7\] _08567_ _08570_ VGND VGND VPWR VPWR _08773_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_35_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25286_ _10885_ VGND VGND VPWR VPWR _02690_ sky130_fd_sc_hd__clkbuf_1
X_22498_ rvcpu.dp.rf.reg_file_arr\[20\]\[10\] rvcpu.dp.rf.reg_file_arr\[21\]\[10\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[10\] rvcpu.dp.rf.reg_file_arr\[23\]\[10\] _09385_
+ _09637_ VGND VGND VPWR VPWR _09654_ sky130_fd_sc_hd__mux4_2
XFILLER_0_35_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_3632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27025_ _11825_ _11899_ VGND VGND VPWR VPWR _11901_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_131_3643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24237_ _09273_ net3342 _10288_ VGND VGND VPWR VPWR _10290_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21449_ rvcpu.dp.rf.reg_file_arr\[28\]\[4\] rvcpu.dp.rf.reg_file_arr\[30\]\[4\] rvcpu.dp.rf.reg_file_arr\[29\]\[4\]
+ rvcpu.dp.rf.reg_file_arr\[31\]\[4\] _08635_ _08637_ VGND VGND VPWR VPWR _08707_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_133_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_2_Left_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_1148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_39_Left_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28976_ _10072_ _12989_ VGND VGND VPWR VPWR _12997_ sky130_fd_sc_hd__and2_1
X_16990_ _04747_ VGND VGND VPWR VPWR _01547_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_34_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27927_ _12415_ VGND VGND VPWR VPWR _03801_ sky130_fd_sc_hd__clkbuf_1
X_15941_ _14306_ VGND VGND VPWR VPWR _02055_ sky130_fd_sc_hd__clkbuf_1
X_22992__698 clknet_1_1__leaf__10084_ VGND VGND VPWR VPWR net824 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_129_3583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_3594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3080 datamem.data_ram\[21\]\[27\] VGND VGND VPWR VPWR net4230 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3091 rvcpu.dp.rf.reg_file_arr\[28\]\[28\] VGND VGND VPWR VPWR net4241 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_30_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18660_ _05427_ _05406_ _05425_ VGND VGND VPWR VPWR _06015_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_30_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27858_ _12377_ VGND VGND VPWR VPWR _03770_ sky130_fd_sc_hd__clkbuf_1
X_15872_ _14268_ VGND VGND VPWR VPWR _02086_ sky130_fd_sc_hd__clkbuf_1
Xhold2390 datamem.data_ram\[48\]\[15\] VGND VGND VPWR VPWR net3540 sky130_fd_sc_hd__dlygate4sd3_1
X_17611_ _13269_ net4095 _05068_ VGND VGND VPWR VPWR _05077_ sky130_fd_sc_hd__mux2_1
X_26809_ _11687_ _11762_ VGND VGND VPWR VPWR _11769_ sky130_fd_sc_hd__and2_1
X_14823_ _13375_ _13285_ VGND VGND VPWR VPWR _13376_ sky130_fd_sc_hd__nor2_1
X_18591_ _05822_ _05949_ _05799_ VGND VGND VPWR VPWR _05950_ sky130_fd_sc_hd__mux2_1
XFILLER_0_215_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_204_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27789_ _10598_ _12335_ _12260_ VGND VGND VPWR VPWR _12336_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_8_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17542_ _05040_ VGND VGND VPWR VPWR _01272_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_48_Left_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29528_ clknet_leaf_272_clk _01263_ VGND VGND VPWR VPWR datamem.data_ram\[5\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_14754_ _13306_ VGND VGND VPWR VPWR _13307_ sky130_fd_sc_hd__buf_4
XFILLER_0_153_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17473_ _14187_ net3675 _04996_ VGND VGND VPWR VPWR _05004_ sky130_fd_sc_hd__mux2_1
X_29459_ net821 _01194_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[30\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_14685_ net2057 _13248_ _13245_ VGND VGND VPWR VPWR _13249_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19212_ _06516_ VGND VGND VPWR VPWR _06520_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16424_ _14578_ VGND VGND VPWR VPWR _01828_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_771 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32470_ clknet_leaf_81_clk _03892_ VGND VGND VPWR VPWR datamem.data_ram\[26\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31421_ clknet_leaf_103_clk _03124_ VGND VGND VPWR VPWR datamem.data_ram\[15\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_19143_ _06445_ _06459_ _06449_ VGND VGND VPWR VPWR _06460_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16355_ net2186 _14453_ _14536_ VGND VGND VPWR VPWR _14542_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_229_6020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15306_ _13423_ _13561_ _13657_ _13794_ _13843_ VGND VGND VPWR VPWR _13844_ sky130_fd_sc_hd__o311a_1
X_19074_ _06399_ VGND VGND VPWR VPWR rvcpu.dp.lAuiPCE\[7\] sky130_fd_sc_hd__clkbuf_1
X_31352_ clknet_leaf_17_clk _03055_ VGND VGND VPWR VPWR rvcpu.dp.plde.ImmExtE\[1\]
+ sky130_fd_sc_hd__dfxtp_4
Xclkbuf_1_0__f__10200_ clknet_0__10200_ VGND VGND VPWR VPWR clknet_1_0__leaf__10200_
+ sky130_fd_sc_hd__clkbuf_16
X_16286_ _14505_ VGND VGND VPWR VPWR _01893_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18025_ _05390_ _05392_ _05394_ VGND VGND VPWR VPWR _05395_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_23_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30303_ net649 _02038_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[5\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_15237_ _13776_ VGND VGND VPWR VPWR _13777_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_57_Left_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31283_ clknet_leaf_110_clk _02986_ VGND VGND VPWR VPWR datamem.data_ram\[34\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f__10131_ clknet_0__10131_ VGND VGND VPWR VPWR clknet_1_0__leaf__10131_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_164_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15168_ _13706_ _13708_ _13711_ VGND VGND VPWR VPWR _13712_ sky130_fd_sc_hd__o21ai_1
X_23865__427 clknet_1_1__leaf__10220_ VGND VGND VPWR VPWR net553 sky130_fd_sc_hd__inv_2
X_30234_ net588 _01969_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[7\]\[21\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_58_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30165_ net527 _01900_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[0\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_15099_ _13524_ _13643_ VGND VGND VPWR VPWR _13644_ sky130_fd_sc_hd__nand2_1
X_19976_ datamem.data_ram\[21\]\[18\] _06661_ _06780_ datamem.data_ram\[17\]\[18\]
+ VGND VGND VPWR VPWR _07270_ sky130_fd_sc_hd__o22a_1
XFILLER_0_120_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18927_ _05633_ _05534_ _05531_ VGND VGND VPWR VPWR _06266_ sky130_fd_sc_hd__o21ai_1
X_30096_ net458 _01831_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[11\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_197_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_207_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18858_ _06141_ _06201_ _05706_ VGND VGND VPWR VPWR _06202_ sky130_fd_sc_hd__mux2_1
X_17809_ _05200_ VGND VGND VPWR VPWR rvcpu.dp.SrcBFW_Mux.y\[30\] sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_66_Left_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18789_ _05721_ _05734_ VGND VGND VPWR VPWR _06137_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32806_ clknet_leaf_158_clk _04228_ VGND VGND VPWR VPWR datamem.data_ram\[13\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_20820_ datamem.data_ram\[27\]\[30\] _06940_ _07863_ datamem.data_ram\[29\]\[30\]
+ VGND VGND VPWR VPWR _08110_ sky130_fd_sc_hd__o22a_1
XFILLER_0_82_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_222_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30998_ clknet_leaf_102_clk _02733_ VGND VGND VPWR VPWR datamem.data_ram\[22\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20751_ _06642_ _08038_ _08039_ _08040_ _06615_ VGND VGND VPWR VPWR _08041_ sky130_fd_sc_hd__a32o_1
XFILLER_0_175_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32737_ clknet_leaf_252_clk _04159_ VGND VGND VPWR VPWR datamem.data_ram\[16\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_214_5621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_214_5632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_214_5643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20682_ datamem.data_ram\[35\]\[5\] _06943_ _06993_ datamem.data_ram\[39\]\[5\] _06602_
+ VGND VGND VPWR VPWR _07973_ sky130_fd_sc_hd__a221o_1
X_32668_ clknet_leaf_253_clk _04090_ VGND VGND VPWR VPWR datamem.data_ram\[19\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22421_ rvcpu.dp.rf.reg_file_arr\[24\]\[6\] rvcpu.dp.rf.reg_file_arr\[25\]\[6\] rvcpu.dp.rf.reg_file_arr\[26\]\[6\]
+ rvcpu.dp.rf.reg_file_arr\[27\]\[6\] _09392_ _09394_ VGND VGND VPWR VPWR _09581_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_210_5529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31619_ clknet_leaf_14_clk net1268 VGND VGND VPWR VPWR rvcpu.dp.plmw.RegWriteW sky130_fd_sc_hd__dfxtp_2
XFILLER_0_116_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32599_ clknet_leaf_274_clk _04021_ VGND VGND VPWR VPWR datamem.data_ram\[21\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_190_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25140_ _10570_ _10630_ _10705_ VGND VGND VPWR VPWR _10802_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_32_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22352_ _09511_ _09514_ VGND VGND VPWR VPWR _09515_ sky130_fd_sc_hd__or2_1
XFILLER_0_198_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21303_ _08532_ VGND VGND VPWR VPWR _08565_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_66_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25071_ _09259_ VGND VGND VPWR VPWR _10766_ sky130_fd_sc_hd__buf_2
X_22283_ rvcpu.dp.rf.reg_file_arr\[20\]\[1\] rvcpu.dp.rf.reg_file_arr\[21\]\[1\] rvcpu.dp.rf.reg_file_arr\[22\]\[1\]
+ rvcpu.dp.rf.reg_file_arr\[23\]\[1\] _09445_ _09447_ VGND VGND VPWR VPWR _09448_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_198_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold230 datamem.data_ram\[40\]\[2\] VGND VGND VPWR VPWR net1380 sky130_fd_sc_hd__dlygate4sd3_1
X_21234_ datamem.data_ram\[52\]\[10\] datamem.data_ram\[52\]\[3\] VGND VGND VPWR VPWR
+ _08497_ sky130_fd_sc_hd__nand2_1
Xhold241 datamem.data_ram\[32\]\[2\] VGND VGND VPWR VPWR net1391 sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 datamem.data_ram\[11\]\[0\] VGND VGND VPWR VPWR net1402 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold263 datamem.data_ram\[48\]\[2\] VGND VGND VPWR VPWR net1413 sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 datamem.data_ram\[55\]\[5\] VGND VGND VPWR VPWR net1424 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_165_4451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28830_ _12758_ net3567 _12914_ VGND VGND VPWR VPWR _12918_ sky130_fd_sc_hd__mux2_1
Xhold285 datamem.data_ram\[12\]\[4\] VGND VGND VPWR VPWR net1435 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_165_4462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21165_ datamem.data_ram\[8\]\[23\] datamem.data_ram\[9\]\[23\] _06933_ VGND VGND
+ VPWR VPWR _08454_ sky130_fd_sc_hd__mux2_1
XFILLER_0_229_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold296 datamem.data_ram\[4\]\[0\] VGND VGND VPWR VPWR net1446 sky130_fd_sc_hd__dlygate4sd3_1
X_24063__590 clknet_1_1__leaf__10247_ VGND VGND VPWR VPWR net716 sky130_fd_sc_hd__inv_2
X_20116_ datamem.data_ram\[25\]\[10\] _06657_ _07406_ _07409_ VGND VGND VPWR VPWR
+ _07410_ sky130_fd_sc_hd__o211a_1
X_28761_ _12694_ net2474 _12877_ VGND VGND VPWR VPWR _12881_ sky130_fd_sc_hd__mux2_1
X_21096_ _08383_ _08384_ _07838_ VGND VGND VPWR VPWR _08385_ sky130_fd_sc_hd__mux2_1
X_25973_ net1652 _11302_ _11300_ _11309_ VGND VGND VPWR VPWR _02953_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_161_4348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_4359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27712_ _12294_ VGND VGND VPWR VPWR _03707_ sky130_fd_sc_hd__clkbuf_1
X_24924_ _10680_ VGND VGND VPWR VPWR _02533_ sky130_fd_sc_hd__clkbuf_1
X_20047_ datamem.data_ram\[10\]\[26\] _06609_ _06617_ datamem.data_ram\[12\]\[26\]
+ _06598_ VGND VGND VPWR VPWR _07341_ sky130_fd_sc_hd__o221a_1
X_28692_ _12844_ VGND VGND VPWR VPWR _04137_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_217_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_198_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27643_ _12136_ net2353 _12251_ VGND VGND VPWR VPWR _12257_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24855_ _10643_ VGND VGND VPWR VPWR _02501_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_3480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_103 _06921_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_114 _07153_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_213_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_125 _07635_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27574_ _12220_ VGND VGND VPWR VPWR _03643_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_64_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24786_ _10605_ VGND VGND VPWR VPWR _02470_ sky130_fd_sc_hd__clkbuf_1
X_21998_ _09220_ _09219_ VGND VGND VPWR VPWR _09228_ sky130_fd_sc_hd__nor2_8
X_26512__64 clknet_1_0__leaf__11602_ VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_913 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_136 _07832_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29313_ clknet_leaf_290_clk _01048_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD1E\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_147 _07868_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26525_ _10070_ _11604_ _11605_ net1297 VGND VGND VPWR VPWR _03209_ sky130_fd_sc_hd__a22o_1
XANTENNA_158 _08464_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20949_ _07071_ _08225_ _08238_ _06713_ VGND VGND VPWR VPWR _08239_ sky130_fd_sc_hd__o211a_1
XANTENNA_169 _08693_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_80_clk clknet_5_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_80_clk sky130_fd_sc_hd__clkbuf_8
Xclkbuf_0__10125_ _10125_ VGND VGND VPWR VPWR clknet_0__10125_ sky130_fd_sc_hd__clkbuf_16
X_29244_ _13142_ VGND VGND VPWR VPWR _04391_ sky130_fd_sc_hd__clkbuf_1
X_26456_ net1877 _11573_ _11582_ _11570_ VGND VGND VPWR VPWR _03163_ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25407_ _10954_ net1756 _10949_ _10958_ VGND VGND VPWR VPWR _02738_ sky130_fd_sc_hd__a31o_1
X_22619_ rvcpu.dp.rf.reg_file_arr\[0\]\[16\] rvcpu.dp.rf.reg_file_arr\[1\]\[16\] rvcpu.dp.rf.reg_file_arr\[2\]\[16\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[16\] _09714_ _09585_ VGND VGND VPWR VPWR _09769_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_107_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26387_ _06587_ VGND VGND VPWR VPWR _11533_ sky130_fd_sc_hd__clkbuf_4
X_29175_ _09235_ net3791 net63 VGND VGND VPWR VPWR _13105_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16140_ net2855 _13260_ _14407_ VGND VGND VPWR VPWR _14413_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25338_ _10762_ net3936 _10909_ VGND VGND VPWR VPWR _10915_ sky130_fd_sc_hd__mux2_1
X_28126_ _12430_ net3941 _12528_ VGND VGND VPWR VPWR _12529_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_23_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_228_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_662 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16071_ _14376_ VGND VGND VPWR VPWR _01987_ sky130_fd_sc_hd__clkbuf_1
X_25269_ _10055_ VGND VGND VPWR VPWR _10876_ sky130_fd_sc_hd__clkbuf_4
X_28057_ _10141_ _12325_ _12482_ VGND VGND VPWR VPWR _12492_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_94_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15022_ _13327_ _13564_ _13566_ _13569_ VGND VGND VPWR VPWR _13570_ sky130_fd_sc_hd__a31o_1
X_27008_ _11889_ net1646 _11885_ _11890_ VGND VGND VPWR VPWR _03407_ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19830_ _06993_ VGND VGND VPWR VPWR _07125_ sky130_fd_sc_hd__buf_8
XFILLER_0_31_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19761_ datamem.data_ram\[52\]\[25\] _06687_ _07054_ _07055_ VGND VGND VPWR VPWR
+ _07056_ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16973_ _04738_ VGND VGND VPWR VPWR _01555_ sky130_fd_sc_hd__clkbuf_1
X_28959_ _12986_ VGND VGND VPWR VPWR _04262_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_53_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18712_ _05449_ _05732_ _06063_ _06064_ VGND VGND VPWR VPWR _06065_ sky130_fd_sc_hd__o211a_1
X_15924_ net2124 _13244_ _14297_ VGND VGND VPWR VPWR _14298_ sky130_fd_sc_hd__mux2_1
X_31970_ clknet_leaf_130_clk _03392_ VGND VGND VPWR VPWR datamem.data_ram\[54\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_19692_ _06586_ _06987_ _06583_ _06588_ VGND VGND VPWR VPWR _06988_ sky130_fd_sc_hd__o22a_2
XFILLER_0_217_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18643_ _05997_ _05599_ _05809_ VGND VGND VPWR VPWR _05999_ sky130_fd_sc_hd__o21a_1
X_30921_ clknet_leaf_220_clk _02656_ VGND VGND VPWR VPWR datamem.data_ram\[40\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15855_ net4019 _13248_ _14258_ VGND VGND VPWR VPWR _14260_ sky130_fd_sc_hd__mux2_1
X_14806_ _13289_ _13336_ VGND VGND VPWR VPWR _13359_ sky130_fd_sc_hd__nor2_2
X_18574_ _05910_ _05591_ _05588_ VGND VGND VPWR VPWR _05933_ sky130_fd_sc_hd__a21oi_1
X_30852_ clknet_leaf_194_clk _02587_ VGND VGND VPWR VPWR datamem.data_ram\[43\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_15786_ _14175_ net2725 _14221_ VGND VGND VPWR VPWR _14223_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17525_ _05031_ VGND VGND VPWR VPWR _01280_ sky130_fd_sc_hd__clkbuf_1
X_14737_ _13282_ _13285_ _13289_ VGND VGND VPWR VPWR _13290_ sky130_fd_sc_hd__or3_1
X_30783_ clknet_leaf_191_clk _02518_ VGND VGND VPWR VPWR datamem.data_ram\[46\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_71_clk clknet_5_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_71_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_143_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32522_ clknet_leaf_258_clk _03944_ VGND VGND VPWR VPWR datamem.data_ram\[24\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17456_ _14170_ net3332 _04985_ VGND VGND VPWR VPWR _04995_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14668_ net4201 _13235_ _13214_ VGND VGND VPWR VPWR _13236_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16407_ _14569_ VGND VGND VPWR VPWR _01836_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_171_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32453_ clknet_leaf_254_clk _03875_ VGND VGND VPWR VPWR datamem.data_ram\[27\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17387_ _04958_ VGND VGND VPWR VPWR _01345_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_171_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14599_ rvcpu.dp.plmw.ALUResultW\[30\] rvcpu.dp.plmw.ReadDataW\[30\] rvcpu.dp.plmw.PCPlus4W\[30\]
+ rvcpu.dp.plmw.lAuiPCW\[30\] _13168_ _13170_ VGND VGND VPWR VPWR _13183_ sky130_fd_sc_hd__mux4_2
XFILLER_0_6_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19126_ _06440_ _06443_ _06444_ VGND VGND VPWR VPWR _06445_ sky130_fd_sc_hd__nand3_1
X_31404_ clknet_leaf_44_clk _03107_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCE\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16338_ net2133 _14436_ _14525_ VGND VGND VPWR VPWR _14533_ sky130_fd_sc_hd__mux2_1
X_32384_ clknet_leaf_165_clk _03806_ VGND VGND VPWR VPWR datamem.data_ram\[2\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19057_ _06384_ rvcpu.dp.plde.ImmExtE\[5\] _06355_ VGND VGND VPWR VPWR _06385_ sky130_fd_sc_hd__mux2_1
X_31335_ clknet_leaf_17_clk _03038_ VGND VGND VPWR VPWR rvcpu.dp.plde.Rs2E\[1\] sky130_fd_sc_hd__dfxtp_1
X_16269_ _14496_ VGND VGND VPWR VPWR _01901_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_207_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_334 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18008_ _05374_ _05377_ VGND VGND VPWR VPWR _05378_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31266_ clknet_leaf_35_clk _02969_ VGND VGND VPWR VPWR rvcpu.dp.plfd.InstrD\[24\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_11_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30217_ net571 _01952_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[7\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31197_ clknet_leaf_46_clk _02900_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCPlus4D\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_19959_ _06716_ _07234_ _07239_ _07252_ _06713_ VGND VGND VPWR VPWR _07253_ sky130_fd_sc_hd__o311a_1
X_30148_ net510 _01883_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[0\]\[7\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_74_Left_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_203_5366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_203_5377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_5270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30079_ net441 _01814_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[11\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_199_5281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21921_ _08692_ _09152_ _09154_ VGND VGND VPWR VPWR _09155_ sky130_fd_sc_hd__a21o_1
XFILLER_0_179_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_195_5167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_195_5178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24640_ _10390_ net3662 _10521_ VGND VGND VPWR VPWR _10524_ sky130_fd_sc_hd__mux2_1
X_21852_ _08842_ _09089_ VGND VGND VPWR VPWR _09090_ sky130_fd_sc_hd__or2_1
XFILLER_0_210_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20803_ datamem.data_ram\[48\]\[30\] _06779_ _06707_ datamem.data_ram\[55\]\[30\]
+ _08092_ VGND VGND VPWR VPWR _08093_ sky130_fd_sc_hd__o221a_1
X_24571_ _10446_ net2605 _10482_ VGND VGND VPWR VPWR _10486_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21783_ _09022_ _09023_ _08743_ VGND VGND VPWR VPWR _09024_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_62_clk clknet_5_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_62_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_72_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26310_ net1871 _11478_ VGND VGND VPWR VPWR _11488_ sky130_fd_sc_hd__and2_1
X_23522_ _10169_ VGND VGND VPWR VPWR _01642_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20734_ datamem.data_ram\[34\]\[6\] datamem.data_ram\[35\]\[6\] _07837_ VGND VGND
+ VPWR VPWR _08024_ sky130_fd_sc_hd__mux2_1
X_27290_ _11972_ _12054_ VGND VGND VPWR VPWR _12058_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26241_ rvcpu.dp.plfd.InstrD\[31\] _11371_ VGND VGND VPWR VPWR _11457_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_83_Left_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_4185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20665_ datamem.data_ram\[63\]\[29\] _06784_ _07952_ _07955_ VGND VGND VPWR VPWR
+ _07956_ sky130_fd_sc_hd__o211a_1
XFILLER_0_162_223 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_4196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_774 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22404_ _09442_ _09560_ _09562_ _09564_ VGND VGND VPWR VPWR _09565_ sky130_fd_sc_hd__o2bb2a_1
X_26172_ _09482_ _11362_ VGND VGND VPWR VPWR _11423_ sky130_fd_sc_hd__and2_1
X_23384_ _10141_ VGND VGND VPWR VPWR _10142_ sky130_fd_sc_hd__buf_8
X_20596_ datamem.data_ram\[2\]\[13\] _07826_ VGND VGND VPWR VPWR _07887_ sky130_fd_sc_hd__or2_1
X_25123_ _10520_ _10601_ _10705_ VGND VGND VPWR VPWR _10793_ sky130_fd_sc_hd__a21oi_2
X_22335_ _09422_ _09498_ _09457_ VGND VGND VPWR VPWR _09499_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_167_4502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_4513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25054_ _10754_ net3704 _10752_ VGND VGND VPWR VPWR _10755_ sky130_fd_sc_hd__mux2_1
X_29931_ net301 _01666_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[16\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22266_ rvcpu.dp.rf.reg_file_arr\[8\]\[0\] rvcpu.dp.rf.reg_file_arr\[10\]\[0\] rvcpu.dp.rf.reg_file_arr\[9\]\[0\]
+ rvcpu.dp.rf.reg_file_arr\[11\]\[0\] _09431_ _09386_ VGND VGND VPWR VPWR _09432_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_104_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21217_ _08487_ _07857_ _08490_ VGND VGND VPWR VPWR _04428_ sky130_fd_sc_hd__o21ai_1
X_29862_ net240 _01597_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[18\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_22197_ _09351_ _09269_ _09361_ VGND VGND VPWR VPWR _09371_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_40_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28813_ _12694_ net3796 _12905_ VGND VGND VPWR VPWR _12909_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_92_Left_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21148_ datamem.data_ram\[20\]\[23\] _06684_ VGND VGND VPWR VPWR _08437_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29793_ net1139 _01528_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[20\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_126_3520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_3531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28744_ _12741_ net3498 net41 VGND VGND VPWR VPWR _12872_ sky130_fd_sc_hd__mux2_1
X_21079_ _06622_ _08362_ _08364_ _08367_ _07858_ VGND VGND VPWR VPWR _08368_ sky130_fd_sc_hd__o311a_1
X_25956_ _11146_ VGND VGND VPWR VPWR _11300_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_122_3417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24907_ _10671_ VGND VGND VPWR VPWR _02525_ sky130_fd_sc_hd__clkbuf_1
X_28675_ _12835_ VGND VGND VPWR VPWR _04129_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_122_3428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25887_ _08620_ _08621_ VGND VGND VPWR VPWR _11261_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_87_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23282__925 clknet_1_1__leaf__10131_ VGND VGND VPWR VPWR net1051 sky130_fd_sc_hd__inv_2
X_27626_ _12091_ net2731 net80 VGND VGND VPWR VPWR _12248_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_1046 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15640_ _14128_ _14129_ VGND VGND VPWR VPWR _14130_ sky130_fd_sc_hd__nand2_2
XFILLER_0_186_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24838_ _10444_ net3830 _10631_ VGND VGND VPWR VPWR _10634_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27557_ _12211_ VGND VGND VPWR VPWR _03635_ sky130_fd_sc_hd__clkbuf_1
X_15571_ net2156 _13173_ _14092_ VGND VGND VPWR VPWR _14093_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24769_ _10594_ VGND VGND VPWR VPWR _02464_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_53_clk clknet_5_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_53_clk sky130_fd_sc_hd__clkbuf_8
X_24113__620 clknet_1_0__leaf__10259_ VGND VGND VPWR VPWR net746 sky130_fd_sc_hd__inv_2
X_17310_ net4275 _13225_ _04913_ VGND VGND VPWR VPWR _04918_ sky130_fd_sc_hd__mux2_1
XFILLER_0_189_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18290_ _05654_ VGND VGND VPWR VPWR _05655_ sky130_fd_sc_hd__clkbuf_4
X_27488_ _12174_ VGND VGND VPWR VPWR _03603_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23593__214 clknet_1_1__leaf__10177_ VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__inv_2
XFILLER_0_138_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__10108_ _10108_ VGND VGND VPWR VPWR clknet_0__10108_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_194_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17241_ _14160_ net3225 _04876_ VGND VGND VPWR VPWR _04881_ sky130_fd_sc_hd__mux2_1
X_29227_ _13133_ VGND VGND VPWR VPWR _04383_ sky130_fd_sc_hd__clkbuf_1
X_26439_ net2375 _11542_ _11569_ _11570_ VGND VGND VPWR VPWR _03158_ sky130_fd_sc_hd__o211a_1
XFILLER_0_181_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29158_ _09235_ net3870 _13094_ VGND VGND VPWR VPWR _13096_ sky130_fd_sc_hd__mux2_1
X_17172_ _04844_ VGND VGND VPWR VPWR _01454_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28109_ _12355_ net3951 net74 VGND VGND VPWR VPWR _12520_ sky130_fd_sc_hd__mux2_1
X_16123_ net2021 _13235_ _14396_ VGND VGND VPWR VPWR _14404_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29089_ _13059_ VGND VGND VPWR VPWR _04319_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31120_ clknet_leaf_110_clk _02855_ VGND VGND VPWR VPWR datamem.data_ram\[35\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_963 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16054_ _14367_ VGND VGND VPWR VPWR _01995_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_55_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15005_ _13341_ _13492_ VGND VGND VPWR VPWR _13553_ sky130_fd_sc_hd__nor2_2
XFILLER_0_20_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31051_ clknet_leaf_210_clk _02786_ VGND VGND VPWR VPWR datamem.data_ram\[9\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24188__28 clknet_1_1__leaf__10266_ VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__inv_2
X_30002_ net372 _01737_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[14\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_19813_ datamem.data_ram\[22\]\[9\] _06630_ _06672_ datamem.data_ram\[23\]\[9\] VGND
+ VGND VPWR VPWR _07108_ sky130_fd_sc_hd__o22a_1
X_19744_ datamem.data_ram\[32\]\[25\] _06821_ _06828_ datamem.data_ram\[35\]\[25\]
+ _06733_ VGND VGND VPWR VPWR _07039_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16956_ _04729_ VGND VGND VPWR VPWR _01563_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_205_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15907_ net2034 _13220_ _14286_ VGND VGND VPWR VPWR _14289_ sky130_fd_sc_hd__mux2_1
X_19675_ datamem.data_ram\[54\]\[0\] _06951_ _06958_ datamem.data_ram\[49\]\[0\] VGND
+ VGND VPWR VPWR _06971_ sky130_fd_sc_hd__a22o_1
X_31953_ clknet_leaf_133_clk _03375_ VGND VGND VPWR VPWR datamem.data_ram\[55\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_139_Right_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16887_ net3810 _14438_ _04684_ VGND VGND VPWR VPWR _04693_ sky130_fd_sc_hd__mux2_1
X_18626_ _05696_ _05702_ _05691_ _05879_ _05982_ VGND VGND VPWR VPWR _05983_ sky130_fd_sc_hd__a311o_1
X_30904_ clknet_leaf_223_clk _02639_ VGND VGND VPWR VPWR datamem.data_ram\[41\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15838_ net2026 _13223_ _14247_ VGND VGND VPWR VPWR _14251_ sky130_fd_sc_hd__mux2_1
X_31884_ clknet_leaf_123_clk _03338_ VGND VGND VPWR VPWR datamem.data_ram\[57\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_177_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_177_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30835_ clknet_leaf_134_clk _02570_ VGND VGND VPWR VPWR datamem.data_ram\[44\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_18557_ _05675_ _05915_ _05916_ VGND VGND VPWR VPWR _05917_ sky130_fd_sc_hd__o21a_1
X_15769_ _14158_ net3552 _14210_ VGND VGND VPWR VPWR _14214_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_44_clk clknet_5_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_44_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_190_5053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_190_5064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17508_ _13217_ net2934 _05021_ VGND VGND VPWR VPWR _05023_ sky130_fd_sc_hd__mux2_1
X_18488_ _05669_ _05847_ _05849_ VGND VGND VPWR VPWR _05850_ sky130_fd_sc_hd__a21oi_1
X_30766_ clknet_leaf_172_clk _02501_ VGND VGND VPWR VPWR datamem.data_ram\[47\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_871 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32505_ clknet_leaf_231_clk _03927_ VGND VGND VPWR VPWR datamem.data_ram\[24\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_16_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_14 _06610_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17439_ _04986_ VGND VGND VPWR VPWR _01321_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_184_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_25 _06632_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_30697_ clknet_leaf_152_clk _02432_ VGND VGND VPWR VPWR datamem.data_ram\[4\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23259__905 clknet_1_0__leaf__10128_ VGND VGND VPWR VPWR net1031 sky130_fd_sc_hd__inv_2
XFILLER_0_16_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_36 _06671_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_47 _06680_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20450_ datamem.data_ram\[11\]\[20\] _06730_ _06705_ datamem.data_ram\[15\]\[20\]
+ VGND VGND VPWR VPWR _07742_ sky130_fd_sc_hd__o22a_1
X_32436_ clknet_leaf_246_clk _03858_ VGND VGND VPWR VPWR datamem.data_ram\[27\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_58 _06714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_69 _06769_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19109_ _06407_ _06413_ _06416_ _06422_ _06414_ VGND VGND VPWR VPWR _06430_ sky130_fd_sc_hd__o311ai_4
XFILLER_0_125_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32367_ clknet_leaf_90_clk _03789_ VGND VGND VPWR VPWR datamem.data_ram\[2\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20381_ datamem.data_ram\[59\]\[28\] _06828_ _07669_ _07672_ VGND VGND VPWR VPWR
+ _07673_ sky130_fd_sc_hd__o211a_1
XFILLER_0_179_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_209_5520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22120_ _09327_ VGND VGND VPWR VPWR _01082_ sky130_fd_sc_hd__clkbuf_1
X_31318_ clknet_leaf_27_clk _03021_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCPlus4E\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32298_ clknet_leaf_160_clk _03720_ VGND VGND VPWR VPWR datamem.data_ram\[32\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_205_5406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22051_ rvcpu.dp.plem.WriteDataM\[1\] _09264_ _09265_ rvcpu.dp.plem.WriteDataM\[9\]
+ VGND VGND VPWR VPWR _09272_ sky130_fd_sc_hd__a22o_4
XTAP_TAPCELL_ROW_205_5417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31249_ clknet_leaf_21_clk _02952_ VGND VGND VPWR VPWR rvcpu.dp.plfd.InstrD\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21002_ datamem.data_ram\[23\]\[15\] _06667_ _06616_ datamem.data_ram\[20\]\[15\]
+ _08290_ VGND VGND VPWR VPWR _08291_ sky130_fd_sc_hd__o221a_1
XFILLER_0_220_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2901 rvcpu.dp.rf.reg_file_arr\[31\]\[17\] VGND VGND VPWR VPWR net4051 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2912 rvcpu.dp.rf.reg_file_arr\[15\]\[7\] VGND VGND VPWR VPWR net4062 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2923 rvcpu.dp.rf.reg_file_arr\[0\]\[13\] VGND VGND VPWR VPWR net4073 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2934 datamem.data_ram\[44\]\[27\] VGND VGND VPWR VPWR net4084 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_197_5218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25810_ net1775 _11181_ _11177_ _11199_ VGND VGND VPWR VPWR _02900_ sky130_fd_sc_hd__o211a_1
Xhold2945 rvcpu.dp.rf.reg_file_arr\[28\]\[3\] VGND VGND VPWR VPWR net4095 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_197_5229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26790_ _11753_ net1625 _11748_ _11757_ VGND VGND VPWR VPWR _03322_ sky130_fd_sc_hd__a31o_1
XFILLER_0_195_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2956 datamem.data_ram\[10\]\[26\] VGND VGND VPWR VPWR net4106 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2967 datamem.data_ram\[17\]\[24\] VGND VGND VPWR VPWR net4117 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2978 rvcpu.dp.rf.reg_file_arr\[15\]\[20\] VGND VGND VPWR VPWR net4128 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_173_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2989 datamem.data_ram\[57\]\[20\] VGND VGND VPWR VPWR net4139 sky130_fd_sc_hd__dlygate4sd3_1
X_25741_ _11146_ VGND VGND VPWR VPWR _11147_ sky130_fd_sc_hd__clkbuf_4
X_22953_ clknet_1_0__leaf__10078_ VGND VGND VPWR VPWR _10079_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_3_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_106_Right_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21904_ rvcpu.dp.rf.reg_file_arr\[8\]\[27\] rvcpu.dp.rf.reg_file_arr\[10\]\[27\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[27\] rvcpu.dp.rf.reg_file_arr\[11\]\[27\] _08534_
+ _08818_ VGND VGND VPWR VPWR _09139_ sky130_fd_sc_hd__mux4_1
X_28460_ _12445_ net4347 _12704_ VGND VGND VPWR VPWR _12712_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25672_ _11104_ VGND VGND VPWR VPWR _11105_ sky130_fd_sc_hd__clkbuf_4
X_22884_ _09481_ _10019_ VGND VGND VPWR VPWR _10020_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap49 _12298_ VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__buf_4
XFILLER_0_78_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27411_ _10668_ _10908_ _11713_ VGND VGND VPWR VPWR _12126_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_214_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24623_ _10514_ VGND VGND VPWR VPWR _02398_ sky130_fd_sc_hd__clkbuf_1
X_21835_ _09065_ _09069_ _09073_ _08624_ VGND VGND VPWR VPWR _01051_ sky130_fd_sc_hd__o31a_1
X_28391_ _12435_ net2999 _12669_ VGND VGND VPWR VPWR _12672_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_156_4236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_35_clk clknet_5_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_35_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_156_4247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_210_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24554_ _10475_ VGND VGND VPWR VPWR _02368_ sky130_fd_sc_hd__clkbuf_1
X_27342_ _12086_ VGND VGND VPWR VPWR _03545_ sky130_fd_sc_hd__clkbuf_1
X_21766_ rvcpu.dp.rf.reg_file_arr\[28\]\[20\] rvcpu.dp.rf.reg_file_arr\[30\]\[20\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[20\] rvcpu.dp.rf.reg_file_arr\[31\]\[20\] _08559_
+ _08636_ VGND VGND VPWR VPWR _09008_ sky130_fd_sc_hd__mux4_1
XFILLER_0_182_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20717_ datamem.data_ram\[19\]\[5\] _07137_ _08004_ _08007_ VGND VGND VPWR VPWR _08008_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_4_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24485_ _09310_ datamem.data_ram\[52\]\[26\] _10430_ VGND VGND VPWR VPWR _10433_
+ sky130_fd_sc_hd__mux2_1
X_27273_ _10820_ net3915 _12043_ VGND VGND VPWR VPWR _12048_ sky130_fd_sc_hd__mux2_1
X_21697_ _08511_ _08942_ VGND VGND VPWR VPWR _08943_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29012_ _10072_ _13010_ VGND VGND VPWR VPWR _13017_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_880 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26224_ rvcpu.c.ad.funct7b5 _11371_ _11444_ VGND VGND VPWR VPWR _11450_ sky130_fd_sc_hd__and3_1
XFILLER_0_149_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20648_ datamem.data_ram\[30\]\[29\] _06682_ _07937_ _07938_ VGND VGND VPWR VPWR
+ _07939_ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_3254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_384 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26155_ _11414_ VGND VGND VPWR VPWR _03030_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_3265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20579_ _07860_ _07861_ _07869_ VGND VGND VPWR VPWR _07870_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_150_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25106_ _10520_ _10640_ _10705_ VGND VGND VPWR VPWR _10784_ sky130_fd_sc_hd__a21oi_4
X_22318_ _09400_ VGND VGND VPWR VPWR _09483_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_186_4955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26086_ rvcpu.dp.plfd.InstrD\[6\] rvcpu.dp.plfd.InstrD\[3\] _11376_ rvcpu.dp.plfd.InstrD\[4\]
+ VGND VGND VPWR VPWR _11377_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_132_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_186_4966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29914_ net284 _01649_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[16\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_25037_ _10470_ net3386 net90 VGND VGND VPWR VPWR _10745_ sky130_fd_sc_hd__mux2_1
X_22249_ _09399_ VGND VGND VPWR VPWR _09415_ sky130_fd_sc_hd__buf_4
XFILLER_0_218_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29845_ net223 _01580_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[18\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_1102 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16810_ _04652_ VGND VGND VPWR VPWR _01632_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_89_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17790_ _05185_ _05175_ VGND VGND VPWR VPWR _05186_ sky130_fd_sc_hd__nor2_1
X_29776_ net1122 _01511_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[20\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26988_ _11878_ VGND VGND VPWR VPWR _03399_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_145_3973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28727_ _12758_ net2817 _12859_ VGND VGND VPWR VPWR _12863_ sky130_fd_sc_hd__mux2_1
X_16741_ net4131 _14428_ _04612_ VGND VGND VPWR VPWR _04616_ sky130_fd_sc_hd__mux2_1
X_25939_ net1877 _11290_ _11286_ _11291_ VGND VGND VPWR VPWR _02937_ sky130_fd_sc_hd__o211a_1
XFILLER_0_191_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19460_ datamem.data_ram\[61\]\[16\] _06722_ _06655_ datamem.data_ram\[57\]\[16\]
+ VGND VGND VPWR VPWR _06756_ sky130_fd_sc_hd__o22a_1
XFILLER_0_92_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_451 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16672_ _04579_ VGND VGND VPWR VPWR _01705_ sky130_fd_sc_hd__clkbuf_1
X_28658_ _12826_ VGND VGND VPWR VPWR _04121_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18411_ _05590_ _05370_ VGND VGND VPWR VPWR _05775_ sky130_fd_sc_hd__nor2_4
XFILLER_0_97_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15623_ net4252 _13260_ _14114_ VGND VGND VPWR VPWR _14120_ sky130_fd_sc_hd__mux2_1
X_27609_ _12153_ net2113 net81 VGND VGND VPWR VPWR _12239_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19391_ _06686_ VGND VGND VPWR VPWR _06687_ sky130_fd_sc_hd__buf_6
X_23601__221 clknet_1_1__leaf__10178_ VGND VGND VPWR VPWR net347 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_48_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28589_ _12789_ VGND VGND VPWR VPWR _04089_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_26_clk clknet_5_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_26_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_48_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23208__859 clknet_1_1__leaf__10112_ VGND VGND VPWR VPWR net985 sky130_fd_sc_hd__inv_2
XFILLER_0_16_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_104_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18342_ _05706_ VGND VGND VPWR VPWR _05707_ sky130_fd_sc_hd__clkbuf_4
X_30620_ clknet_leaf_147_clk _02355_ VGND VGND VPWR VPWR datamem.data_ram\[52\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_15554_ _13455_ _14077_ _13442_ VGND VGND VPWR VPWR _14078_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_104_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18273_ _05637_ _05546_ VGND VGND VPWR VPWR _05638_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_44_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30551_ clknet_leaf_182_clk _02286_ VGND VGND VPWR VPWR datamem.data_ram\[55\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_15485_ _13541_ _13560_ _13880_ _13332_ VGND VGND VPWR VPWR _14014_ sky130_fd_sc_hd__a211o_1
XFILLER_0_140_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17224_ _14143_ net2646 _04865_ VGND VGND VPWR VPWR _04872_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30482_ net160 _02217_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[19\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32221_ clknet_leaf_222_clk _03643_ VGND VGND VPWR VPWR datamem.data_ram\[35\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17155_ _04835_ VGND VGND VPWR VPWR _01462_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold807 rvcpu.dp.rf.reg_file_arr\[8\]\[21\] VGND VGND VPWR VPWR net1957 sky130_fd_sc_hd__dlygate4sd3_1
X_16106_ net2044 _13210_ _14385_ VGND VGND VPWR VPWR _14395_ sky130_fd_sc_hd__mux2_1
Xhold818 rvcpu.dp.rf.reg_file_arr\[6\]\[21\] VGND VGND VPWR VPWR net1968 sky130_fd_sc_hd__dlygate4sd3_1
X_32152_ clknet_leaf_208_clk _03574_ VGND VGND VPWR VPWR datamem.data_ram\[38\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_760 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17086_ _14141_ net2458 _04793_ VGND VGND VPWR VPWR _04799_ sky130_fd_sc_hd__mux2_1
Xhold829 datamem.data_ram\[18\]\[9\] VGND VGND VPWR VPWR net1979 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31103_ clknet_leaf_108_clk _02838_ VGND VGND VPWR VPWR datamem.data_ram\[19\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_208_Right_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16037_ _14358_ VGND VGND VPWR VPWR _02003_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_204_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32083_ clknet_leaf_62_clk _03505_ VGND VGND VPWR VPWR datamem.data_ram\[47\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31034_ clknet_leaf_102_clk _02769_ VGND VGND VPWR VPWR datamem.data_ram\[12\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2208 datamem.data_ram\[36\]\[14\] VGND VGND VPWR VPWR net3358 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2219 rvcpu.dp.rf.reg_file_arr\[12\]\[1\] VGND VGND VPWR VPWR net3369 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_200_5303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1507 rvcpu.dp.rf.reg_file_arr\[15\]\[28\] VGND VGND VPWR VPWR net2657 sky130_fd_sc_hd__dlygate4sd3_1
X_17988_ rvcpu.dp.plde.RD1E\[5\] _05266_ _05270_ _13262_ _05357_ VGND VGND VPWR VPWR
+ _05358_ sky130_fd_sc_hd__a221o_4
Xhold1518 datamem.data_ram\[40\]\[11\] VGND VGND VPWR VPWR net2668 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1529 datamem.data_ram\[36\]\[18\] VGND VGND VPWR VPWR net2679 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19727_ datamem.data_ram\[13\]\[25\] _07019_ _07021_ datamem.data_ram\[15\]\[25\]
+ VGND VGND VPWR VPWR _07022_ sky130_fd_sc_hd__o22a_1
X_16939_ net2080 _14420_ _04720_ VGND VGND VPWR VPWR _04721_ sky130_fd_sc_hd__mux2_1
X_32985_ clknet_leaf_206_clk _04407_ VGND VGND VPWR VPWR datamem.data_ram\[62\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_192_5104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31936_ clknet_leaf_111_clk _03358_ VGND VGND VPWR VPWR datamem.data_ram\[59\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_19658_ _06953_ VGND VGND VPWR VPWR _06954_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_192_5115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18609_ _05871_ _05966_ _05799_ VGND VGND VPWR VPWR _05967_ sky130_fd_sc_hd__mux2_2
X_31867_ clknet_leaf_122_clk _03321_ VGND VGND VPWR VPWR datamem.data_ram\[63\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19589_ datamem.data_ram\[43\]\[8\] _06634_ _06881_ _06884_ VGND VGND VPWR VPWR _06885_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_176_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_17_clk clknet_5_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_181_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21620_ rvcpu.dp.rf.reg_file_arr\[28\]\[12\] rvcpu.dp.rf.reg_file_arr\[30\]\[12\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[12\] rvcpu.dp.rf.reg_file_arr\[31\]\[12\] _08533_
+ _08536_ VGND VGND VPWR VPWR _08870_ sky130_fd_sc_hd__mux4_1
XFILLER_0_48_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_622 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30818_ clknet_leaf_180_clk _02553_ VGND VGND VPWR VPWR datamem.data_ram\[45\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_31798_ clknet_leaf_209_clk _03252_ VGND VGND VPWR VPWR datamem.data_ram\[2\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_627 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21551_ rvcpu.dp.rf.reg_file_arr\[24\]\[9\] rvcpu.dp.rf.reg_file_arr\[25\]\[9\] rvcpu.dp.rf.reg_file_arr\[26\]\[9\]
+ rvcpu.dp.rf.reg_file_arr\[27\]\[9\] _08548_ _08526_ VGND VGND VPWR VPWR _08804_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_151_4111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30749_ clknet_leaf_179_clk _02484_ VGND VGND VPWR VPWR datamem.data_ram\[48\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_151_4122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20502_ datamem.data_ram\[46\]\[21\] _06630_ _06701_ datamem.data_ram\[41\]\[21\]
+ VGND VGND VPWR VPWR _07793_ sky130_fd_sc_hd__o22a_1
XFILLER_0_173_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24270_ _09224_ net3939 _10307_ VGND VGND VPWR VPWR _10308_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21482_ _08565_ _08736_ _08738_ _08576_ VGND VGND VPWR VPWR _08739_ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_530 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32419_ clknet_leaf_77_clk _03841_ VGND VGND VPWR VPWR datamem.data_ram\[28\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_20433_ datamem.data_ram\[16\]\[12\] _06646_ _06618_ datamem.data_ram\[20\]\[12\]
+ VGND VGND VPWR VPWR _07725_ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_703 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload250 clknet_leaf_153_clk VGND VGND VPWR VPWR clkload250/Y sky130_fd_sc_hd__clkinv_4
X_20364_ datamem.data_ram\[2\]\[28\] _06692_ _07652_ _07655_ VGND VGND VPWR VPWR _07656_
+ sky130_fd_sc_hd__o211a_1
Xclkload261 clknet_leaf_148_clk VGND VGND VPWR VPWR clkload261/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_228_5962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload272 clknet_leaf_137_clk VGND VGND VPWR VPWR clkload272/Y sky130_fd_sc_hd__inv_6
XFILLER_0_141_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_228_5973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22103_ _09313_ VGND VGND VPWR VPWR _09314_ sky130_fd_sc_hd__buf_2
Xclkload283 clknet_1_1__leaf__10247_ VGND VGND VPWR VPWR clkload283/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_149_4062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27960_ _12433_ net3384 _12431_ VGND VGND VPWR VPWR _12434_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload294 clknet_1_1__leaf__10223_ VGND VGND VPWR VPWR clkload294/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_149_4073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20295_ datamem.data_ram\[10\]\[19\] _06754_ _06742_ _07587_ VGND VGND VPWR VPWR
+ _07588_ sky130_fd_sc_hd__o211a_1
XFILLER_0_80_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26911_ _11803_ _11823_ VGND VGND VPWR VPWR _11832_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_181_4830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22034_ _09257_ VGND VGND VPWR VPWR _01066_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_181_4841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27891_ _12391_ net1755 _12393_ _12396_ VGND VGND VPWR VPWR _03784_ sky130_fd_sc_hd__a31o_1
X_23313__954 clknet_1_1__leaf__10133_ VGND VGND VPWR VPWR net1080 sky130_fd_sc_hd__inv_2
XFILLER_0_41_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_220_1172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29630_ clknet_leaf_142_clk _01365_ VGND VGND VPWR VPWR datamem.data_ram\[5\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2720 datamem.data_ram\[7\]\[17\] VGND VGND VPWR VPWR net3870 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_71_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26842_ _11681_ _11786_ VGND VGND VPWR VPWR _11789_ sky130_fd_sc_hd__and2_1
Xhold2731 datamem.data_ram\[34\]\[12\] VGND VGND VPWR VPWR net3881 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2742 datamem.data_ram\[23\]\[26\] VGND VGND VPWR VPWR net3892 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2753 datamem.data_ram\[38\]\[21\] VGND VGND VPWR VPWR net3903 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2764 datamem.data_ram\[18\]\[16\] VGND VGND VPWR VPWR net3914 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2775 datamem.data_ram\[38\]\[14\] VGND VGND VPWR VPWR net3925 sky130_fd_sc_hd__dlygate4sd3_1
X_29561_ net915 _01296_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[27\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_26773_ _11735_ net1851 _11737_ _11746_ VGND VGND VPWR VPWR _03316_ sky130_fd_sc_hd__a31o_1
Xhold2786 datamem.data_ram\[39\]\[21\] VGND VGND VPWR VPWR net3936 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2797 datamem.data_ram\[48\]\[20\] VGND VGND VPWR VPWR net3947 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_108_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28512_ _09281_ VGND VGND VPWR VPWR _12743_ sky130_fd_sc_hd__clkbuf_2
X_25724_ _10816_ net2917 _11133_ VGND VGND VPWR VPWR _11136_ sky130_fd_sc_hd__mux2_1
X_22936_ rvcpu.dp.plem.WriteDataM\[4\] VGND VGND VPWR VPWR _10066_ sky130_fd_sc_hd__buf_4
X_29492_ net854 _01227_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[2\]\[31\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_179_4781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_179_4792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28443_ _12702_ net3241 _12688_ VGND VGND VPWR VPWR _12703_ sky130_fd_sc_hd__mux2_1
X_25655_ _10070_ _11094_ _11095_ net1312 VGND VGND VPWR VPWR _02849_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_80_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22867_ _09388_ _09995_ _09999_ _10003_ VGND VGND VPWR VPWR _10004_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_80_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23739__330 clknet_1_1__leaf__10199_ VGND VGND VPWR VPWR net456 sky130_fd_sc_hd__inv_2
XFILLER_0_38_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24606_ _10505_ VGND VGND VPWR VPWR _02390_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_195_465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xwire91 _10678_ VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__buf_4
X_21818_ rvcpu.dp.rf.reg_file_arr\[16\]\[23\] rvcpu.dp.rf.reg_file_arr\[17\]\[23\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[23\] rvcpu.dp.rf.reg_file_arr\[19\]\[23\] _08631_
+ _08721_ VGND VGND VPWR VPWR _09057_ sky130_fd_sc_hd__mux4_1
X_28374_ _12662_ VGND VGND VPWR VPWR _04001_ sky130_fd_sc_hd__clkbuf_1
X_25586_ _10405_ _11055_ VGND VGND VPWR VPWR _11056_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_175_4689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22798_ _09936_ _09937_ _09449_ VGND VGND VPWR VPWR _09938_ sky130_fd_sc_hd__mux2_2
XFILLER_0_112_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27325_ _07191_ _10042_ _10044_ VGND VGND VPWR VPWR _12078_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_117_3305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24537_ _10400_ net4389 _10456_ VGND VGND VPWR VPWR _10464_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21749_ _08742_ _08991_ VGND VGND VPWR VPWR _08992_ sky130_fd_sc_hd__or2_1
XFILLER_0_186_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15270_ _13401_ _13451_ VGND VGND VPWR VPWR _13809_ sky130_fd_sc_hd__nor2_1
X_27256_ _10048_ net52 _12042_ net1367 VGND VGND VPWR VPWR _03503_ sky130_fd_sc_hd__a22o_1
X_24468_ _09310_ net4227 _10421_ VGND VGND VPWR VPWR _10424_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_184_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_227_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26207_ _11361_ _11371_ VGND VGND VPWR VPWR _11442_ sky130_fd_sc_hd__and2_1
XFILLER_0_145_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27187_ _11991_ net1430 _11995_ _12001_ VGND VGND VPWR VPWR _03475_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_78_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24399_ _09276_ net2311 _10376_ VGND VGND VPWR VPWR _10379_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26138_ net1892 _11397_ VGND VGND VPWR VPWR _11405_ sky130_fd_sc_hd__and2_1
XFILLER_0_22_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18960_ _05715_ _05699_ _05677_ VGND VGND VPWR VPWR _06297_ sky130_fd_sc_hd__mux2_1
X_26069_ _11364_ VGND VGND VPWR VPWR _03029_ sky130_fd_sc_hd__buf_1
XFILLER_0_131_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_219_820 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17911_ _05283_ VGND VGND VPWR VPWR _05284_ sky130_fd_sc_hd__inv_2
X_18891_ _05694_ _05967_ _05866_ VGND VGND VPWR VPWR _06233_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_37_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17842_ _05222_ VGND VGND VPWR VPWR rvcpu.dp.SrcBFW_Mux.y\[17\] sky130_fd_sc_hd__buf_1
XFILLER_0_20_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29828_ net206 _01563_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[1\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23288__931 clknet_1_1__leaf__10131_ VGND VGND VPWR VPWR net1057 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_7_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17773_ _05158_ _05164_ _05167_ _05170_ VGND VGND VPWR VPWR _05171_ sky130_fd_sc_hd__nor4b_1
X_29759_ net1105 _01494_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[21\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_14985_ _13374_ VGND VGND VPWR VPWR _13533_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_156_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19512_ datamem.data_ram\[48\]\[24\] _06807_ _06726_ datamem.data_ram\[55\]\[24\]
+ VGND VGND VPWR VPWR _06808_ sky130_fd_sc_hd__o22a_1
XFILLER_0_221_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16724_ _04606_ VGND VGND VPWR VPWR _01680_ sky130_fd_sc_hd__clkbuf_1
X_32770_ clknet_leaf_212_clk _04192_ VGND VGND VPWR VPWR datamem.data_ram\[14\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19443_ _06738_ VGND VGND VPWR VPWR _06739_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_18_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31721_ net170 _03179_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[9\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16655_ _14187_ net4003 _04562_ VGND VGND VPWR VPWR _04570_ sky130_fd_sc_hd__mux2_1
XFILLER_0_202_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15606_ net2131 _13235_ _14103_ VGND VGND VPWR VPWR _14111_ sky130_fd_sc_hd__mux2_1
X_31652_ clknet_leaf_67_clk net1293 VGND VGND VPWR VPWR rvcpu.dp.plmw.ALUResultW\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_19374_ _06669_ VGND VGND VPWR VPWR _06670_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_146_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16586_ _14187_ net2153 _04525_ VGND VGND VPWR VPWR _04533_ sky130_fd_sc_hd__mux2_1
XFILLER_0_174_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18325_ _05685_ _05687_ _05689_ VGND VGND VPWR VPWR _05690_ sky130_fd_sc_hd__mux2_1
X_30603_ clknet_leaf_195_clk _02338_ VGND VGND VPWR VPWR datamem.data_ram\[53\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15537_ _13512_ _14061_ _14062_ _13319_ VGND VGND VPWR VPWR _14063_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_85_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31583_ clknet_leaf_65_clk net1163 VGND VGND VPWR VPWR rvcpu.dp.plmw.PCPlus4W\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18256_ rvcpu.dp.plde.RD1E\[21\] _05564_ _05468_ VGND VGND VPWR VPWR _05621_ sky130_fd_sc_hd__o21ai_2
X_30534_ clknet_leaf_218_clk _02269_ VGND VGND VPWR VPWR datamem.data_ram\[55\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_15468_ _13341_ _13302_ _13581_ _13328_ VGND VGND VPWR VPWR _13998_ sky130_fd_sc_hd__or4b_1
XFILLER_0_170_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23491__137 clknet_1_1__leaf__10160_ VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__inv_2
X_17207_ _04862_ VGND VGND VPWR VPWR _01437_ sky130_fd_sc_hd__clkbuf_1
X_18187_ _05551_ _05535_ _05529_ VGND VGND VPWR VPWR _05552_ sky130_fd_sc_hd__a21o_1
X_30465_ net143 _02200_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[19\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_15399_ _13572_ _13925_ _13931_ VGND VGND VPWR VPWR _13932_ sky130_fd_sc_hd__a21o_1
XFILLER_0_170_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_1332 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32204_ clknet_leaf_161_clk _03626_ VGND VGND VPWR VPWR datamem.data_ram\[36\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold604 datamem.data_ram\[62\]\[1\] VGND VGND VPWR VPWR net1754 sky130_fd_sc_hd__dlygate4sd3_1
X_17138_ _14193_ net2918 _04792_ VGND VGND VPWR VPWR _04826_ sky130_fd_sc_hd__mux2_1
Xhold615 rvcpu.dp.plfd.PCPlus4D\[19\] VGND VGND VPWR VPWR net1765 sky130_fd_sc_hd__dlygate4sd3_1
Xhold626 rvcpu.dp.plfd.PCPlus4D\[8\] VGND VGND VPWR VPWR net1776 sky130_fd_sc_hd__dlygate4sd3_1
X_23571__194 clknet_1_0__leaf__10175_ VGND VGND VPWR VPWR net320 sky130_fd_sc_hd__inv_2
XFILLER_0_64_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30396_ net734 _02131_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[31\]\[7\] sky130_fd_sc_hd__dfxtp_1
Xhold637 datamem.data_ram\[54\]\[5\] VGND VGND VPWR VPWR net1787 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_229_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold648 datamem.data_ram\[8\]\[7\] VGND VGND VPWR VPWR net1798 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32135_ clknet_leaf_209_clk _03557_ VGND VGND VPWR VPWR datamem.data_ram\[10\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold659 datamem.data_ram\[36\]\[5\] VGND VGND VPWR VPWR net1809 sky130_fd_sc_hd__dlygate4sd3_1
X_17069_ _04789_ VGND VGND VPWR VPWR _01502_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_6_clk clknet_5_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23909__466 clknet_1_1__leaf__10225_ VGND VGND VPWR VPWR net592 sky130_fd_sc_hd__inv_2
X_32066_ clknet_leaf_122_clk _03488_ VGND VGND VPWR VPWR datamem.data_ram\[29\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_20080_ datamem.data_ram\[34\]\[10\] _06803_ _06805_ datamem.data_ram\[36\]\[10\]
+ _07373_ VGND VGND VPWR VPWR _07374_ sky130_fd_sc_hd__o221a_1
XFILLER_0_0_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2005 rvcpu.dp.rf.reg_file_arr\[25\]\[5\] VGND VGND VPWR VPWR net3155 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2016 rvcpu.dp.rf.reg_file_arr\[12\]\[27\] VGND VGND VPWR VPWR net3166 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2027 datamem.data_ram\[63\]\[17\] VGND VGND VPWR VPWR net3177 sky130_fd_sc_hd__dlygate4sd3_1
X_31017_ clknet_leaf_190_clk _02752_ VGND VGND VPWR VPWR datamem.data_ram\[42\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2038 datamem.data_ram\[49\]\[17\] VGND VGND VPWR VPWR net3188 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_176_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1304 rvcpu.dp.rf.reg_file_arr\[27\]\[0\] VGND VGND VPWR VPWR net2454 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_191_Right_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2049 datamem.data_ram\[56\]\[22\] VGND VGND VPWR VPWR net3199 sky130_fd_sc_hd__dlygate4sd3_1
X_23608__227 clknet_1_1__leaf__10179_ VGND VGND VPWR VPWR net353 sky130_fd_sc_hd__inv_2
Xhold1315 datamem.data_ram\[37\]\[17\] VGND VGND VPWR VPWR net2465 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1326 datamem.data_ram\[59\]\[25\] VGND VGND VPWR VPWR net2476 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_224_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1337 rvcpu.dp.rf.reg_file_arr\[9\]\[6\] VGND VGND VPWR VPWR net2487 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1348 datamem.data_ram\[34\]\[23\] VGND VGND VPWR VPWR net2498 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1359 datamem.data_ram\[33\]\[25\] VGND VGND VPWR VPWR net2509 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_224_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32968_ clknet_leaf_202_clk _04390_ VGND VGND VPWR VPWR datamem.data_ram\[63\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_20982_ datamem.data_ram\[14\]\[15\] datamem.data_ram\[15\]\[15\] _06650_ VGND VGND
+ VPWR VPWR _08271_ sky130_fd_sc_hd__mux2_1
XFILLER_0_178_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_174_1288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22721_ _09476_ _09863_ _09865_ _09474_ VGND VGND VPWR VPWR _09866_ sky130_fd_sc_hd__o211a_1
X_31919_ _04431_ net119 VGND VGND VPWR VPWR datamem.rd_data_mem\[24\] sky130_fd_sc_hd__dlxtn_1
XFILLER_0_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32899_ clknet_leaf_210_clk _04321_ VGND VGND VPWR VPWR datamem.data_ram\[0\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25440_ _10976_ VGND VGND VPWR VPWR _02753_ sky130_fd_sc_hd__clkbuf_1
X_22652_ _09798_ _09799_ _09421_ VGND VGND VPWR VPWR _09800_ sky130_fd_sc_hd__mux2_2
XFILLER_0_177_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_217_5696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21603_ _08795_ _08847_ _08849_ _08853_ _08808_ VGND VGND VPWR VPWR _08854_ sky130_fd_sc_hd__a311o_1
X_25371_ _10405_ _10936_ VGND VGND VPWR VPWR _10937_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22583_ rvcpu.dp.rf.reg_file_arr\[12\]\[14\] rvcpu.dp.rf.reg_file_arr\[13\]\[14\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[14\] rvcpu.dp.rf.reg_file_arr\[15\]\[14\] _09386_
+ _09419_ VGND VGND VPWR VPWR _09735_ sky130_fd_sc_hd__mux4_2
XFILLER_0_1_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27110_ _11109_ _10778_ VGND VGND VPWR VPWR _11953_ sky130_fd_sc_hd__nor2_1
XFILLER_0_164_159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21534_ rvcpu.dp.rf.reg_file_arr\[0\]\[8\] rvcpu.dp.rf.reg_file_arr\[1\]\[8\] rvcpu.dp.rf.reg_file_arr\[2\]\[8\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[8\] _08550_ _08554_ VGND VGND VPWR VPWR _08788_ sky130_fd_sc_hd__mux4_1
X_24322_ _10336_ VGND VGND VPWR VPWR _02275_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_170_4564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28090_ _12509_ VGND VGND VPWR VPWR _03870_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_170_4575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_4586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27041_ _11909_ VGND VGND VPWR VPWR _11910_ sky130_fd_sc_hd__clkbuf_2
X_24253_ _09298_ net2753 _10298_ VGND VGND VPWR VPWR _10299_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21465_ rvcpu.dp.rf.reg_file_arr\[16\]\[5\] rvcpu.dp.rf.reg_file_arr\[17\]\[5\] rvcpu.dp.rf.reg_file_arr\[18\]\[5\]
+ rvcpu.dp.rf.reg_file_arr\[19\]\[5\] _08703_ _08721_ VGND VGND VPWR VPWR _08722_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_65_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_209_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23204_ _09260_ net3979 _10115_ VGND VGND VPWR VPWR _10123_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20416_ datamem.data_ram\[53\]\[12\] _06662_ _07243_ datamem.data_ram\[49\]\[12\]
+ VGND VGND VPWR VPWR _07708_ sky130_fd_sc_hd__o22a_1
X_24184_ clknet_1_0__leaf__10079_ VGND VGND VPWR VPWR _10266_ sky130_fd_sc_hd__buf_1
X_21396_ _08654_ _08655_ _08541_ VGND VGND VPWR VPWR _08656_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20347_ datamem.data_ram\[48\]\[4\] _06990_ _06976_ datamem.data_ram\[52\]\[4\] VGND
+ VGND VPWR VPWR _07639_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_73_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28992_ _13005_ VGND VGND VPWR VPWR _04276_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_73_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23237__885 clknet_1_1__leaf__10126_ VGND VGND VPWR VPWR net1011 sky130_fd_sc_hd__inv_2
XFILLER_0_105_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27943_ _12361_ net3406 _12421_ VGND VGND VPWR VPWR _12424_ sky130_fd_sc_hd__mux2_1
X_23066_ _09273_ net3971 _10093_ VGND VGND VPWR VPWR _10095_ sky130_fd_sc_hd__mux2_1
X_20278_ datamem.data_ram\[43\]\[19\] _06738_ _07570_ _06742_ VGND VGND VPWR VPWR
+ _07571_ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold3240 rvcpu.dp.rf.reg_file_arr\[29\]\[25\] VGND VGND VPWR VPWR net4390 sky130_fd_sc_hd__dlygate4sd3_1
X_22017_ _09243_ VGND VGND VPWR VPWR _09244_ sky130_fd_sc_hd__clkbuf_2
Xhold3251 rvcpu.dp.rf.reg_file_arr\[20\]\[27\] VGND VGND VPWR VPWR net4401 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3262 datamem.data_ram\[27\]\[14\] VGND VGND VPWR VPWR net4412 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3273 datamem.data_ram\[53\]\[9\] VGND VGND VPWR VPWR net4423 sky130_fd_sc_hd__dlygate4sd3_1
X_27874_ _12149_ net2647 net77 VGND VGND VPWR VPWR _12386_ sky130_fd_sc_hd__mux2_1
Xhold3284 rvcpu.dp.rf.reg_file_arr\[13\]\[11\] VGND VGND VPWR VPWR net4434 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1097 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_5_26__f_clk clknet_2_3_0_clk VGND VGND VPWR VPWR clknet_5_26__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_142_3910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3295 datamem.data_ram\[1\]\[12\] VGND VGND VPWR VPWR net4445 sky130_fd_sc_hd__dlygate4sd3_1
X_29613_ net967 _01348_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[25\]\[16\] sky130_fd_sc_hd__dfxtp_1
Xhold2550 datamem.data_ram\[63\]\[13\] VGND VGND VPWR VPWR net3700 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26825_ _11767_ net1665 _11773_ _11778_ VGND VGND VPWR VPWR _03336_ sky130_fd_sc_hd__a31o_1
Xhold2561 datamem.data_ram\[5\]\[24\] VGND VGND VPWR VPWR net3711 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2572 datamem.data_ram\[50\]\[13\] VGND VGND VPWR VPWR net3722 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_106_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2583 rvcpu.dp.rf.reg_file_arr\[27\]\[24\] VGND VGND VPWR VPWR net3733 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2594 datamem.data_ram\[53\]\[7\] VGND VGND VPWR VPWR net3744 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29544_ net898 _01279_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[27\]\[11\] sky130_fd_sc_hd__dfxtp_1
Xhold1860 datamem.data_ram\[30\]\[30\] VGND VGND VPWR VPWR net3010 sky130_fd_sc_hd__dlygate4sd3_1
X_26756_ _11736_ VGND VGND VPWR VPWR _11737_ sky130_fd_sc_hd__buf_2
X_14770_ _13321_ _13322_ VGND VGND VPWR VPWR _13323_ sky130_fd_sc_hd__nor2_4
Xhold1871 rvcpu.dp.rf.reg_file_arr\[23\]\[1\] VGND VGND VPWR VPWR net3021 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1882 datamem.data_ram\[0\]\[8\] VGND VGND VPWR VPWR net3032 sky130_fd_sc_hd__dlygate4sd3_1
X_23968_ clknet_1_1__leaf__10224_ VGND VGND VPWR VPWR _10238_ sky130_fd_sc_hd__buf_1
Xhold1893 datamem.data_ram\[34\]\[17\] VGND VGND VPWR VPWR net3043 sky130_fd_sc_hd__dlygate4sd3_1
X_25707_ _10816_ net2895 _11124_ VGND VGND VPWR VPWR _11127_ sky130_fd_sc_hd__mux2_1
X_22919_ _09299_ _10049_ _10052_ VGND VGND VPWR VPWR _10053_ sky130_fd_sc_hd__and3_2
XFILLER_0_168_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29475_ net837 _01210_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[2\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26687_ _11683_ net1678 _11693_ _11697_ VGND VGND VPWR VPWR _03279_ sky130_fd_sc_hd__a31o_1
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16440_ net2102 _14470_ _04451_ VGND VGND VPWR VPWR _04455_ sky130_fd_sc_hd__mux2_1
X_28426_ _12691_ VGND VGND VPWR VPWR _04024_ sky130_fd_sc_hd__clkbuf_1
X_25638_ _11047_ _11079_ VGND VGND VPWR VPWR _11088_ sky130_fd_sc_hd__and2_1
XFILLER_0_169_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28357_ _12653_ VGND VGND VPWR VPWR _03993_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16371_ _14550_ VGND VGND VPWR VPWR _01853_ sky130_fd_sc_hd__clkbuf_1
X_25569_ _10410_ _11042_ VGND VGND VPWR VPWR _11045_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_699 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18110_ _05477_ VGND VGND VPWR VPWR rvcpu.dp.SrcBFW_Mux.y\[20\] sky130_fd_sc_hd__clkbuf_2
X_27308_ _11970_ _12066_ VGND VGND VPWR VPWR _12069_ sky130_fd_sc_hd__and2_1
X_15322_ _13292_ _13301_ _13510_ VGND VGND VPWR VPWR _13859_ sky130_fd_sc_hd__or3_1
X_19090_ rvcpu.dp.plde.ImmExtE\[10\] rvcpu.dp.plde.PCE\[10\] VGND VGND VPWR VPWR _06413_
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_136_3758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_3769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28288_ _12616_ VGND VGND VPWR VPWR _03961_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18041_ rvcpu.dp.plem.ALUResultM\[10\] _05272_ VGND VGND VPWR VPWR _05411_ sky130_fd_sc_hd__and2_1
X_15253_ _13284_ _13307_ _13289_ _13403_ VGND VGND VPWR VPWR _13793_ sky130_fd_sc_hd__and4_1
X_27239_ _11968_ _12031_ VGND VGND VPWR VPWR _12033_ sky130_fd_sc_hd__and2_1
X_22997__703 clknet_1_1__leaf__10084_ VGND VGND VPWR VPWR net829 sky130_fd_sc_hd__inv_2
XFILLER_0_41_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30250_ net604 _01985_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[6\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_15184_ _13324_ _13489_ _13589_ _13431_ _13429_ VGND VGND VPWR VPWR _13727_ sky130_fd_sc_hd__o221a_1
XFILLER_0_1_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19992_ datamem.data_ram\[3\]\[2\] _06942_ _07285_ _06601_ VGND VGND VPWR VPWR _07286_
+ sky130_fd_sc_hd__a211o_1
X_30181_ net535 _01916_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[8\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18943_ _05549_ _06280_ VGND VGND VPWR VPWR _06281_ sky130_fd_sc_hd__xor2_1
XFILLER_0_120_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_197_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18874_ _05469_ _05475_ _05484_ _05490_ _05666_ _05670_ VGND VGND VPWR VPWR _06217_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_218_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17825_ _13203_ rvcpu.dp.plde.RD2E\[24\] _05196_ VGND VGND VPWR VPWR _05211_ sky130_fd_sc_hd__mux2_1
Xhold1 rvcpu.dp.plem.PCPlus4M\[18\] VGND VGND VPWR VPWR net1151 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_179_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32822_ clknet_leaf_237_clk _04244_ VGND VGND VPWR VPWR datamem.data_ram\[12\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_222_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_206_388 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17756_ _13175_ rvcpu.dp.plde.Rs2E\[3\] _05153_ VGND VGND VPWR VPWR _05154_ sky130_fd_sc_hd__o21a_2
XFILLER_0_222_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14968_ _13292_ VGND VGND VPWR VPWR _13517_ sky130_fd_sc_hd__clkbuf_4
X_16707_ _04597_ VGND VGND VPWR VPWR _01688_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32753_ clknet_leaf_160_clk _04175_ VGND VGND VPWR VPWR datamem.data_ram\[15\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f__11601_ clknet_0__11601_ VGND VGND VPWR VPWR clknet_1_0__leaf__11601_
+ sky130_fd_sc_hd__clkbuf_16
X_17687_ _14129_ _04538_ VGND VGND VPWR VPWR _05117_ sky130_fd_sc_hd__nand2_2
X_14899_ _13449_ _13402_ VGND VGND VPWR VPWR _13450_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31704_ clknet_leaf_29_clk _03162_ VGND VGND VPWR VPWR rvcpu.dp.pcreg.q\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19426_ _06721_ VGND VGND VPWR VPWR _06722_ sky130_fd_sc_hd__buf_6
XFILLER_0_71_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_186_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16638_ _14170_ net2587 _04551_ VGND VGND VPWR VPWR _04561_ sky130_fd_sc_hd__mux2_1
XFILLER_0_175_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32684_ clknet_leaf_79_clk _04106_ VGND VGND VPWR VPWR datamem.data_ram\[18\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31635_ clknet_leaf_48_clk net1246 VGND VGND VPWR VPWR rvcpu.dp.plmw.lAuiPCW\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19357_ _06652_ _06642_ VGND VGND VPWR VPWR _06653_ sky130_fd_sc_hd__nand2_8
XFILLER_0_31_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23342__980 clknet_1_1__leaf__10136_ VGND VGND VPWR VPWR net1106 sky130_fd_sc_hd__inv_2
X_16569_ _14170_ net3363 _04514_ VGND VGND VPWR VPWR _04524_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18308_ _05446_ _05412_ _05441_ _05421_ _05665_ _05670_ VGND VGND VPWR VPWR _05673_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_169_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31566_ clknet_leaf_64_clk datamem.rd_data_mem\[16\] VGND VGND VPWR VPWR rvcpu.dp.plmw.ReadDataW\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_19288_ net1 VGND VGND VPWR VPWR _06584_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_155_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_212_5582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_212_5593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30517_ clknet_leaf_144_clk _02252_ VGND VGND VPWR VPWR datamem.data_ram\[56\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_18239_ rvcpu.dp.plem.ALUResultM\[8\] _05272_ _05267_ rvcpu.dp.plde.RD1E\[8\] _05420_
+ VGND VGND VPWR VPWR _05604_ sky130_fd_sc_hd__a221oi_4
XFILLER_0_115_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31497_ clknet_leaf_29_clk rvcpu.dp.lAuiPCE\[23\] VGND VGND VPWR VPWR rvcpu.dp.plem.lAuiPCM\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21250_ rvcpu.dp.plfd.InstrD\[18\] VGND VGND VPWR VPWR _08512_ sky130_fd_sc_hd__clkbuf_4
Xhold401 datamem.data_ram\[60\]\[7\] VGND VGND VPWR VPWR net1551 sky130_fd_sc_hd__dlygate4sd3_1
X_30448_ net786 _02183_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[29\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold412 datamem.data_ram\[54\]\[4\] VGND VGND VPWR VPWR net1562 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold423 datamem.data_ram\[13\]\[2\] VGND VGND VPWR VPWR net1573 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20201_ datamem.data_ram\[59\]\[11\] _06730_ _06765_ datamem.data_ram\[60\]\[11\]
+ VGND VGND VPWR VPWR _07494_ sky130_fd_sc_hd__o22a_1
Xhold434 datamem.data_ram\[58\]\[4\] VGND VGND VPWR VPWR net1584 sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 datamem.data_ram\[32\]\[7\] VGND VGND VPWR VPWR net1595 sky130_fd_sc_hd__dlygate4sd3_1
X_21181_ _06583_ _08466_ _08467_ _08469_ VGND VGND VPWR VPWR _04444_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_187_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_4010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30379_ net725 _02114_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[3\]\[30\] sky130_fd_sc_hd__dfxtp_1
Xhold456 datamem.data_ram\[29\]\[4\] VGND VGND VPWR VPWR net1606 sky130_fd_sc_hd__dlygate4sd3_1
Xhold467 datamem.data_ram\[58\]\[3\] VGND VGND VPWR VPWR net1617 sky130_fd_sc_hd__dlygate4sd3_1
Xhold478 datamem.data_ram\[23\]\[6\] VGND VGND VPWR VPWR net1628 sky130_fd_sc_hd__dlygate4sd3_1
X_32118_ clknet_leaf_98_clk _03540_ VGND VGND VPWR VPWR datamem.data_ram\[0\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_20132_ _06602_ _07422_ _07424_ VGND VGND VPWR VPWR _07425_ sky130_fd_sc_hd__and3_1
Xhold489 datamem.data_ram\[48\]\[7\] VGND VGND VPWR VPWR net1639 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_221_5807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32049_ clknet_leaf_131_clk _03471_ VGND VGND VPWR VPWR datamem.data_ram\[30\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24940_ _10442_ net2754 _10687_ VGND VGND VPWR VPWR _10689_ sky130_fd_sc_hd__mux2_1
X_20063_ datamem.data_ram\[58\]\[26\] _06608_ VGND VGND VPWR VPWR _07357_ sky130_fd_sc_hd__or2_1
XFILLER_0_176_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1101 rvcpu.dp.rf.reg_file_arr\[1\]\[24\] VGND VGND VPWR VPWR net2251 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1112 rvcpu.dp.rf.reg_file_arr\[27\]\[7\] VGND VGND VPWR VPWR net2262 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1123 rvcpu.dp.rf.reg_file_arr\[19\]\[10\] VGND VGND VPWR VPWR net2273 sky130_fd_sc_hd__dlygate4sd3_1
X_23440__91 clknet_1_0__leaf__10155_ VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__inv_2
XFILLER_0_225_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24871_ _10468_ net3248 net92 VGND VGND VPWR VPWR _10652_ sky130_fd_sc_hd__mux2_1
XFILLER_0_224_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1134 datamem.data_ram\[12\]\[16\] VGND VGND VPWR VPWR net2284 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1145 rvcpu.dp.rf.reg_file_arr\[8\]\[7\] VGND VGND VPWR VPWR net2295 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1156 datamem.data_ram\[60\]\[15\] VGND VGND VPWR VPWR net2306 sky130_fd_sc_hd__dlygate4sd3_1
X_26610_ _10816_ net3213 _11650_ VGND VGND VPWR VPWR _11653_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23822_ clknet_1_1__leaf__10203_ VGND VGND VPWR VPWR _10208_ sky130_fd_sc_hd__buf_1
Xhold1167 rvcpu.dp.rf.reg_file_arr\[7\]\[10\] VGND VGND VPWR VPWR net2317 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27590_ _12134_ net4173 _12224_ VGND VGND VPWR VPWR _12229_ sky130_fd_sc_hd__mux2_1
Xhold1178 rvcpu.dp.rf.reg_file_arr\[13\]\[22\] VGND VGND VPWR VPWR net2328 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1189 datamem.data_ram\[6\]\[22\] VGND VGND VPWR VPWR net2339 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_36_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_307 _14158_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__10110_ clknet_0__10110_ VGND VGND VPWR VPWR clknet_1_1__leaf__10110_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_219_5747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26541_ _11517_ net1457 _11608_ _11614_ VGND VGND VPWR VPWR _03216_ sky130_fd_sc_hd__a31o_1
XANTENNA_318 _14185_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_219_5758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20965_ _08242_ _08247_ _08253_ VGND VGND VPWR VPWR _08254_ sky130_fd_sc_hd__a21o_1
XANTENNA_329 _14457_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22704_ _09849_ VGND VGND VPWR VPWR _01144_ sky130_fd_sc_hd__clkbuf_1
X_29260_ _09266_ net4317 _13150_ VGND VGND VPWR VPWR _13151_ sky130_fd_sc_hd__mux2_1
X_26472_ _11535_ rvcpu.ALUResultE\[29\] _11288_ VGND VGND VPWR VPWR _11593_ sky130_fd_sc_hd__a21o_1
XFILLER_0_32_1008 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20896_ datamem.data_ram\[4\]\[22\] datamem.data_ram\[5\]\[22\] _07836_ VGND VGND
+ VPWR VPWR _08186_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_172_4615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_177_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_4626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_424 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28211_ _10838_ _12325_ _12573_ VGND VGND VPWR VPWR _12574_ sky130_fd_sc_hd__a21oi_1
X_25423_ _10967_ VGND VGND VPWR VPWR _02745_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_901 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29191_ _13113_ VGND VGND VPWR VPWR _04367_ sky130_fd_sc_hd__clkbuf_1
X_22635_ _09390_ _09783_ VGND VGND VPWR VPWR _09784_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28142_ _10777_ _12345_ _12482_ VGND VGND VPWR VPWR _12537_ sky130_fd_sc_hd__a21oi_1
X_25354_ _10410_ _10923_ VGND VGND VPWR VPWR _10926_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22566_ _09622_ _09715_ _09718_ VGND VGND VPWR VPWR _09719_ sky130_fd_sc_hd__a21o_1
XFILLER_0_134_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24305_ _10326_ net107 VGND VGND VPWR VPWR _10327_ sky130_fd_sc_hd__nor2_8
X_21517_ _08663_ _08769_ _08771_ _08575_ VGND VGND VPWR VPWR _08772_ sky130_fd_sc_hd__o211a_1
X_28073_ _12500_ VGND VGND VPWR VPWR _03862_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_161_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22497_ _09422_ _09652_ VGND VGND VPWR VPWR _09653_ sky130_fd_sc_hd__nor2_1
X_25285_ _10737_ net2459 _10878_ VGND VGND VPWR VPWR _10885_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27024_ _11889_ net1583 _11897_ _11900_ VGND VGND VPWR VPWR _03413_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_131_3633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_3644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21448_ _08704_ _08705_ _08541_ VGND VGND VPWR VPWR _08706_ sky130_fd_sc_hd__mux2_1
X_24236_ _10289_ VGND VGND VPWR VPWR _02236_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_224_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21379_ rvcpu.dp.rf.reg_file_arr\[24\]\[1\] rvcpu.dp.rf.reg_file_arr\[25\]\[1\] rvcpu.dp.rf.reg_file_arr\[26\]\[1\]
+ rvcpu.dp.rf.reg_file_arr\[27\]\[1\] _08517_ _08519_ VGND VGND VPWR VPWR _08640_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_31_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28975_ _12995_ net1800 _12988_ _12996_ VGND VGND VPWR VPWR _04268_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_34_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold990 datamem.data_ram\[11\]\[28\] VGND VGND VPWR VPWR net2140 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_34_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27926_ _12130_ net4307 _12412_ VGND VGND VPWR VPWR _12415_ sky130_fd_sc_hd__mux2_1
X_15940_ net2185 _13269_ _14297_ VGND VGND VPWR VPWR _14306_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_129_3584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3070 datamem.data_ram\[49\]\[28\] VGND VGND VPWR VPWR net4220 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3081 rvcpu.dp.rf.reg_file_arr\[26\]\[27\] VGND VGND VPWR VPWR net4231 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_30_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3092 datamem.data_ram\[12\]\[11\] VGND VGND VPWR VPWR net4242 sky130_fd_sc_hd__dlygate4sd3_1
X_27857_ _12132_ net4025 _12373_ VGND VGND VPWR VPWR _12377_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15871_ net2047 _13272_ _14258_ VGND VGND VPWR VPWR _14268_ sky130_fd_sc_hd__mux2_1
Xhold2380 datamem.data_ram\[38\]\[29\] VGND VGND VPWR VPWR net3530 sky130_fd_sc_hd__dlygate4sd3_1
X_17610_ _05076_ VGND VGND VPWR VPWR _01232_ sky130_fd_sc_hd__clkbuf_1
X_14822_ _13305_ _13321_ VGND VGND VPWR VPWR _13375_ sky130_fd_sc_hd__nand2_1
X_26808_ _11767_ net1477 _11761_ _11768_ VGND VGND VPWR VPWR _03329_ sky130_fd_sc_hd__a31o_1
Xhold2391 datamem.data_ram\[14\]\[21\] VGND VGND VPWR VPWR net3541 sky130_fd_sc_hd__dlygate4sd3_1
X_18590_ _05832_ VGND VGND VPWR VPWR _05949_ sky130_fd_sc_hd__inv_2
X_27788_ _08125_ _09228_ VGND VGND VPWR VPWR _12335_ sky130_fd_sc_hd__nor2_8
XFILLER_0_25_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17541_ _13266_ net3532 _05032_ VGND VGND VPWR VPWR _05040_ sky130_fd_sc_hd__mux2_1
Xhold1690 datamem.data_ram\[18\]\[10\] VGND VGND VPWR VPWR net2840 sky130_fd_sc_hd__dlygate4sd3_1
X_29527_ clknet_leaf_264_clk _01262_ VGND VGND VPWR VPWR datamem.data_ram\[5\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26739_ _11700_ net1748 _11724_ _11727_ VGND VGND VPWR VPWR _03301_ sky130_fd_sc_hd__a31o_1
X_14753_ rvcpu.dp.pcreg.q\[4\] rvcpu.dp.pcreg.q\[2\] VGND VGND VPWR VPWR _13306_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_103_Left_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_138_3809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29458_ net820 _01193_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[30\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_17472_ _05003_ VGND VGND VPWR VPWR _01305_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1__f__10239_ clknet_0__10239_ VGND VGND VPWR VPWR clknet_1_1__leaf__10239_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_168_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14684_ _13247_ VGND VGND VPWR VPWR _13248_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_86_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19211_ _06519_ VGND VGND VPWR VPWR rvcpu.dp.lAuiPCE\[24\] sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_28_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28409_ _12681_ VGND VGND VPWR VPWR _04017_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16423_ net1990 _14453_ _14572_ VGND VGND VPWR VPWR _14578_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29389_ clknet_leaf_0_clk _01124_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD2E\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31420_ clknet_leaf_53_clk _03123_ VGND VGND VPWR VPWR datamem.data_ram\[15\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_19142_ _06458_ VGND VGND VPWR VPWR _06459_ sky130_fd_sc_hd__inv_2
XFILLER_0_144_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16354_ _14541_ VGND VGND VPWR VPWR _01861_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_60_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_229_6010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_229_6021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15305_ _13312_ _13841_ _13842_ VGND VGND VPWR VPWR _13843_ sky130_fd_sc_hd__and3_1
XFILLER_0_171_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19073_ _06398_ rvcpu.dp.plde.ImmExtE\[7\] _06355_ VGND VGND VPWR VPWR _06399_ sky130_fd_sc_hd__mux2_1
X_31351_ clknet_leaf_18_clk _03054_ VGND VGND VPWR VPWR rvcpu.dp.plde.ImmExtE\[0\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_87_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16285_ net3479 _14451_ _14500_ VGND VGND VPWR VPWR _14505_ sky130_fd_sc_hd__mux2_1
X_23179__850 clknet_1_1__leaf__10111_ VGND VGND VPWR VPWR net976 sky130_fd_sc_hd__inv_2
X_18024_ rvcpu.dp.plde.RD1E\[0\] _05265_ _05269_ _13277_ _05393_ VGND VGND VPWR VPWR
+ _05394_ sky130_fd_sc_hd__a221oi_4
X_30302_ net648 _02037_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[5\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_15236_ _13346_ _13393_ _13592_ _13285_ VGND VGND VPWR VPWR _13776_ sky130_fd_sc_hd__a31o_2
XFILLER_0_164_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31282_ clknet_leaf_110_clk _02985_ VGND VGND VPWR VPWR datamem.data_ram\[34\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__10130_ clknet_0__10130_ VGND VGND VPWR VPWR clknet_1_0__leaf__10130_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_2_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_112_Left_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_75_Right_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30233_ net587 _01968_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[7\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_15167_ _13533_ _13709_ _13710_ _13573_ _13466_ VGND VGND VPWR VPWR _13711_ sky130_fd_sc_hd__o221a_1
XFILLER_0_140_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30164_ net526 _01899_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[0\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_15098_ _13399_ _13642_ VGND VGND VPWR VPWR _13643_ sky130_fd_sc_hd__or2_1
X_19975_ datamem.data_ram\[23\]\[18\] _06706_ _07230_ datamem.data_ram\[20\]\[18\]
+ VGND VGND VPWR VPWR _07269_ sky130_fd_sc_hd__o22a_1
XFILLER_0_201_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18926_ _05531_ _06263_ VGND VGND VPWR VPWR _06265_ sky130_fd_sc_hd__or2_1
XFILLER_0_157_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30095_ net457 _01830_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[11\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_197_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18857_ _05475_ _05484_ _05490_ _05500_ _05665_ _05670_ VGND VGND VPWR VPWR _06201_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_222_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_179_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_230_clk clknet_5_20__leaf_clk VGND VGND VPWR VPWR clknet_leaf_230_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_94_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17808_ rvcpu.dp.plem.ALUResultM\[30\] _05199_ _05178_ VGND VGND VPWR VPWR _05200_
+ sky130_fd_sc_hd__mux2_1
X_18788_ _05658_ _05749_ VGND VGND VPWR VPWR _06136_ sky130_fd_sc_hd__nand2_2
XFILLER_0_82_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_121_Left_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_84_Right_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_210_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32805_ clknet_leaf_164_clk _04227_ VGND VGND VPWR VPWR datamem.data_ram\[13\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17739_ _13257_ net2562 _05140_ VGND VGND VPWR VPWR _05145_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30997_ clknet_leaf_101_clk _02732_ VGND VGND VPWR VPWR datamem.data_ram\[22\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_20750_ datamem.data_ram\[12\]\[6\] datamem.data_ram\[13\]\[6\] _07836_ VGND VGND
+ VPWR VPWR _08040_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32736_ clknet_leaf_167_clk _04158_ VGND VGND VPWR VPWR datamem.data_ram\[16\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_214_5622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_214_5633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19409_ _06704_ VGND VGND VPWR VPWR _06705_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_46_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20681_ datamem.data_ram\[38\]\[5\] _06978_ _06949_ datamem.data_ram\[33\]\[5\] VGND
+ VGND VPWR VPWR _07972_ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32667_ clknet_leaf_251_clk _04089_ VGND VGND VPWR VPWR datamem.data_ram\[19\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_23497__143 clknet_1_1__leaf__10160_ VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__inv_2
XFILLER_0_175_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22420_ rvcpu.dp.rf.reg_file_arr\[28\]\[6\] rvcpu.dp.rf.reg_file_arr\[30\]\[6\] rvcpu.dp.rf.reg_file_arr\[29\]\[6\]
+ rvcpu.dp.rf.reg_file_arr\[31\]\[6\] _09446_ _09402_ VGND VGND VPWR VPWR _09580_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_162_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31618_ clknet_leaf_13_clk net1271 VGND VGND VPWR VPWR rvcpu.dp.plmw.RdW\[4\] sky130_fd_sc_hd__dfxtp_1
X_32598_ clknet_leaf_271_clk _04020_ VGND VGND VPWR VPWR datamem.data_ram\[21\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22351_ rvcpu.dp.rf.reg_file_arr\[16\]\[3\] rvcpu.dp.rf.reg_file_arr\[17\]\[3\] rvcpu.dp.rf.reg_file_arr\[18\]\[3\]
+ rvcpu.dp.rf.reg_file_arr\[19\]\[3\] _09512_ _09513_ VGND VGND VPWR VPWR _09514_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31549_ clknet_leaf_67_clk net1207 VGND VGND VPWR VPWR rvcpu.dp.plmw.ResultSrcW\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_130_Left_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21302_ _08547_ _08556_ _08558_ _08563_ VGND VGND VPWR VPWR _08564_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_93_Right_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25070_ _10765_ VGND VGND VPWR VPWR _02594_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22282_ _09446_ VGND VGND VPWR VPWR _09447_ sky130_fd_sc_hd__buf_4
XFILLER_0_170_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_206_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold220 datamem.data_ram\[47\]\[4\] VGND VGND VPWR VPWR net1370 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21233_ datamem.data_ram\[52\]\[27\] datamem.data_ram\[52\]\[19\] datamem.data_ram\[53\]\[11\]
+ datamem.data_ram\[52\]\[11\] VGND VGND VPWR VPWR _08496_ sky130_fd_sc_hd__or4b_1
XFILLER_0_131_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold231 datamem.data_ram\[38\]\[6\] VGND VGND VPWR VPWR net1381 sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 datamem.data_ram\[5\]\[7\] VGND VGND VPWR VPWR net1392 sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 datamem.data_ram\[3\]\[0\] VGND VGND VPWR VPWR net1403 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__10259_ clknet_0__10259_ VGND VGND VPWR VPWR clknet_1_0__leaf__10259_
+ sky130_fd_sc_hd__clkbuf_16
Xhold264 datamem.data_ram\[33\]\[4\] VGND VGND VPWR VPWR net1414 sky130_fd_sc_hd__dlygate4sd3_1
X_21164_ datamem.data_ram\[1\]\[23\] _07242_ _08452_ _07844_ VGND VGND VPWR VPWR _08453_
+ sky130_fd_sc_hd__o22a_1
Xhold275 datamem.data_ram\[31\]\[3\] VGND VGND VPWR VPWR net1425 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_165_4452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold286 datamem.data_ram\[2\]\[0\] VGND VGND VPWR VPWR net1436 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_165_4463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold297 datamem.data_ram\[59\]\[3\] VGND VGND VPWR VPWR net1447 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20115_ datamem.data_ram\[27\]\[10\] _06731_ _07408_ _06741_ VGND VGND VPWR VPWR
+ _07409_ sky130_fd_sc_hd__o211a_1
X_28760_ _12880_ VGND VGND VPWR VPWR _04169_ sky130_fd_sc_hd__clkbuf_1
X_25972_ _14002_ _11268_ VGND VGND VPWR VPWR _11309_ sky130_fd_sc_hd__nand2_1
X_21095_ datamem.data_ram\[4\]\[7\] datamem.data_ram\[5\]\[7\] _07911_ VGND VGND VPWR
+ VPWR _08384_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_226_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_161_4349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27711_ _12151_ net2867 _12289_ VGND VGND VPWR VPWR _12294_ sky130_fd_sc_hd__mux2_1
X_24923_ _10468_ net3281 net91 VGND VGND VPWR VPWR _10680_ sky130_fd_sc_hd__mux2_1
X_20046_ datamem.data_ram\[8\]\[26\] _06820_ _06632_ datamem.data_ram\[11\]\[26\]
+ VGND VGND VPWR VPWR _07340_ sky130_fd_sc_hd__o22a_1
XFILLER_0_217_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28691_ _12739_ net3617 net42 VGND VGND VPWR VPWR _12844_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_221_clk clknet_5_21__leaf_clk VGND VGND VPWR VPWR clknet_leaf_221_clk
+ sky130_fd_sc_hd__clkbuf_8
X_27642_ _12256_ VGND VGND VPWR VPWR _03675_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_68_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24854_ _10388_ net2800 _10641_ VGND VGND VPWR VPWR _10643_ sky130_fd_sc_hd__mux2_1
X_23349__986 clknet_1_1__leaf__10137_ VGND VGND VPWR VPWR net1112 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_124_3470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_3481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_104 _06924_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27573_ _12089_ net3203 net82 VGND VGND VPWR VPWR _12220_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_115 _07182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24785_ _10470_ net2864 net94 VGND VGND VPWR VPWR _10605_ sky130_fd_sc_hd__mux2_1
XANTENNA_126 _07791_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_200_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21997_ _06603_ _08355_ VGND VGND VPWR VPWR _09227_ sky130_fd_sc_hd__nand2_8
XTAP_TAPCELL_ROW_64_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_217_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29312_ clknet_leaf_290_clk _01047_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD1E\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_137 _07832_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26524_ _10782_ _11604_ _11605_ net1304 VGND VGND VPWR VPWR _03208_ sky130_fd_sc_hd__a22o_1
XFILLER_0_185_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_148 _07872_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_159 _08499_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20948_ _08226_ _08231_ _08237_ _06753_ VGND VGND VPWR VPWR _08238_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_120_3378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__10124_ _10124_ VGND VGND VPWR VPWR clknet_0__10124_ sky130_fd_sc_hd__clkbuf_16
X_29243_ _09223_ net3510 _13141_ VGND VGND VPWR VPWR _13142_ sky130_fd_sc_hd__mux2_1
X_26455_ _11576_ _11218_ _11540_ _06512_ _11581_ VGND VGND VPWR VPWR _11582_ sky130_fd_sc_hd__a221o_1
XFILLER_0_166_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23667_ clknet_1_0__leaf__10192_ VGND VGND VPWR VPWR _10193_ sky130_fd_sc_hd__buf_1
XFILLER_0_37_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20879_ datamem.data_ram\[44\]\[14\] datamem.data_ram\[45\]\[14\] _07827_ VGND VGND
+ VPWR VPWR _08169_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25406_ _10418_ _10950_ VGND VGND VPWR VPWR _10958_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29174_ _13104_ VGND VGND VPWR VPWR _04359_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22618_ _09510_ _09761_ _09763_ _09767_ _09525_ VGND VGND VPWR VPWR _09768_ sky130_fd_sc_hd__a311o_2
X_26386_ _11524_ rvcpu.ALUResultE\[4\] _06377_ _11522_ _11531_ VGND VGND VPWR VPWR
+ _11532_ sky130_fd_sc_hd__a221o_1
XFILLER_0_180_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28125_ _10777_ _12335_ _12482_ VGND VGND VPWR VPWR _12528_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_23_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_288_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_288_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_181_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25337_ _10914_ VGND VGND VPWR VPWR _02712_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_23_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22549_ _09627_ _09700_ _09702_ _09438_ VGND VGND VPWR VPWR _09703_ sky130_fd_sc_hd__a211o_1
XFILLER_0_180_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28056_ _12491_ VGND VGND VPWR VPWR _03854_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16070_ net2033 _13257_ _14371_ VGND VGND VPWR VPWR _14376_ sky130_fd_sc_hd__mux2_1
X_25268_ _10538_ net1437 _10867_ _10875_ VGND VGND VPWR VPWR _02682_ sky130_fd_sc_hd__a31o_1
XFILLER_0_84_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15021_ _13517_ _13567_ _13568_ VGND VGND VPWR VPWR _13569_ sky130_fd_sc_hd__a21oi_1
X_27007_ _11827_ _11886_ VGND VGND VPWR VPWR _11890_ sky130_fd_sc_hd__and2_1
X_24219_ _10280_ VGND VGND VPWR VPWR _02228_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25199_ _10837_ VGND VGND VPWR VPWR _02651_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16972_ net2810 _14455_ _04731_ VGND VGND VPWR VPWR _04738_ sky130_fd_sc_hd__mux2_1
X_19760_ datamem.data_ram\[53\]\[25\] _06723_ _06731_ datamem.data_ram\[51\]\[25\]
+ _06733_ VGND VGND VPWR VPWR _07055_ sky130_fd_sc_hd__o221a_1
X_28958_ _12749_ net2046 _12978_ VGND VGND VPWR VPWR _12986_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_1214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18711_ _05410_ _05726_ _05785_ _05447_ VGND VGND VPWR VPWR _06064_ sky130_fd_sc_hd__o2bb2a_1
X_15923_ _14274_ VGND VGND VPWR VPWR _14297_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_53_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19691_ _06582_ VGND VGND VPWR VPWR _06987_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27909_ _12147_ net4107 net47 VGND VGND VPWR VPWR _12406_ sky130_fd_sc_hd__mux2_1
X_28889_ _12766_ net3295 _12941_ VGND VGND VPWR VPWR _12949_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_212_clk clknet_5_22__leaf_clk VGND VGND VPWR VPWR clknet_leaf_212_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_189_814 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18642_ _05997_ _05599_ VGND VGND VPWR VPWR _05998_ sky130_fd_sc_hd__nand2_1
X_30920_ clknet_leaf_221_clk _02655_ VGND VGND VPWR VPWR datamem.data_ram\[40\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_15854_ _14259_ VGND VGND VPWR VPWR _02095_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_204_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14805_ _13331_ VGND VGND VPWR VPWR _13358_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_157_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18573_ _05931_ _05588_ VGND VGND VPWR VPWR _05932_ sky130_fd_sc_hd__xnor2_1
X_30851_ clknet_leaf_193_clk _02586_ VGND VGND VPWR VPWR datamem.data_ram\[43\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15785_ _14222_ VGND VGND VPWR VPWR _02135_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_204_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17524_ _13241_ net2648 _05021_ VGND VGND VPWR VPWR _05031_ sky130_fd_sc_hd__mux2_1
X_14736_ _13287_ _13288_ VGND VGND VPWR VPWR _13289_ sky130_fd_sc_hd__nand2b_4
XFILLER_0_157_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30782_ clknet_leaf_155_clk _02517_ VGND VGND VPWR VPWR datamem.data_ram\[46\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32521_ clknet_leaf_247_clk _03943_ VGND VGND VPWR VPWR datamem.data_ram\[24\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17455_ _04994_ VGND VGND VPWR VPWR _01313_ sky130_fd_sc_hd__clkbuf_1
X_14667_ _13234_ VGND VGND VPWR VPWR _13235_ sky130_fd_sc_hd__buf_4
XFILLER_0_200_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16406_ net2588 _14436_ _14561_ VGND VGND VPWR VPWR _14569_ sky130_fd_sc_hd__mux2_1
XFILLER_0_223_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32452_ clknet_leaf_254_clk _03874_ VGND VGND VPWR VPWR datamem.data_ram\[27\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17386_ _14168_ net3618 _04949_ VGND VGND VPWR VPWR _04958_ sky130_fd_sc_hd__mux2_1
X_14598_ _13182_ VGND VGND VPWR VPWR _03203_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_229_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19125_ _06421_ _06429_ _06430_ _06435_ _06427_ VGND VGND VPWR VPWR _06444_ sky130_fd_sc_hd__a311o_1
X_31403_ clknet_leaf_43_clk _03106_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCE\[20\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_279_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_279_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_15_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16337_ _14532_ VGND VGND VPWR VPWR _01869_ sky130_fd_sc_hd__clkbuf_1
X_32383_ clknet_leaf_90_clk _03805_ VGND VGND VPWR VPWR datamem.data_ram\[2\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_723 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19056_ _06380_ _06383_ VGND VGND VPWR VPWR _06384_ sky130_fd_sc_hd__xnor2_2
X_31334_ clknet_leaf_16_clk _03037_ VGND VGND VPWR VPWR rvcpu.dp.plde.Rs2E\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_11_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16268_ net2350 _14434_ _14489_ VGND VGND VPWR VPWR _14496_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23650__250 clknet_1_1__leaf__10181_ VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__inv_2
X_18007_ _05375_ _05376_ VGND VGND VPWR VPWR _05377_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15219_ _13372_ _13630_ VGND VGND VPWR VPWR _13760_ sky130_fd_sc_hd__or2_1
X_31265_ clknet_leaf_16_clk _02968_ VGND VGND VPWR VPWR rvcpu.dp.plfd.InstrD\[23\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_112_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16199_ _13225_ VGND VGND VPWR VPWR _14451_ sky130_fd_sc_hd__buf_4
XFILLER_0_26_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24047__575 clknet_1_1__leaf__10246_ VGND VGND VPWR VPWR net701 sky130_fd_sc_hd__inv_2
XFILLER_0_199_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30216_ net570 _01951_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[7\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_31196_ clknet_leaf_46_clk _02899_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCPlus4D\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_207_5470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30147_ net509 _01882_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[0\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_19958_ _06752_ _07246_ _07251_ VGND VGND VPWR VPWR _07252_ sky130_fd_sc_hd__or3_1
X_22975__683 clknet_1_0__leaf__10082_ VGND VGND VPWR VPWR net809 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_203_5356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18909_ _05525_ _05537_ VGND VGND VPWR VPWR _06249_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_203_5367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_5260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30078_ net440 _01813_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[11\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_203_5378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19889_ datamem.data_ram\[28\]\[17\] _07182_ _06659_ datamem.data_ram\[25\]\[17\]
+ _07183_ VGND VGND VPWR VPWR _07184_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_199_5271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_5282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_203_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_203_clk
+ sky130_fd_sc_hd__clkbuf_8
X_21920_ _08813_ _09153_ _08579_ VGND VGND VPWR VPWR _09154_ sky130_fd_sc_hd__a21o_1
XFILLER_0_184_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_1180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_195_5168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_195_5179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21851_ rvcpu.dp.rf.reg_file_arr\[0\]\[24\] rvcpu.dp.rf.reg_file_arr\[1\]\[24\] rvcpu.dp.rf.reg_file_arr\[2\]\[24\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[24\] _08550_ _08554_ VGND VGND VPWR VPWR _09089_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_222_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23505__150 clknet_1_0__leaf__10161_ VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__inv_2
XFILLER_0_210_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20802_ datamem.data_ram\[53\]\[30\] _06663_ _07230_ datamem.data_ram\[52\]\[30\]
+ VGND VGND VPWR VPWR _08092_ sky130_fd_sc_hd__o22a_1
X_24570_ _10485_ VGND VGND VPWR VPWR _02374_ sky130_fd_sc_hd__clkbuf_1
X_21782_ rvcpu.dp.rf.reg_file_arr\[20\]\[21\] rvcpu.dp.rf.reg_file_arr\[21\]\[21\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[21\] rvcpu.dp.rf.reg_file_arr\[23\]\[21\] _08778_
+ _08825_ VGND VGND VPWR VPWR _09023_ sky130_fd_sc_hd__mux4_1
XFILLER_0_148_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23521_ _09256_ net3430 _10162_ VGND VGND VPWR VPWR _10169_ sky130_fd_sc_hd__mux2_1
X_20733_ _08015_ _08017_ _06797_ _08022_ VGND VGND VPWR VPWR _08023_ sky130_fd_sc_hd__o211a_1
X_32719_ clknet_leaf_285_clk _04141_ VGND VGND VPWR VPWR datamem.data_ram\[17\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26240_ _11379_ _03046_ _11454_ VGND VGND VPWR VPWR _03073_ sky130_fd_sc_hd__a21o_1
XFILLER_0_133_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20664_ datamem.data_ram\[57\]\[29\] _06789_ _07953_ _07954_ VGND VGND VPWR VPWR
+ _07955_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_154_4186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_4197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22403_ _09422_ _09563_ _09457_ VGND VGND VPWR VPWR _09564_ sky130_fd_sc_hd__o21ai_1
X_23383_ _07137_ VGND VGND VPWR VPWR _10141_ sky130_fd_sc_hd__buf_12
X_26171_ _11422_ VGND VGND VPWR VPWR _03038_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_208_Left_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20595_ datamem.data_ram\[0\]\[13\] datamem.data_ram\[1\]\[13\] _07827_ VGND VGND
+ VPWR VPWR _07886_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25122_ _10792_ VGND VGND VPWR VPWR _02619_ sky130_fd_sc_hd__clkbuf_1
X_22334_ rvcpu.dp.rf.reg_file_arr\[24\]\[2\] rvcpu.dp.rf.reg_file_arr\[25\]\[2\] rvcpu.dp.rf.reg_file_arr\[26\]\[2\]
+ rvcpu.dp.rf.reg_file_arr\[27\]\[2\] _09385_ _09431_ VGND VGND VPWR VPWR _09498_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_171_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_167_4503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_167_4514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23848__412 clknet_1_1__leaf__10208_ VGND VGND VPWR VPWR net538 sky130_fd_sc_hd__inv_2
XFILLER_0_170_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25053_ _09235_ VGND VGND VPWR VPWR _10754_ sky130_fd_sc_hd__buf_2
X_29930_ net300 _01665_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[16\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22265_ _09430_ VGND VGND VPWR VPWR _09431_ sky130_fd_sc_hd__clkbuf_8
X_21216_ _08487_ _07781_ _08490_ VGND VGND VPWR VPWR _04427_ sky130_fd_sc_hd__o21ai_1
X_29861_ net239 _01596_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[18\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_22196_ _09370_ VGND VGND VPWR VPWR _01115_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_228_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21147_ _08423_ _08428_ _08435_ VGND VGND VPWR VPWR _08436_ sky130_fd_sc_hd__a21o_1
X_28812_ _12908_ VGND VGND VPWR VPWR _04193_ sky130_fd_sc_hd__clkbuf_1
X_29792_ net1138 _01527_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[20\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_3510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_126_3521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28743_ _12871_ VGND VGND VPWR VPWR _04161_ sky130_fd_sc_hd__clkbuf_1
X_25955_ net1795 _11290_ _11286_ _11299_ VGND VGND VPWR VPWR _02945_ sky130_fd_sc_hd__o211a_1
X_21078_ _05371_ _08365_ _08366_ rvcpu.dp.plem.ALUResultM\[4\] VGND VGND VPWR VPWR
+ _08367_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_217_Left_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_226_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20029_ _06911_ _07322_ _06588_ VGND VGND VPWR VPWR _07323_ sky130_fd_sc_hd__or3b_1
X_24906_ _10388_ net3657 _10669_ VGND VGND VPWR VPWR _10671_ sky130_fd_sc_hd__mux2_1
XFILLER_0_214_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28674_ _12756_ net3350 _12832_ VGND VGND VPWR VPWR _12835_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_122_3418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25886_ net1371 _11153_ VGND VGND VPWR VPWR _11260_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_122_3429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27625_ _12247_ VGND VGND VPWR VPWR _03667_ sky130_fd_sc_hd__clkbuf_1
X_24837_ _10633_ VGND VGND VPWR VPWR _02493_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_87_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15570_ _14091_ VGND VGND VPWR VPWR _14092_ sky130_fd_sc_hd__buf_4
X_27556_ _12151_ net2593 net98 VGND VGND VPWR VPWR _12211_ sky130_fd_sc_hd__mux2_1
X_23894__454 clknet_1_0__leaf__10222_ VGND VGND VPWR VPWR net580 sky130_fd_sc_hd__inv_2
X_24768_ _10474_ net4018 _10589_ VGND VGND VPWR VPWR _10594_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_185_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27487_ _12134_ net3316 _12169_ VGND VGND VPWR VPWR _12174_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24699_ _10448_ net4333 _10552_ VGND VGND VPWR VPWR _10557_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_563 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__10107_ _10107_ VGND VGND VPWR VPWR clknet_0__10107_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_138_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17240_ _04880_ VGND VGND VPWR VPWR _01422_ sky130_fd_sc_hd__clkbuf_1
X_29226_ _09297_ net2437 _13132_ VGND VGND VPWR VPWR _13133_ sky130_fd_sc_hd__mux2_1
X_26438_ _11533_ VGND VGND VPWR VPWR _11570_ sky130_fd_sc_hd__buf_2
XFILLER_0_3_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_226_Left_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_193_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29157_ _13095_ VGND VGND VPWR VPWR _04351_ sky130_fd_sc_hd__clkbuf_1
X_17171_ _14158_ net3776 _04840_ VGND VGND VPWR VPWR _04844_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26369_ _11091_ _11511_ VGND VGND VPWR VPWR _11519_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16122_ _14403_ VGND VGND VPWR VPWR _01963_ sky130_fd_sc_hd__clkbuf_1
X_28108_ _10777_ _12325_ _12482_ VGND VGND VPWR VPWR _12519_ sky130_fd_sc_hd__a21oi_2
X_29088_ _09297_ net2330 net40 VGND VGND VPWR VPWR _13059_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28039_ _10500_ VGND VGND VPWR VPWR _12482_ sky130_fd_sc_hd__clkbuf_8
X_16053_ net2411 _13232_ _14360_ VGND VGND VPWR VPWR _14367_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15004_ _13364_ VGND VGND VPWR VPWR _13552_ sky130_fd_sc_hd__inv_2
XFILLER_0_150_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31050_ clknet_leaf_238_clk _02785_ VGND VGND VPWR VPWR datamem.data_ram\[9\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30001_ net371 _01736_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[14\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_19812_ datamem.data_ram\[18\]\[9\] _06613_ VGND VGND VPWR VPWR _07107_ sky130_fd_sc_hd__or2_1
XFILLER_0_208_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19743_ datamem.data_ram\[39\]\[25\] _06726_ _06656_ datamem.data_ram\[33\]\[25\]
+ VGND VGND VPWR VPWR _07038_ sky130_fd_sc_hd__o22a_1
X_16955_ net3437 _14438_ _04720_ VGND VGND VPWR VPWR _04729_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15906_ _14288_ VGND VGND VPWR VPWR _02072_ sky130_fd_sc_hd__clkbuf_1
X_19674_ _06969_ VGND VGND VPWR VPWR _06970_ sky130_fd_sc_hd__clkbuf_4
X_31952_ clknet_leaf_132_clk _03374_ VGND VGND VPWR VPWR datamem.data_ram\[55\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16886_ _04692_ VGND VGND VPWR VPWR _01596_ sky130_fd_sc_hd__clkbuf_1
X_23680__276 clknet_1_0__leaf__10194_ VGND VGND VPWR VPWR net402 sky130_fd_sc_hd__inv_2
XFILLER_0_194_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18625_ _05346_ _05726_ _05974_ _05344_ _05981_ VGND VGND VPWR VPWR _05982_ sky130_fd_sc_hd__a221o_1
X_15837_ _14250_ VGND VGND VPWR VPWR _02103_ sky130_fd_sc_hd__clkbuf_1
X_30903_ clknet_leaf_202_clk _02638_ VGND VGND VPWR VPWR datamem.data_ram\[41\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_31883_ clknet_leaf_124_clk _03337_ VGND VGND VPWR VPWR datamem.data_ram\[57\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26488__42 clknet_1_1__leaf__10267_ VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__inv_2
XFILLER_0_56_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_189_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30834_ clknet_leaf_135_clk _02569_ VGND VGND VPWR VPWR datamem.data_ram\[44\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18556_ _05398_ _05668_ _05663_ _05394_ VGND VGND VPWR VPWR _05916_ sky130_fd_sc_hd__or4_1
X_15768_ _14213_ VGND VGND VPWR VPWR _02143_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_220_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23144__819 clknet_1_0__leaf__10107_ VGND VGND VPWR VPWR net945 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_190_5054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14719_ rvcpu.dp.plmw.ALUResultW\[1\] rvcpu.dp.plmw.ReadDataW\[1\] rvcpu.dp.plmw.PCPlus4W\[1\]
+ rvcpu.dp.plmw.lAuiPCW\[1\] rvcpu.dp.plmw.ResultSrcW\[0\] rvcpu.dp.plmw.ResultSrcW\[1\]
+ VGND VGND VPWR VPWR _13274_ sky130_fd_sc_hd__mux4_2
XFILLER_0_75_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17507_ _05022_ VGND VGND VPWR VPWR _01289_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_190_5065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18487_ _05342_ _05769_ _05848_ _05689_ VGND VGND VPWR VPWR _05849_ sky130_fd_sc_hd__o211a_1
X_30765_ clknet_leaf_265_clk _02500_ VGND VGND VPWR VPWR datamem.data_ram\[47\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_15699_ _13240_ VGND VGND VPWR VPWR _14170_ sky130_fd_sc_hd__buf_4
XANTENNA_490 _09750_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_883 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17438_ _14151_ net3467 _04985_ VGND VGND VPWR VPWR _04986_ sky130_fd_sc_hd__mux2_1
X_32504_ clknet_leaf_275_clk _03926_ VGND VGND VPWR VPWR datamem.data_ram\[25\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_31747__124 VGND VGND VPWR VPWR _31747__124/HI net124 sky130_fd_sc_hd__conb_1
X_30696_ clknet_leaf_154_clk _02431_ VGND VGND VPWR VPWR datamem.data_ram\[4\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_15 _06612_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_26 _06632_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_37 _06671_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_48 _06680_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32435_ clknet_leaf_240_clk _03857_ VGND VGND VPWR VPWR datamem.data_ram\[27\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17369_ _04937_ VGND VGND VPWR VPWR _04949_ sky130_fd_sc_hd__buf_4
XANTENNA_59 _06714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19108_ _06427_ _06428_ VGND VGND VPWR VPWR _06429_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32366_ clknet_leaf_93_clk _03788_ VGND VGND VPWR VPWR datamem.data_ram\[2\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_20380_ datamem.data_ram\[63\]\[28\] _06669_ _07671_ _06599_ VGND VGND VPWR VPWR
+ _07672_ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_209_5510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_209_5521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19039_ _06367_ _06368_ VGND VGND VPWR VPWR _06369_ sky130_fd_sc_hd__nand2_1
XFILLER_0_179_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31317_ clknet_leaf_28_clk _03020_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCPlus4E\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32297_ clknet_leaf_161_clk _03719_ VGND VGND VPWR VPWR datamem.data_ram\[32\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22050_ _09271_ VGND VGND VPWR VPWR _01068_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_205_5407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31248_ clknet_leaf_21_clk _02951_ VGND VGND VPWR VPWR rvcpu.dp.plfd.InstrD\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_205_5418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21001_ datamem.data_ram\[21\]\[15\] _06660_ _06643_ datamem.data_ram\[16\]\[15\]
+ VGND VGND VPWR VPWR _08290_ sky130_fd_sc_hd__o22a_1
XFILLER_0_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2902 datamem.data_ram\[57\]\[28\] VGND VGND VPWR VPWR net4052 sky130_fd_sc_hd__dlygate4sd3_1
X_31179_ clknet_leaf_188_clk _02882_ VGND VGND VPWR VPWR datamem.data_ram\[5\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_5_7__f_clk clknet_2_0_0_clk VGND VGND VPWR VPWR clknet_5_7__leaf_clk sky130_fd_sc_hd__clkbuf_16
Xhold2913 rvcpu.dp.rf.reg_file_arr\[27\]\[27\] VGND VGND VPWR VPWR net4063 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2924 datamem.data_ram\[17\]\[16\] VGND VGND VPWR VPWR net4074 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2935 datamem.data_ram\[33\]\[26\] VGND VGND VPWR VPWR net4085 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_197_5219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2946 datamem.data_ram\[59\]\[19\] VGND VGND VPWR VPWR net4096 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2957 datamem.data_ram\[2\]\[10\] VGND VGND VPWR VPWR net4107 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2968 rvcpu.dp.rf.reg_file_arr\[26\]\[24\] VGND VGND VPWR VPWR net4118 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_214_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25740_ _11145_ VGND VGND VPWR VPWR _11146_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_177_1275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2979 datamem.data_ram\[0\]\[17\] VGND VGND VPWR VPWR net4129 sky130_fd_sc_hd__dlygate4sd3_1
X_22952_ clknet_5_4__leaf_clk VGND VGND VPWR VPWR _10078_ sky130_fd_sc_hd__buf_1
XFILLER_0_98_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21903_ _08692_ _09135_ _09137_ VGND VGND VPWR VPWR _09138_ sky130_fd_sc_hd__a21o_1
XFILLER_0_218_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25671_ _06587_ VGND VGND VPWR VPWR _11104_ sky130_fd_sc_hd__buf_2
XFILLER_0_223_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22883_ rvcpu.dp.rf.reg_file_arr\[12\]\[30\] rvcpu.dp.rf.reg_file_arr\[13\]\[30\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[30\] rvcpu.dp.rf.reg_file_arr\[15\]\[30\] _09462_
+ _09465_ VGND VGND VPWR VPWR _10019_ sky130_fd_sc_hd__mux4_1
Xmax_cap39 _13085_ VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__buf_4
X_27410_ _09223_ VGND VGND VPWR VPWR _12125_ sky130_fd_sc_hd__buf_2
X_24622_ _10444_ net2993 _10511_ VGND VGND VPWR VPWR _10514_ sky130_fd_sc_hd__mux2_1
X_28390_ _12671_ VGND VGND VPWR VPWR _04008_ sky130_fd_sc_hd__clkbuf_1
X_21834_ _08547_ _09070_ _09072_ _08576_ VGND VGND VPWR VPWR _09073_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_156_4237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_156_4248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27341_ _12085_ net2762 _12081_ VGND VGND VPWR VPWR _12086_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_195_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24553_ _10474_ net3672 net60 VGND VGND VPWR VPWR _10475_ sky130_fd_sc_hd__mux2_1
X_21765_ _08522_ _09006_ VGND VGND VPWR VPWR _09007_ sky130_fd_sc_hd__or2_1
XFILLER_0_109_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20716_ datamem.data_ram\[23\]\[5\] _06927_ _08005_ _08006_ VGND VGND VPWR VPWR _08007_
+ sky130_fd_sc_hd__a211o_1
X_23657__256 clknet_1_1__leaf__10191_ VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__inv_2
X_27272_ _12047_ VGND VGND VPWR VPWR _03514_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24484_ _10432_ VGND VGND VPWR VPWR _02341_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21696_ _08627_ _08937_ _08939_ _08941_ VGND VGND VPWR VPWR _08942_ sky130_fd_sc_hd__o2bb2a_1
X_29011_ _12995_ net1715 _13009_ _13016_ VGND VGND VPWR VPWR _04284_ sky130_fd_sc_hd__a31o_1
XFILLER_0_34_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26223_ _11449_ VGND VGND VPWR VPWR _03063_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20647_ datamem.data_ram\[26\]\[29\] _06803_ _06789_ datamem.data_ram\[25\]\[29\]
+ _06851_ VGND VGND VPWR VPWR _07938_ sky130_fd_sc_hd__o221a_1
XFILLER_0_19_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_191_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26154_ rvcpu.dp.plfd.InstrD\[13\] _11413_ VGND VGND VPWR VPWR _11414_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_115_3255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20578_ _07863_ _07864_ _07865_ _07868_ VGND VGND VPWR VPWR _07869_ sky130_fd_sc_hd__o22a_1
XFILLER_0_190_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25105_ _10783_ _10779_ _10781_ net1361 VGND VGND VPWR VPWR _02611_ sky130_fd_sc_hd__a22o_1
X_22317_ _09481_ VGND VGND VPWR VPWR _09482_ sky130_fd_sc_hd__buf_4
XFILLER_0_108_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26085_ rvcpu.dp.plfd.InstrD\[2\] rvcpu.dp.plfd.InstrD\[0\] VGND VGND VPWR VPWR _11376_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_186_4956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_186_4967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_225_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29913_ net283 _01648_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[16\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_25036_ _10744_ VGND VGND VPWR VPWR _02581_ sky130_fd_sc_hd__clkbuf_1
X_24143__647 clknet_1_0__leaf__10262_ VGND VGND VPWR VPWR net773 sky130_fd_sc_hd__inv_2
XFILLER_0_104_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22248_ _09397_ _09405_ _09410_ _09412_ _09413_ VGND VGND VPWR VPWR _09414_ sky130_fd_sc_hd__a221o_1
X_22179_ _09230_ VGND VGND VPWR VPWR _09361_ sky130_fd_sc_hd__buf_8
X_29844_ net222 _01579_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[18\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_50_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26987_ _10756_ net2542 _11875_ VGND VGND VPWR VPWR _11878_ sky130_fd_sc_hd__mux2_1
X_29775_ net1121 _01510_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[20\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_219_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_145_3974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16740_ _04615_ VGND VGND VPWR VPWR _01673_ sky130_fd_sc_hd__clkbuf_1
X_25938_ net1843 _11279_ VGND VGND VPWR VPWR _11291_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_145_3985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28726_ _12862_ VGND VGND VPWR VPWR _04153_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_199_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23902__461 clknet_1_0__leaf__10223_ VGND VGND VPWR VPWR net587 sky130_fd_sc_hd__inv_2
X_16671_ _14135_ net2866 _04576_ VGND VGND VPWR VPWR _04579_ sky130_fd_sc_hd__mux2_1
X_28657_ _12692_ net3548 _12823_ VGND VGND VPWR VPWR _12826_ sky130_fd_sc_hd__mux2_1
XFILLER_0_202_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25869_ rvcpu.dp.pcreg.q\[30\] rvcpu.dp.pcreg.q\[29\] _11239_ VGND VGND VPWR VPWR
+ _11247_ sky130_fd_sc_hd__and3_1
XFILLER_0_198_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18410_ _05768_ _05770_ _05773_ _05707_ VGND VGND VPWR VPWR _05774_ sky130_fd_sc_hd__o211a_1
X_15622_ _14119_ VGND VGND VPWR VPWR _02195_ sky130_fd_sc_hd__clkbuf_1
X_19390_ _06685_ VGND VGND VPWR VPWR _06686_ sky130_fd_sc_hd__buf_8
X_27608_ _12238_ VGND VGND VPWR VPWR _03659_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_185_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28588_ _12739_ net4325 _12786_ VGND VGND VPWR VPWR _12789_ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18341_ _05705_ VGND VGND VPWR VPWR _05706_ sky130_fd_sc_hd__buf_2
XFILLER_0_9_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15553_ _13378_ _13767_ _13780_ _13398_ VGND VGND VPWR VPWR _14077_ sky130_fd_sc_hd__o22a_1
X_27539_ _12134_ net3469 _12197_ VGND VGND VPWR VPWR _12202_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_104_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_104_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18272_ rvcpu.dp.plde.RD1E\[26\] _05564_ _05544_ VGND VGND VPWR VPWR _05637_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_127_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30550_ clknet_leaf_178_clk _02285_ VGND VGND VPWR VPWR datamem.data_ram\[55\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_13_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15484_ _14010_ _13501_ _13409_ _14012_ VGND VGND VPWR VPWR _14013_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_16_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17223_ _04871_ VGND VGND VPWR VPWR _01430_ sky130_fd_sc_hd__clkbuf_1
X_29209_ _10047_ _13123_ VGND VGND VPWR VPWR _13124_ sky130_fd_sc_hd__and2_1
XFILLER_0_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_583 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30481_ net159 _02216_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[19\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32220_ clknet_leaf_227_clk _03642_ VGND VGND VPWR VPWR datamem.data_ram\[35\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17154_ _14141_ net2886 _04829_ VGND VGND VPWR VPWR _04835_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16105_ _14394_ VGND VGND VPWR VPWR _01971_ sky130_fd_sc_hd__clkbuf_1
Xhold808 datamem.data_ram\[38\]\[22\] VGND VGND VPWR VPWR net1958 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32151_ clknet_leaf_209_clk _03573_ VGND VGND VPWR VPWR datamem.data_ram\[38\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold819 datamem.data_ram\[44\]\[15\] VGND VGND VPWR VPWR net1969 sky130_fd_sc_hd__dlygate4sd3_1
X_17085_ _04798_ VGND VGND VPWR VPWR _01495_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_172_Right_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31102_ clknet_leaf_106_clk _02837_ VGND VGND VPWR VPWR datamem.data_ram\[19\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16036_ net1913 _13207_ _14349_ VGND VGND VPWR VPWR _14358_ sky130_fd_sc_hd__mux2_1
X_32082_ clknet_leaf_62_clk _03504_ VGND VGND VPWR VPWR datamem.data_ram\[47\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31033_ clknet_leaf_55_clk _02768_ VGND VGND VPWR VPWR datamem.data_ram\[12\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_196_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2209 rvcpu.dp.rf.reg_file_arr\[25\]\[8\] VGND VGND VPWR VPWR net3359 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1508 datamem.data_ram\[54\]\[14\] VGND VGND VPWR VPWR net2658 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_200_5304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17987_ rvcpu.dp.plem.ALUResultM\[5\] _05272_ VGND VGND VPWR VPWR _05357_ sky130_fd_sc_hd__and2_1
X_23762__351 clknet_1_0__leaf__10201_ VGND VGND VPWR VPWR net477 sky130_fd_sc_hd__inv_2
Xhold1519 datamem.data_ram\[14\]\[25\] VGND VGND VPWR VPWR net2669 sky130_fd_sc_hd__dlygate4sd3_1
X_19726_ _07020_ VGND VGND VPWR VPWR _07021_ sky130_fd_sc_hd__buf_6
XFILLER_0_165_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16938_ _04719_ VGND VGND VPWR VPWR _04720_ sky130_fd_sc_hd__buf_4
X_32984_ clknet_leaf_173_clk _04406_ VGND VGND VPWR VPWR datamem.data_ram\[63\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31935_ clknet_leaf_123_clk _03357_ VGND VGND VPWR VPWR datamem.data_ram\[59\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_192_5105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19657_ _06666_ _06917_ VGND VGND VPWR VPWR _06953_ sky130_fd_sc_hd__nor2_8
X_16869_ _14089_ _14347_ VGND VGND VPWR VPWR _04683_ sky130_fd_sc_hd__nor2_2
XFILLER_0_149_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18608_ _05914_ _05965_ _05768_ VGND VGND VPWR VPWR _05966_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31866_ clknet_leaf_110_clk _03320_ VGND VGND VPWR VPWR datamem.data_ram\[63\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_19588_ datamem.data_ram\[47\]\[8\] _06670_ _06883_ _06851_ VGND VGND VPWR VPWR _06884_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_149_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18539_ _05625_ _05632_ _05633_ _05637_ _05667_ _05663_ VGND VGND VPWR VPWR _05900_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_133_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30817_ clknet_leaf_261_clk _02552_ VGND VGND VPWR VPWR datamem.data_ram\[45\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31797_ clknet_leaf_209_clk _03251_ VGND VGND VPWR VPWR datamem.data_ram\[2\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21550_ rvcpu.dp.rf.reg_file_arr\[28\]\[9\] rvcpu.dp.rf.reg_file_arr\[30\]\[9\] rvcpu.dp.rf.reg_file_arr\[29\]\[9\]
+ rvcpu.dp.rf.reg_file_arr\[31\]\[9\] _08559_ _08636_ VGND VGND VPWR VPWR _08803_
+ sky130_fd_sc_hd__mux4_1
X_30748_ clknet_leaf_130_clk _02483_ VGND VGND VPWR VPWR datamem.data_ram\[48\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_151_4112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_4123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20501_ datamem.data_ram\[47\]\[21\] _07791_ _07182_ datamem.data_ram\[44\]\[21\]
+ VGND VGND VPWR VPWR _07792_ sky130_fd_sc_hd__o22a_1
XFILLER_0_69_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21481_ _08572_ _08737_ VGND VGND VPWR VPWR _08738_ sky130_fd_sc_hd__or2_1
X_30679_ clknet_leaf_96_clk _02414_ VGND VGND VPWR VPWR datamem.data_ram\[4\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_209_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20432_ datamem.data_ram\[10\]\[12\] _06612_ _07720_ _07723_ VGND VGND VPWR VPWR
+ _07724_ sky130_fd_sc_hd__o211a_1
X_32418_ clknet_leaf_81_clk _03840_ VGND VGND VPWR VPWR datamem.data_ram\[28\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_715 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload240 clknet_leaf_120_clk VGND VGND VPWR VPWR clkload240/Y sky130_fd_sc_hd__clkinv_4
X_23151_ clknet_1_1__leaf__10108_ VGND VGND VPWR VPWR _10109_ sky130_fd_sc_hd__buf_1
X_20363_ datamem.data_ram\[5\]\[28\] _06702_ _07653_ _07654_ VGND VGND VPWR VPWR _07655_
+ sky130_fd_sc_hd__o211a_1
Xclkload251 clknet_leaf_154_clk VGND VGND VPWR VPWR clkload251/Y sky130_fd_sc_hd__bufinv_16
X_32349_ clknet_leaf_170_clk _03771_ VGND VGND VPWR VPWR datamem.data_ram\[30\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_23447__97 clknet_1_1__leaf__10156_ VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_228_5963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload262 clknet_leaf_195_clk VGND VGND VPWR VPWR clkload262/Y sky130_fd_sc_hd__bufinv_16
Xclkload273 clknet_leaf_127_clk VGND VGND VPWR VPWR clkload273/Y sky130_fd_sc_hd__clkinv_1
X_22102_ rvcpu.dp.plem.WriteDataM\[27\] _09221_ _09295_ rvcpu.dp.plem.WriteDataM\[11\]
+ _09312_ VGND VGND VPWR VPWR _09313_ sky130_fd_sc_hd__a221o_4
XFILLER_0_114_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_110_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_228_5974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload284 clknet_1_1__leaf__10246_ VGND VGND VPWR VPWR clkload284/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_110_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_4063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20294_ datamem.data_ram\[15\]\[19\] _06726_ _06766_ datamem.data_ram\[12\]\[19\]
+ _07586_ VGND VGND VPWR VPWR _07587_ sky130_fd_sc_hd__o221a_1
Xclkload295 clknet_1_1__leaf__10221_ VGND VGND VPWR VPWR clkload295/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_149_4074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_282 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26910_ _11752_ VGND VGND VPWR VPWR _11831_ sky130_fd_sc_hd__clkbuf_4
X_22033_ _09256_ net3531 _09232_ VGND VGND VPWR VPWR _09257_ sky130_fd_sc_hd__mux2_1
X_27890_ _11968_ _12394_ VGND VGND VPWR VPWR _12396_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_181_4831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_181_4842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2710 datamem.data_ram\[51\]\[25\] VGND VGND VPWR VPWR net3860 sky130_fd_sc_hd__dlygate4sd3_1
X_26841_ _11781_ net1738 _11785_ _11788_ VGND VGND VPWR VPWR _03342_ sky130_fd_sc_hd__a31o_1
Xhold2721 datamem.data_ram\[23\]\[21\] VGND VGND VPWR VPWR net3871 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_71_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23090__770 clknet_1_0__leaf__10102_ VGND VGND VPWR VPWR net896 sky130_fd_sc_hd__inv_2
Xhold2732 rvcpu.dp.rf.reg_file_arr\[16\]\[22\] VGND VGND VPWR VPWR net3882 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2743 datamem.data_ram\[31\]\[14\] VGND VGND VPWR VPWR net3893 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2754 rvcpu.dp.rf.reg_file_arr\[20\]\[4\] VGND VGND VPWR VPWR net3904 sky130_fd_sc_hd__dlygate4sd3_1
X_29560_ net914 _01295_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[27\]\[27\] sky130_fd_sc_hd__dfxtp_1
Xhold2765 datamem.data_ram\[8\]\[28\] VGND VGND VPWR VPWR net3915 sky130_fd_sc_hd__dlygate4sd3_1
X_26772_ _11672_ _11738_ VGND VGND VPWR VPWR _11746_ sky130_fd_sc_hd__and2_1
X_23012__716 clknet_1_0__leaf__10086_ VGND VGND VPWR VPWR net842 sky130_fd_sc_hd__inv_2
Xhold2776 datamem.data_ram\[4\]\[13\] VGND VGND VPWR VPWR net3926 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2787 datamem.data_ram\[28\]\[8\] VGND VGND VPWR VPWR net3937 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_216_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28511_ _12742_ VGND VGND VPWR VPWR _04058_ sky130_fd_sc_hd__clkbuf_1
Xhold2798 datamem.data_ram\[12\]\[9\] VGND VGND VPWR VPWR net3948 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_108_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25723_ _11135_ VGND VGND VPWR VPWR _02877_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_108_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22935_ _10056_ net1472 _10046_ _10065_ VGND VGND VPWR VPWR _01159_ sky130_fd_sc_hd__a31o_1
X_29491_ net853 _01226_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[2\]\[30\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_84_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_179_4782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28442_ _09329_ VGND VGND VPWR VPWR _12702_ sky130_fd_sc_hd__clkbuf_2
X_25654_ _10782_ _11094_ _11095_ net1452 VGND VGND VPWR VPWR _02848_ sky130_fd_sc_hd__a22o_1
XFILLER_0_190_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_179_4793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22866_ _09452_ _10000_ _10002_ _09795_ VGND VGND VPWR VPWR _10003_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_80_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24605_ _10470_ net3513 _10502_ VGND VGND VPWR VPWR _10505_ sky130_fd_sc_hd__mux2_1
X_21817_ _09056_ VGND VGND VPWR VPWR _01050_ sky130_fd_sc_hd__clkbuf_1
X_28373_ _12361_ net3753 _12659_ VGND VGND VPWR VPWR _12662_ sky130_fd_sc_hd__mux2_1
X_25585_ _09299_ _11054_ _10052_ VGND VGND VPWR VPWR _11055_ sky130_fd_sc_hd__and3_2
XFILLER_0_195_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22797_ rvcpu.dp.rf.reg_file_arr\[20\]\[26\] rvcpu.dp.rf.reg_file_arr\[21\]\[26\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[26\] rvcpu.dp.rf.reg_file_arr\[23\]\[26\] _09434_
+ _09558_ VGND VGND VPWR VPWR _09937_ sky130_fd_sc_hd__mux4_1
XFILLER_0_39_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27324_ _10058_ _12076_ _12077_ net1537 VGND VGND VPWR VPWR _03536_ sky130_fd_sc_hd__a22o_1
XFILLER_0_182_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24536_ _10463_ VGND VGND VPWR VPWR _02362_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_3306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21748_ rvcpu.dp.rf.reg_file_arr\[24\]\[19\] rvcpu.dp.rf.reg_file_arr\[25\]\[19\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[19\] rvcpu.dp.rf.reg_file_arr\[27\]\[19\] _08548_
+ _08526_ VGND VGND VPWR VPWR _08991_ sky130_fd_sc_hd__mux4_1
XFILLER_0_136_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27255_ _09231_ net52 VGND VGND VPWR VPWR _12042_ sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_159_Left_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24467_ _10423_ VGND VGND VPWR VPWR _02333_ sky130_fd_sc_hd__clkbuf_1
X_21679_ rvcpu.dp.rf.reg_file_arr\[0\]\[15\] rvcpu.dp.rf.reg_file_arr\[1\]\[15\] rvcpu.dp.rf.reg_file_arr\[2\]\[15\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[15\] _08810_ _08811_ VGND VGND VPWR VPWR _08926_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_0_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23932__487 clknet_1_0__leaf__10227_ VGND VGND VPWR VPWR net613 sky130_fd_sc_hd__inv_2
XFILLER_0_151_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26206_ net1864 _02993_ _03037_ _11441_ VGND VGND VPWR VPWR _03054_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27186_ _11946_ _11996_ VGND VGND VPWR VPWR _12001_ sky130_fd_sc_hd__and2_1
XFILLER_0_62_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24398_ _10378_ VGND VGND VPWR VPWR _02309_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_78_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26137_ _11404_ VGND VGND VPWR VPWR _03021_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23631__248 clknet_1_0__leaf__10181_ VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__inv_2
XFILLER_0_120_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26068_ rvcpu.dp.plfd.InstrD\[12\] _08622_ VGND VGND VPWR VPWR _11364_ sky130_fd_sc_hd__and2_1
XFILLER_0_104_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_219_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17910_ _05281_ _05282_ VGND VGND VPWR VPWR _05283_ sky130_fd_sc_hd__and2_1
X_25019_ _09281_ VGND VGND VPWR VPWR _10733_ sky130_fd_sc_hd__buf_2
X_18890_ _05694_ _06113_ _06231_ _06109_ VGND VGND VPWR VPWR _06232_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_119_28 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_37_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_168_Left_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17841_ rvcpu.dp.plem.ALUResultM\[17\] _05221_ _05177_ VGND VGND VPWR VPWR _05222_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_7_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29827_ net205 _01562_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[1\]\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_7_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14984_ _13425_ _13531_ _13470_ VGND VGND VPWR VPWR _13532_ sky130_fd_sc_hd__a21oi_1
X_17772_ rvcpu.dp.plem.RdM\[1\] _05165_ _05168_ _05169_ rvcpu.dp.plem.RegWriteM VGND
+ VGND VPWR VPWR _05170_ sky130_fd_sc_hd__o221a_1
X_29758_ net1104 _01493_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[21\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19511_ _06695_ VGND VGND VPWR VPWR _06807_ sky130_fd_sc_hd__buf_6
XFILLER_0_135_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16723_ _14187_ net2469 _04598_ VGND VGND VPWR VPWR _04606_ sky130_fd_sc_hd__mux2_1
X_28709_ _12853_ VGND VGND VPWR VPWR _04145_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29689_ net1035 _01424_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[23\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23525__153 clknet_1_1__leaf__10161_ VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__inv_2
XFILLER_0_159_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19442_ _06737_ VGND VGND VPWR VPWR _06738_ sky130_fd_sc_hd__buf_6
X_16654_ _04569_ VGND VGND VPWR VPWR _01713_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_18_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31720_ net169 _03178_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[9\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_198_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15605_ _14110_ VGND VGND VPWR VPWR _02203_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_201_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31651_ clknet_leaf_26_clk net1189 VGND VGND VPWR VPWR rvcpu.dp.plmw.lAuiPCW\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_16585_ _04532_ VGND VGND VPWR VPWR _01753_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19373_ _06668_ VGND VGND VPWR VPWR _06669_ sky130_fd_sc_hd__buf_4
XFILLER_0_97_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15536_ _13512_ _13965_ _13823_ VGND VGND VPWR VPWR _14062_ sky130_fd_sc_hd__o21ai_1
X_18324_ _05688_ VGND VGND VPWR VPWR _05689_ sky130_fd_sc_hd__clkbuf_4
X_30602_ clknet_leaf_217_clk _02337_ VGND VGND VPWR VPWR datamem.data_ram\[53\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_31582_ clknet_leaf_67_clk net1222 VGND VGND VPWR VPWR rvcpu.dp.plmw.PCPlus4W\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_210_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23792__377 clknet_1_1__leaf__10205_ VGND VGND VPWR VPWR net503 sky130_fd_sc_hd__inv_2
XFILLER_0_155_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18255_ _05461_ _05467_ _05473_ VGND VGND VPWR VPWR _05620_ sky130_fd_sc_hd__nor3_1
XFILLER_0_60_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30533_ clknet_leaf_206_clk _02268_ VGND VGND VPWR VPWR datamem.data_ram\[55\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_15467_ _13381_ _13996_ _13706_ VGND VGND VPWR VPWR _13997_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_154_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_503 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24011__544 clknet_1_1__leaf__10241_ VGND VGND VPWR VPWR net670 sky130_fd_sc_hd__inv_2
XFILLER_0_155_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17206_ _14193_ net3533 _04828_ VGND VGND VPWR VPWR _04862_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18186_ _05530_ VGND VGND VPWR VPWR _05551_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30464_ net142 _02199_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[19\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_15398_ _13928_ _13930_ _13897_ _13864_ VGND VGND VPWR VPWR _13931_ sky130_fd_sc_hd__and4b_1
XFILLER_0_181_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32203_ clknet_leaf_167_clk _03625_ VGND VGND VPWR VPWR datamem.data_ram\[36\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_17137_ _04825_ VGND VGND VPWR VPWR _01470_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold605 datamem.data_ram\[2\]\[1\] VGND VGND VPWR VPWR net1755 sky130_fd_sc_hd__dlygate4sd3_1
X_30395_ net733 _02130_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[31\]\[6\] sky130_fd_sc_hd__dfxtp_1
Xhold616 datamem.data_ram\[10\]\[3\] VGND VGND VPWR VPWR net1766 sky130_fd_sc_hd__dlygate4sd3_1
Xhold627 rvcpu.dp.plfd.PCPlus4D\[27\] VGND VGND VPWR VPWR net1777 sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 datamem.data_ram\[36\]\[3\] VGND VGND VPWR VPWR net1788 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32134_ clknet_leaf_236_clk _03556_ VGND VGND VPWR VPWR datamem.data_ram\[10\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold649 datamem.data_ram\[24\]\[6\] VGND VGND VPWR VPWR net1799 sky130_fd_sc_hd__dlygate4sd3_1
X_17068_ net2288 _14482_ _04779_ VGND VGND VPWR VPWR _04789_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16019_ _14348_ VGND VGND VPWR VPWR _14349_ sky130_fd_sc_hd__buf_4
X_32065_ clknet_leaf_121_clk _03487_ VGND VGND VPWR VPWR datamem.data_ram\[29\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_228_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2006 datamem.data_ram\[26\]\[17\] VGND VGND VPWR VPWR net3156 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31016_ clknet_leaf_155_clk _02751_ VGND VGND VPWR VPWR datamem.data_ram\[42\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23686__282 clknet_1_1__leaf__10194_ VGND VGND VPWR VPWR net408 sky130_fd_sc_hd__inv_2
XFILLER_0_209_353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2017 datamem.data_ram\[16\]\[17\] VGND VGND VPWR VPWR net3167 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2028 datamem.data_ram\[59\]\[8\] VGND VGND VPWR VPWR net3178 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2039 rvcpu.dp.rf.reg_file_arr\[28\]\[7\] VGND VGND VPWR VPWR net3189 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1305 rvcpu.dp.rf.reg_file_arr\[0\]\[27\] VGND VGND VPWR VPWR net2455 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1316 datamem.data_ram\[34\]\[19\] VGND VGND VPWR VPWR net2466 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1327 datamem.data_ram\[63\]\[15\] VGND VGND VPWR VPWR net2477 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1338 datamem.data_ram\[2\]\[11\] VGND VGND VPWR VPWR net2488 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1349 rvcpu.dp.rf.reg_file_arr\[17\]\[3\] VGND VGND VPWR VPWR net2499 sky130_fd_sc_hd__dlygate4sd3_1
X_19709_ datamem.data_ram\[21\]\[0\] _06920_ _06954_ datamem.data_ram\[20\]\[0\] VGND
+ VGND VPWR VPWR _07005_ sky130_fd_sc_hd__a22o_1
XFILLER_0_174_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_224_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20981_ datamem.data_ram\[12\]\[15\] datamem.data_ram\[13\]\[15\] _06650_ VGND VGND
+ VPWR VPWR _08270_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32967_ clknet_leaf_200_clk _04389_ VGND VGND VPWR VPWR datamem.data_ram\[63\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22720_ _09482_ _09864_ VGND VGND VPWR VPWR _09865_ sky130_fd_sc_hd__or2_1
X_31918_ _04430_ net119 VGND VGND VPWR VPWR datamem.rd_data_mem\[23\] sky130_fd_sc_hd__dlxtn_1
XFILLER_0_149_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32898_ clknet_leaf_211_clk _04320_ VGND VGND VPWR VPWR datamem.data_ram\[0\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22651_ rvcpu.dp.rf.reg_file_arr\[20\]\[18\] rvcpu.dp.rf.reg_file_arr\[21\]\[18\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[18\] rvcpu.dp.rf.reg_file_arr\[23\]\[18\] _09401_
+ _09430_ VGND VGND VPWR VPWR _09799_ sky130_fd_sc_hd__mux4_1
X_31849_ clknet_leaf_124_clk _03303_ VGND VGND VPWR VPWR datamem.data_ram\[61\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_217_5697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21602_ _08531_ _08850_ _08852_ _08806_ VGND VGND VPWR VPWR _08853_ sky130_fd_sc_hd__o211a_1
X_25370_ _09299_ _10935_ _10052_ VGND VGND VPWR VPWR _10936_ sky130_fd_sc_hd__and3_2
XFILLER_0_36_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22582_ _09441_ _09733_ VGND VGND VPWR VPWR _09734_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24321_ _09330_ net3486 _10328_ VGND VGND VPWR VPWR _10336_ sky130_fd_sc_hd__mux2_1
XFILLER_0_173_650 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21533_ rvcpu.dp.rf.reg_file_arr\[4\]\[8\] rvcpu.dp.rf.reg_file_arr\[5\]\[8\] rvcpu.dp.rf.reg_file_arr\[6\]\[8\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[8\] _08551_ _08555_ VGND VGND VPWR VPWR _08787_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_170_4565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_170_4576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27040_ _10402_ _11039_ VGND VGND VPWR VPWR _11909_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_170_4587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24252_ _10297_ _09301_ _10269_ VGND VGND VPWR VPWR _10298_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_181_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21464_ _08559_ VGND VGND VPWR VPWR _08721_ sky130_fd_sc_hd__buf_4
XFILLER_0_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23122__799 clknet_1_1__leaf__10105_ VGND VGND VPWR VPWR net925 sky130_fd_sc_hd__inv_2
X_23203_ _10122_ VGND VGND VPWR VPWR _01370_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20415_ datamem.data_ram\[59\]\[12\] _06737_ _07703_ _07706_ VGND VGND VPWR VPWR
+ _07707_ sky130_fd_sc_hd__o211a_1
X_21395_ rvcpu.dp.rf.reg_file_arr\[20\]\[2\] rvcpu.dp.rf.reg_file_arr\[21\]\[2\] rvcpu.dp.rf.reg_file_arr\[22\]\[2\]
+ rvcpu.dp.rf.reg_file_arr\[23\]\[2\] _08631_ _08632_ VGND VGND VPWR VPWR _08655_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_222_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23769__357 clknet_1_0__leaf__10202_ VGND VGND VPWR VPWR net483 sky130_fd_sc_hd__inv_2
X_20346_ datamem.data_ram\[63\]\[4\] _07125_ _07634_ _07637_ VGND VGND VPWR VPWR _07638_
+ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_73_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28991_ _12698_ net2410 _12999_ VGND VGND VPWR VPWR _13005_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_73_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20277_ datamem.data_ram\[45\]\[19\] _06768_ _06696_ datamem.data_ram\[40\]\[19\]
+ _07569_ VGND VGND VPWR VPWR _07570_ sky130_fd_sc_hd__o221a_1
X_27942_ _12423_ VGND VGND VPWR VPWR _03808_ sky130_fd_sc_hd__clkbuf_1
X_23065_ _10094_ VGND VGND VPWR VPWR _01260_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold3230 datamem.data_ram\[2\]\[23\] VGND VGND VPWR VPWR net4380 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3241 datamem.data_ram\[55\]\[30\] VGND VGND VPWR VPWR net4391 sky130_fd_sc_hd__dlygate4sd3_1
X_22016_ rvcpu.dp.plem.WriteDataM\[3\] _09215_ _09219_ _09242_ VGND VGND VPWR VPWR
+ _09243_ sky130_fd_sc_hd__a31o_4
X_27873_ _12385_ VGND VGND VPWR VPWR _03777_ sky130_fd_sc_hd__clkbuf_1
Xhold3252 rvcpu.dp.rf.reg_file_arr\[24\]\[14\] VGND VGND VPWR VPWR net4402 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3263 rvcpu.dp.rf.reg_file_arr\[24\]\[5\] VGND VGND VPWR VPWR net4413 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3274 rvcpu.dp.plde.ImmExtE\[14\] VGND VGND VPWR VPWR net4424 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_175_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold3285 datamem.data_ram\[2\]\[16\] VGND VGND VPWR VPWR net4435 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2540 rvcpu.dp.rf.reg_file_arr\[30\]\[4\] VGND VGND VPWR VPWR net3690 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3296 rvcpu.dp.plfd.InstrD\[8\] VGND VGND VPWR VPWR net4446 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2551 datamem.data_ram\[1\]\[11\] VGND VGND VPWR VPWR net3701 sky130_fd_sc_hd__dlygate4sd3_1
X_29612_ net966 _01347_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[25\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_26824_ _11684_ _11774_ VGND VGND VPWR VPWR _11778_ sky130_fd_sc_hd__and2_1
XFILLER_0_192_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2562 datamem.data_ram\[34\]\[11\] VGND VGND VPWR VPWR net3712 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2573 datamem.data_ram\[15\]\[25\] VGND VGND VPWR VPWR net3723 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_879 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2584 rvcpu.dp.rf.reg_file_arr\[23\]\[16\] VGND VGND VPWR VPWR net3734 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2595 datamem.data_ram\[20\]\[24\] VGND VGND VPWR VPWR net3745 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1850 datamem.data_ram\[8\]\[14\] VGND VGND VPWR VPWR net3000 sky130_fd_sc_hd__dlygate4sd3_1
X_26755_ _11725_ _10947_ VGND VGND VPWR VPWR _11736_ sky130_fd_sc_hd__or2_1
X_29543_ net897 _01278_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[27\]\[10\] sky130_fd_sc_hd__dfxtp_1
Xhold1861 datamem.data_ram\[60\]\[25\] VGND VGND VPWR VPWR net3011 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1872 datamem.data_ram\[25\]\[16\] VGND VGND VPWR VPWR net3022 sky130_fd_sc_hd__dlygate4sd3_1
X_23967_ _10237_ VGND VGND VPWR VPWR _02019_ sky130_fd_sc_hd__clkbuf_1
Xhold1883 rvcpu.dp.rf.reg_file_arr\[16\]\[9\] VGND VGND VPWR VPWR net3033 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1894 datamem.data_ram\[51\]\[27\] VGND VGND VPWR VPWR net3044 sky130_fd_sc_hd__dlygate4sd3_1
X_25706_ _11126_ VGND VGND VPWR VPWR _02869_ sky130_fd_sc_hd__clkbuf_1
X_22918_ _10051_ VGND VGND VPWR VPWR _10052_ sky130_fd_sc_hd__buf_2
X_26686_ _11681_ _11694_ VGND VGND VPWR VPWR _11697_ sky130_fd_sc_hd__and2_1
X_29474_ net836 _01209_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[2\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25637_ _11085_ net1407 _11077_ _11087_ VGND VGND VPWR VPWR _02839_ sky130_fd_sc_hd__a31o_1
XFILLER_0_195_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28425_ _12690_ net4122 _12688_ VGND VGND VPWR VPWR _12691_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22849_ _09978_ _09982_ _09986_ _09389_ VGND VGND VPWR VPWR _01152_ sky130_fd_sc_hd__o31a_1
XFILLER_0_13_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28356_ _12452_ net4116 net95 VGND VGND VPWR VPWR _12653_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16370_ net1931 _14468_ _14547_ VGND VGND VPWR VPWR _14550_ sky130_fd_sc_hd__mux2_1
X_25568_ _11018_ net1433 _11041_ _11044_ VGND VGND VPWR VPWR _02813_ sky130_fd_sc_hd__a31o_1
XFILLER_0_94_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27307_ _12061_ net1759 _12065_ _12068_ VGND VGND VPWR VPWR _03528_ sky130_fd_sc_hd__a31o_1
X_15321_ _13307_ _13350_ VGND VGND VPWR VPWR _13858_ sky130_fd_sc_hd__or2_2
XFILLER_0_186_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_3748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24519_ _09259_ VGND VGND VPWR VPWR _10454_ sky130_fd_sc_hd__buf_2
XFILLER_0_93_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_3759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28287_ _12435_ net2237 _12613_ VGND VGND VPWR VPWR _12616_ sky130_fd_sc_hd__mux2_1
XFILLER_0_192_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25499_ _11004_ VGND VGND VPWR VPWR _02784_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_62_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18040_ net103 _05409_ VGND VGND VPWR VPWR _05410_ sky130_fd_sc_hd__xnor2_4
XTAP_TAPCELL_ROW_62_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15252_ _13539_ _13791_ VGND VGND VPWR VPWR _13792_ sky130_fd_sc_hd__nand2_1
X_27238_ _12022_ net1565 _12030_ _12032_ VGND VGND VPWR VPWR _03495_ sky130_fd_sc_hd__a31o_1
XFILLER_0_164_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24149__653 clknet_1_1__leaf__10262_ VGND VGND VPWR VPWR net779 sky130_fd_sc_hd__inv_2
X_23555__179 clknet_1_0__leaf__10174_ VGND VGND VPWR VPWR net305 sky130_fd_sc_hd__inv_2
XFILLER_0_62_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15183_ _13431_ _13289_ _13403_ _13307_ _13646_ VGND VGND VPWR VPWR _13726_ sky130_fd_sc_hd__o2111a_1
X_27169_ _11974_ net1729 _11983_ _11990_ VGND VGND VPWR VPWR _03468_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23097__776 clknet_1_0__leaf__10103_ VGND VGND VPWR VPWR net902 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_39_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30180_ clknet_leaf_203_clk _01915_ VGND VGND VPWR VPWR datamem.data_ram\[58\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_19991_ datamem.data_ram\[6\]\[2\] _06950_ _06924_ datamem.data_ram\[7\]\[2\] _07284_
+ VGND VGND VPWR VPWR _07285_ sky130_fd_sc_hd__a221o_1
X_23426__78 clknet_1_1__leaf__10154_ VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__inv_2
XFILLER_0_104_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_176_Left_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_197_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18942_ _05531_ _05537_ _06251_ _05635_ VGND VGND VPWR VPWR _06280_ sky130_fd_sc_hd__o31a_1
XFILLER_0_197_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18873_ _05694_ _05941_ VGND VGND VPWR VPWR _06216_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17824_ _05210_ VGND VGND VPWR VPWR rvcpu.dp.SrcBFW_Mux.y\[25\] sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_20_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2 rvcpu.dp.plem.lAuiPCM\[19\] VGND VGND VPWR VPWR net1152 sky130_fd_sc_hd__dlygate4sd3_1
X_32821_ clknet_leaf_236_clk _04243_ VGND VGND VPWR VPWR datamem.data_ram\[12\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_14967_ _13504_ _13508_ _13515_ _13456_ VGND VGND VPWR VPWR _13516_ sky130_fd_sc_hd__a211oi_1
X_17755_ _13176_ rvcpu.dp.plde.Rs2E\[4\] VGND VGND VPWR VPWR _05153_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_221_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16706_ _14170_ net3262 _04587_ VGND VGND VPWR VPWR _04597_ sky130_fd_sc_hd__mux2_1
X_32752_ clknet_leaf_189_clk _04174_ VGND VGND VPWR VPWR datamem.data_ram\[15\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_14898_ _13397_ _13387_ VGND VGND VPWR VPWR _13449_ sky130_fd_sc_hd__and2_2
X_17686_ _05116_ VGND VGND VPWR VPWR _01196_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_187_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_185_Left_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31703_ clknet_leaf_42_clk _03161_ VGND VGND VPWR VPWR rvcpu.dp.pcreg.q\[21\] sky130_fd_sc_hd__dfxtp_1
X_19425_ _06660_ VGND VGND VPWR VPWR _06721_ sky130_fd_sc_hd__buf_6
X_16637_ _04560_ VGND VGND VPWR VPWR _01721_ sky130_fd_sc_hd__clkbuf_1
X_32683_ clknet_leaf_171_clk _04105_ VGND VGND VPWR VPWR datamem.data_ram\[18\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31634_ clknet_leaf_47_clk net1209 VGND VGND VPWR VPWR rvcpu.dp.plmw.lAuiPCW\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_19356_ _06651_ VGND VGND VPWR VPWR _06652_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_70_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16568_ _04523_ VGND VGND VPWR VPWR _01761_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_174_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18307_ _05313_ _05334_ _05320_ _05327_ _05666_ _05671_ VGND VGND VPWR VPWR _05672_
+ sky130_fd_sc_hd__mux4_1
X_15519_ _13737_ _13656_ VGND VGND VPWR VPWR _14046_ sky130_fd_sc_hd__nand2_1
X_31565_ clknet_leaf_71_clk datamem.rd_data_mem\[15\] VGND VGND VPWR VPWR rvcpu.dp.plmw.ReadDataW\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_19287_ _06580_ _06582_ VGND VGND VPWR VPWR _06583_ sky130_fd_sc_hd__nand2_2
XFILLER_0_143_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16499_ net4182 _14459_ _04478_ VGND VGND VPWR VPWR _04487_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_212_5572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23041__742 clknet_1_0__leaf__10089_ VGND VGND VPWR VPWR net868 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_212_5583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18238_ rvcpu.dp.plde.RD1E\[15\] _05266_ _05271_ _13231_ _05312_ VGND VGND VPWR VPWR
+ _05603_ sky130_fd_sc_hd__a221oi_4
X_30516_ clknet_leaf_203_clk _02251_ VGND VGND VPWR VPWR datamem.data_ram\[56\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_212_5594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31496_ clknet_leaf_29_clk rvcpu.dp.lAuiPCE\[22\] VGND VGND VPWR VPWR rvcpu.dp.plem.lAuiPCM\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30447_ net785 _02182_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[29\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_18169_ rvcpu.dp.plde.ImmExtE\[24\] rvcpu.dp.SrcBFW_Mux.y\[24\] _05279_ VGND VGND
+ VPWR VPWR _05534_ sky130_fd_sc_hd__mux2_1
Xhold402 datamem.data_ram\[45\]\[7\] VGND VGND VPWR VPWR net1552 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap110 net111 VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__clkbuf_2
Xhold413 datamem.data_ram\[21\]\[2\] VGND VGND VPWR VPWR net1563 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_225_5900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_194_Left_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20200_ datamem.data_ram\[62\]\[11\] _06763_ _06702_ datamem.data_ram\[61\]\[11\]
+ VGND VGND VPWR VPWR _07493_ sky130_fd_sc_hd__o22a_1
Xhold424 datamem.data_ram\[31\]\[6\] VGND VGND VPWR VPWR net1574 sky130_fd_sc_hd__dlygate4sd3_1
X_21180_ _08468_ _08408_ VGND VGND VPWR VPWR _08469_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold435 datamem.data_ram\[45\]\[6\] VGND VGND VPWR VPWR net1585 sky130_fd_sc_hd__dlygate4sd3_1
X_30378_ net724 _02113_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[3\]\[29\] sky130_fd_sc_hd__dfxtp_1
Xhold446 datamem.data_ram\[37\]\[6\] VGND VGND VPWR VPWR net1596 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_4000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold457 datamem.data_ram\[6\]\[4\] VGND VGND VPWR VPWR net1607 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_4011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold468 datamem.data_ram\[63\]\[3\] VGND VGND VPWR VPWR net1618 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20131_ datamem.data_ram\[14\]\[27\] _06682_ _06671_ datamem.data_ram\[15\]\[27\]
+ _07423_ VGND VGND VPWR VPWR _07424_ sky130_fd_sc_hd__o221a_1
X_32117_ clknet_leaf_98_clk _03539_ VGND VGND VPWR VPWR datamem.data_ram\[0\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold479 datamem.data_ram\[31\]\[1\] VGND VGND VPWR VPWR net1629 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_221_5808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32048_ clknet_leaf_132_clk _03470_ VGND VGND VPWR VPWR datamem.data_ram\[49\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_20062_ datamem.data_ram\[60\]\[26\] _06684_ _07242_ datamem.data_ram\[57\]\[26\]
+ _07355_ VGND VGND VPWR VPWR _07356_ sky130_fd_sc_hd__o221a_1
XFILLER_0_29_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_176_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1102 rvcpu.dp.rf.reg_file_arr\[4\]\[0\] VGND VGND VPWR VPWR net2252 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1113 datamem.data_ram\[50\]\[22\] VGND VGND VPWR VPWR net2263 sky130_fd_sc_hd__dlygate4sd3_1
X_24870_ _10651_ VGND VGND VPWR VPWR _02508_ sky130_fd_sc_hd__clkbuf_1
Xhold1124 rvcpu.dp.rf.reg_file_arr\[19\]\[11\] VGND VGND VPWR VPWR net2274 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1135 datamem.data_ram\[56\]\[25\] VGND VGND VPWR VPWR net2285 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1146 rvcpu.dp.rf.reg_file_arr\[1\]\[17\] VGND VGND VPWR VPWR net2296 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1157 datamem.data_ram\[3\]\[15\] VGND VGND VPWR VPWR net2307 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1168 rvcpu.dp.rf.reg_file_arr\[11\]\[1\] VGND VGND VPWR VPWR net2318 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1179 rvcpu.dp.rf.reg_file_arr\[4\]\[22\] VGND VGND VPWR VPWR net2329 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26540_ _11086_ _11610_ VGND VGND VPWR VPWR _11614_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_219_5748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_308 _14160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_219_5759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_176_4730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20964_ datamem.data_ram\[56\]\[15\] _06644_ _08249_ _08252_ VGND VGND VPWR VPWR
+ _08253_ sky130_fd_sc_hd__o211a_1
XANTENNA_319 _14187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0__10140_ _10140_ VGND VGND VPWR VPWR clknet_0__10140_ sky130_fd_sc_hd__clkbuf_16
X_22703_ _09705_ _09840_ _09844_ _09848_ VGND VGND VPWR VPWR _09849_ sky130_fd_sc_hd__and4_1
X_26471_ net1860 _11573_ _11592_ _10041_ VGND VGND VPWR VPWR _03168_ sky130_fd_sc_hd__o211a_1
XFILLER_0_152_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_4616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20895_ datamem.data_ram\[0\]\[22\] _06649_ _08184_ _07851_ _06681_ VGND VGND VPWR
+ VPWR _08185_ sky130_fd_sc_hd__o221a_1
XFILLER_0_137_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28210_ _06591_ VGND VGND VPWR VPWR _12573_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_172_4627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25422_ _10762_ net3861 _10961_ VGND VGND VPWR VPWR _10967_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29190_ _09297_ net2590 _13112_ VGND VGND VPWR VPWR _13113_ sky130_fd_sc_hd__mux2_1
X_22634_ rvcpu.dp.rf.reg_file_arr\[24\]\[17\] rvcpu.dp.rf.reg_file_arr\[25\]\[17\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[17\] rvcpu.dp.rf.reg_file_arr\[27\]\[17\] _09392_
+ _09394_ VGND VGND VPWR VPWR _09783_ sky130_fd_sc_hd__mux4_1
XFILLER_0_165_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28141_ _12536_ VGND VGND VPWR VPWR _03894_ sky130_fd_sc_hd__clkbuf_1
X_25353_ _10876_ net1473 _10920_ _10925_ VGND VGND VPWR VPWR _02717_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_957 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22565_ _09528_ _09717_ _09426_ VGND VGND VPWR VPWR _09718_ sky130_fd_sc_hd__a21o_1
XFILLER_0_180_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24304_ _06681_ _08355_ VGND VGND VPWR VPWR _10326_ sky130_fd_sc_hd__nand2_8
XFILLER_0_111_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23474__122 clknet_1_1__leaf__10158_ VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__inv_2
XFILLER_0_134_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28072_ _12371_ net3139 _12492_ VGND VGND VPWR VPWR _12500_ sky130_fd_sc_hd__mux2_1
X_21516_ _08542_ _08770_ VGND VGND VPWR VPWR _08771_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25284_ _10884_ VGND VGND VPWR VPWR _02689_ sky130_fd_sc_hd__clkbuf_1
X_22496_ rvcpu.dp.rf.reg_file_arr\[16\]\[10\] rvcpu.dp.rf.reg_file_arr\[17\]\[10\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[10\] rvcpu.dp.rf.reg_file_arr\[19\]\[10\] _09385_
+ _09637_ VGND VGND VPWR VPWR _09652_ sky130_fd_sc_hd__mux4_2
XFILLER_0_32_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27023_ _11822_ _11899_ VGND VGND VPWR VPWR _11900_ sky130_fd_sc_hd__and2_1
XFILLER_0_146_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_3634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24235_ _09267_ net3621 _10288_ VGND VGND VPWR VPWR _10289_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_131_3645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21447_ rvcpu.dp.rf.reg_file_arr\[20\]\[4\] rvcpu.dp.rf.reg_file_arr\[21\]\[4\] rvcpu.dp.rf.reg_file_arr\[22\]\[4\]
+ rvcpu.dp.rf.reg_file_arr\[23\]\[4\] _08631_ _08632_ VGND VGND VPWR VPWR _08705_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_20_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21378_ _08532_ _08638_ VGND VGND VPWR VPWR _08639_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_9_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23117_ clknet_1_1__leaf__10087_ VGND VGND VPWR VPWR _10105_ sky130_fd_sc_hd__buf_1
X_20329_ _07071_ _07615_ _07620_ _06713_ VGND VGND VPWR VPWR _07621_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_92_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28974_ _10069_ _12989_ VGND VGND VPWR VPWR _12996_ sky130_fd_sc_hd__and2_1
X_23018__722 clknet_1_1__leaf__10086_ VGND VGND VPWR VPWR net848 sky130_fd_sc_hd__inv_2
Xhold980 datamem.data_ram\[38\]\[23\] VGND VGND VPWR VPWR net2130 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold991 rvcpu.dp.rf.reg_file_arr\[8\]\[8\] VGND VGND VPWR VPWR net2141 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_34_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27925_ _12414_ VGND VGND VPWR VPWR _03800_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_34_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3060 datamem.data_ram\[11\]\[14\] VGND VGND VPWR VPWR net4210 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3071 datamem.data_ram\[60\]\[23\] VGND VGND VPWR VPWR net4221 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_3596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3082 rvcpu.dp.rf.reg_file_arr\[10\]\[17\] VGND VGND VPWR VPWR net4232 sky130_fd_sc_hd__dlygate4sd3_1
X_15870_ _14267_ VGND VGND VPWR VPWR _02087_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_215_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27856_ _12376_ VGND VGND VPWR VPWR _03769_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_30_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3093 datamem.data_ram\[24\]\[10\] VGND VGND VPWR VPWR net4243 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2370 rvcpu.dp.rf.reg_file_arr\[4\]\[26\] VGND VGND VPWR VPWR net3520 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14821_ _13373_ VGND VGND VPWR VPWR _13374_ sky130_fd_sc_hd__clkbuf_4
Xhold2381 datamem.data_ram\[62\]\[22\] VGND VGND VPWR VPWR net3531 sky130_fd_sc_hd__dlygate4sd3_1
X_26807_ _11645_ _11762_ VGND VGND VPWR VPWR _11768_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2392 rvcpu.dp.rf.reg_file_arr\[19\]\[23\] VGND VGND VPWR VPWR net3542 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_1104 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24999_ _10720_ VGND VGND VPWR VPWR _02568_ sky130_fd_sc_hd__clkbuf_1
X_27787_ _12334_ VGND VGND VPWR VPWR _03742_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_192_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_203_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1680 datamem.data_ram\[5\]\[31\] VGND VGND VPWR VPWR net2830 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14752_ _13288_ VGND VGND VPWR VPWR _13305_ sky130_fd_sc_hd__buf_4
X_17540_ _05039_ VGND VGND VPWR VPWR _01273_ sky130_fd_sc_hd__clkbuf_1
Xhold1691 rvcpu.dp.rf.reg_file_arr\[14\]\[13\] VGND VGND VPWR VPWR net2841 sky130_fd_sc_hd__dlygate4sd3_1
X_29526_ clknet_leaf_271_clk _01261_ VGND VGND VPWR VPWR datamem.data_ram\[5\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_26738_ _11676_ _11726_ VGND VGND VPWR VPWR _11727_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17471_ _14185_ net3659 _04996_ VGND VGND VPWR VPWR _05003_ sky130_fd_sc_hd__mux2_1
X_26669_ _11645_ _11677_ VGND VGND VPWR VPWR _11686_ sky130_fd_sc_hd__and2_1
X_14683_ rvcpu.dp.plmw.ALUResultW\[10\] rvcpu.dp.plmw.ReadDataW\[10\] rvcpu.dp.plmw.PCPlus4W\[10\]
+ rvcpu.dp.plmw.lAuiPCW\[10\] _13169_ _13171_ VGND VGND VPWR VPWR _13247_ sky130_fd_sc_hd__mux4_2
X_23326__965 clknet_1_1__leaf__10135_ VGND VGND VPWR VPWR net1091 sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__10238_ clknet_0__10238_ VGND VGND VPWR VPWR clknet_1_1__leaf__10238_
+ sky130_fd_sc_hd__clkbuf_16
X_29457_ net819 _01192_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[30\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19210_ _06518_ rvcpu.dp.plde.ImmExtE\[24\] _06493_ VGND VGND VPWR VPWR _06519_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28408_ _12452_ net3192 _12678_ VGND VGND VPWR VPWR _12681_ sky130_fd_sc_hd__mux2_1
X_16422_ _14577_ VGND VGND VPWR VPWR _01829_ sky130_fd_sc_hd__clkbuf_1
X_23938__493 clknet_1_0__leaf__10227_ VGND VGND VPWR VPWR net619 sky130_fd_sc_hd__inv_2
X_29388_ clknet_leaf_174_clk _01123_ VGND VGND VPWR VPWR datamem.data_ram\[60\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19141_ _06441_ _06450_ VGND VGND VPWR VPWR _06458_ sky130_fd_sc_hd__nand2_1
XFILLER_0_144_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16353_ net4232 _14451_ _14536_ VGND VGND VPWR VPWR _14541_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28339_ _12435_ net3636 _12641_ VGND VGND VPWR VPWR _12644_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_229_6000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_229_6011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15304_ _13487_ _13350_ _13513_ VGND VGND VPWR VPWR _13842_ sky130_fd_sc_hd__a21o_1
XFILLER_0_26_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19072_ _06396_ _06397_ VGND VGND VPWR VPWR _06398_ sky130_fd_sc_hd__xor2_2
X_31350_ clknet_leaf_68_clk _03053_ VGND VGND VPWR VPWR rvcpu.dp.plde.ResultSrcE\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_229_6022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16284_ _14504_ VGND VGND VPWR VPWR _01894_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30301_ net647 _02036_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[5\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_15235_ _13762_ _13765_ _13770_ _13775_ _13572_ VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__o32a_1
XFILLER_0_180_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18023_ _05391_ _05293_ VGND VGND VPWR VPWR _05393_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31281_ clknet_leaf_126_clk _02984_ VGND VGND VPWR VPWR datamem.data_ram\[24\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30232_ net586 _01967_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[7\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_15166_ _13308_ _13565_ _13577_ VGND VGND VPWR VPWR _13710_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_58_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30163_ net525 _01898_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[0\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_15097_ _13454_ _13477_ VGND VGND VPWR VPWR _13642_ sky130_fd_sc_hd__or2_1
X_19974_ datamem.data_ram\[31\]\[18\] _06707_ _07264_ _07267_ VGND VGND VPWR VPWR
+ _07268_ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18925_ _05531_ _06263_ VGND VGND VPWR VPWR _06264_ sky130_fd_sc_hd__nand2_1
X_30094_ net456 _01829_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[11\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18856_ _05693_ _05925_ _05927_ _06136_ VGND VGND VPWR VPWR _06200_ sky130_fd_sc_hd__a211o_1
XFILLER_0_59_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_206_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17807_ _13183_ rvcpu.dp.plde.RD2E\[30\] _05196_ VGND VGND VPWR VPWR _05199_ sky130_fd_sc_hd__mux2_1
XFILLER_0_222_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18787_ _05513_ _05616_ VGND VGND VPWR VPWR _06135_ sky130_fd_sc_hd__nand2_1
X_15999_ _14337_ VGND VGND VPWR VPWR _02028_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_206_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32804_ clknet_leaf_163_clk _04226_ VGND VGND VPWR VPWR datamem.data_ram\[13\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_222_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17738_ _05144_ VGND VGND VPWR VPWR _01172_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_221_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30996_ clknet_leaf_99_clk _02731_ VGND VGND VPWR VPWR datamem.data_ram\[13\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23798__383 clknet_1_1__leaf__10205_ VGND VGND VPWR VPWR net509 sky130_fd_sc_hd__inv_2
XFILLER_0_221_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32735_ clknet_leaf_86_clk _04157_ VGND VGND VPWR VPWR datamem.data_ram\[16\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_1307 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_187_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17669_ net2703 _13253_ _05104_ VGND VGND VPWR VPWR _05108_ sky130_fd_sc_hd__mux2_1
XFILLER_0_202_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_214_5623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_392 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19408_ _06667_ VGND VGND VPWR VPWR _06704_ sky130_fd_sc_hd__buf_8
XFILLER_0_58_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_214_5634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20680_ datamem.data_ram\[37\]\[5\] _07132_ _07123_ datamem.data_ram\[36\]\[5\] VGND
+ VGND VPWR VPWR _07971_ sky130_fd_sc_hd__a22o_1
XFILLER_0_169_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32666_ clknet_leaf_285_clk _04088_ VGND VGND VPWR VPWR datamem.data_ram\[19\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31617_ clknet_leaf_14_clk net1262 VGND VGND VPWR VPWR rvcpu.dp.plmw.RdW\[3\] sky130_fd_sc_hd__dfxtp_4
X_19339_ _06634_ VGND VGND VPWR VPWR _06635_ sky130_fd_sc_hd__buf_6
XFILLER_0_70_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32597_ clknet_leaf_288_clk _04019_ VGND VGND VPWR VPWR datamem.data_ram\[21\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22350_ _09394_ VGND VGND VPWR VPWR _09513_ sky130_fd_sc_hd__buf_4
XFILLER_0_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31548_ clknet_leaf_67_clk net1159 VGND VGND VPWR VPWR rvcpu.dp.plmw.ResultSrcW\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_116_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21301_ _08542_ _08562_ VGND VGND VPWR VPWR _08563_ sky130_fd_sc_hd__or2_1
X_22281_ _08595_ VGND VGND VPWR VPWR _09446_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_206_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31479_ clknet_leaf_48_clk rvcpu.dp.lAuiPCE\[5\] VGND VGND VPWR VPWR rvcpu.dp.plem.lAuiPCM\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold210 datamem.data_ram\[47\]\[2\] VGND VGND VPWR VPWR net1360 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21232_ _08492_ _08493_ _08494_ VGND VGND VPWR VPWR _08495_ sky130_fd_sc_hd__or3_1
XFILLER_0_206_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold221 rvcpu.dp.plfd.PCD\[2\] VGND VGND VPWR VPWR net1371 sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 datamem.data_ram\[13\]\[6\] VGND VGND VPWR VPWR net1382 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__10258_ clknet_0__10258_ VGND VGND VPWR VPWR clknet_1_0__leaf__10258_
+ sky130_fd_sc_hd__clkbuf_16
Xhold243 datamem.data_ram\[39\]\[0\] VGND VGND VPWR VPWR net1393 sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 datamem.data_ram\[3\]\[3\] VGND VGND VPWR VPWR net1404 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold265 datamem.data_ram\[43\]\[1\] VGND VGND VPWR VPWR net1415 sky130_fd_sc_hd__dlygate4sd3_1
X_21163_ _08450_ _08451_ _07819_ VGND VGND VPWR VPWR _08452_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold276 datamem.data_ram\[56\]\[1\] VGND VGND VPWR VPWR net1426 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_165_4453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold287 datamem.data_ram\[3\]\[6\] VGND VGND VPWR VPWR net1437 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_165_4464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold298 datamem.data_ram\[2\]\[6\] VGND VGND VPWR VPWR net1448 sky130_fd_sc_hd__dlygate4sd3_1
X_20114_ datamem.data_ram\[30\]\[10\] _06626_ _06669_ datamem.data_ram\[31\]\[10\]
+ _07407_ VGND VGND VPWR VPWR _07408_ sky130_fd_sc_hd__o221a_1
X_21094_ datamem.data_ram\[6\]\[7\] datamem.data_ram\[7\]\[7\] _07824_ VGND VGND VPWR
+ VPWR _08383_ sky130_fd_sc_hd__mux2_1
X_25971_ net4451 _11302_ _11300_ _11308_ VGND VGND VPWR VPWR _02952_ sky130_fd_sc_hd__o211a_1
X_24922_ _10679_ VGND VGND VPWR VPWR _02532_ sky130_fd_sc_hd__clkbuf_1
X_27710_ _12293_ VGND VGND VPWR VPWR _03706_ sky130_fd_sc_hd__clkbuf_1
X_20045_ datamem.data_ram\[14\]\[26\] _06744_ _07243_ datamem.data_ram\[9\]\[26\]
+ VGND VGND VPWR VPWR _07339_ sky130_fd_sc_hd__o22a_1
X_28690_ _12843_ VGND VGND VPWR VPWR _04136_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_217_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_198_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_225_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27641_ _12134_ net2548 _12251_ VGND VGND VPWR VPWR _12256_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24853_ _10642_ VGND VGND VPWR VPWR _02500_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_68_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_3460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_3471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_3482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27572_ _12219_ VGND VGND VPWR VPWR _03642_ sky130_fd_sc_hd__clkbuf_1
X_24784_ _10604_ VGND VGND VPWR VPWR _02469_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_105 _06934_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_213_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_212_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_116 _07182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21996_ _09225_ VGND VGND VPWR VPWR _09226_ sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_64_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_127 _07808_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26523_ _10064_ _11604_ _11605_ net1321 VGND VGND VPWR VPWR _03207_ sky130_fd_sc_hd__a22o_1
X_29311_ clknet_leaf_290_clk _01046_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD1E\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_64_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_138 _07832_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20947_ _07823_ _08233_ _08236_ _07081_ VGND VGND VPWR VPWR _08237_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_120_3368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23048__748 clknet_1_0__leaf__10090_ VGND VGND VPWR VPWR net874 sky130_fd_sc_hd__inv_2
XANTENNA_149 _07874_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26454_ _11535_ rvcpu.ALUResultE\[23\] _11288_ VGND VGND VPWR VPWR _11581_ sky130_fd_sc_hd__a21o_1
XFILLER_0_166_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29242_ _12601_ _09229_ _09230_ VGND VGND VPWR VPWR _13141_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_49_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23666_ clknet_1_0__leaf__10078_ VGND VGND VPWR VPWR _10192_ sky130_fd_sc_hd__buf_1
XFILLER_0_95_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20878_ datamem.data_ram\[40\]\[14\] _06648_ _08167_ _07851_ VGND VGND VPWR VPWR
+ _08168_ sky130_fd_sc_hd__o22a_1
X_25405_ _10954_ net1716 _10949_ _10957_ VGND VGND VPWR VPWR _02737_ sky130_fd_sc_hd__a31o_1
XFILLER_0_187_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29173_ _09223_ net4053 net63 VGND VGND VPWR VPWR _13104_ sky130_fd_sc_hd__mux2_1
X_22617_ _09451_ _09764_ _09766_ _09523_ VGND VGND VPWR VPWR _09767_ sky130_fd_sc_hd__o211a_1
X_26385_ _08620_ _08621_ _11154_ _11157_ VGND VGND VPWR VPWR _11531_ sky130_fd_sc_hd__a31o_1
XFILLER_0_165_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24070__596 clknet_1_1__leaf__10248_ VGND VGND VPWR VPWR net722 sky130_fd_sc_hd__inv_2
XFILLER_0_76_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28124_ _12527_ VGND VGND VPWR VPWR _03886_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_187_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25336_ _10760_ net4292 _10909_ VGND VGND VPWR VPWR _10914_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_98_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22548_ _09534_ _09701_ VGND VGND VPWR VPWR _09702_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_23_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_180_269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28055_ _12462_ net4097 _12483_ VGND VGND VPWR VPWR _12491_ sky130_fd_sc_hd__mux2_1
X_25267_ _10418_ _10868_ VGND VGND VPWR VPWR _10875_ sky130_fd_sc_hd__and2_1
XFILLER_0_224_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22479_ _09391_ VGND VGND VPWR VPWR _09636_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_94_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23710__304 clknet_1_1__leaf__10196_ VGND VGND VPWR VPWR net430 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_94_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15020_ _13333_ _13420_ _13525_ _13357_ VGND VGND VPWR VPWR _13568_ sky130_fd_sc_hd__a31o_1
X_27006_ _11752_ VGND VGND VPWR VPWR _11889_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_161_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24218_ _09224_ net4136 _10279_ VGND VGND VPWR VPWR _10280_ sky130_fd_sc_hd__mux2_1
X_25198_ _10739_ net3114 _10829_ VGND VGND VPWR VPWR _10837_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16971_ _04737_ VGND VGND VPWR VPWR _01556_ sky130_fd_sc_hd__clkbuf_1
X_28957_ _12985_ VGND VGND VPWR VPWR _04261_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18710_ _05693_ _05864_ _05820_ VGND VGND VPWR VPWR _06063_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27908_ _12405_ VGND VGND VPWR VPWR _03792_ sky130_fd_sc_hd__clkbuf_1
X_15922_ _14296_ VGND VGND VPWR VPWR _02064_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_200_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19690_ _06916_ _06965_ _06984_ _06985_ VGND VGND VPWR VPWR _06986_ sky130_fd_sc_hd__a211o_1
X_28888_ _12948_ VGND VGND VPWR VPWR _04229_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18641_ _05425_ _05426_ VGND VGND VPWR VPWR _05997_ sky130_fd_sc_hd__or2_1
X_27839_ _12365_ net4323 _12357_ VGND VGND VPWR VPWR _12366_ sky130_fd_sc_hd__mux2_1
X_15853_ net2110 _13244_ _14258_ VGND VGND VPWR VPWR _14259_ sky130_fd_sc_hd__mux2_1
XFILLER_0_203_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_189_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_204_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14804_ _13356_ VGND VGND VPWR VPWR _13357_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_157_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18572_ _05368_ _05401_ _05366_ VGND VGND VPWR VPWR _05931_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30850_ clknet_leaf_221_clk _02585_ VGND VGND VPWR VPWR datamem.data_ram\[43\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_15784_ _14172_ net2567 _14221_ VGND VGND VPWR VPWR _14222_ sky130_fd_sc_hd__mux2_1
X_26503__55 clknet_1_1__leaf__11602_ VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__inv_2
XFILLER_0_87_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17523_ _05030_ VGND VGND VPWR VPWR _01281_ sky130_fd_sc_hd__clkbuf_1
X_29509_ net871 _01244_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[28\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_14735_ rvcpu.dp.pcreg.q\[3\] VGND VGND VPWR VPWR _13288_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_143_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30781_ clknet_leaf_154_clk _02516_ VGND VGND VPWR VPWR datamem.data_ram\[46\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_197_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32520_ clknet_leaf_4_clk _03942_ VGND VGND VPWR VPWR datamem.data_ram\[24\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_14666_ rvcpu.dp.plmw.ALUResultW\[14\] rvcpu.dp.plmw.ReadDataW\[14\] rvcpu.dp.plmw.PCPlus4W\[14\]
+ rvcpu.dp.plmw.lAuiPCW\[14\] _13192_ _13193_ VGND VGND VPWR VPWR _13234_ sky130_fd_sc_hd__mux4_2
XFILLER_0_184_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17454_ _14168_ net2388 _04985_ VGND VGND VPWR VPWR _04994_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23871__433 clknet_1_0__leaf__10220_ VGND VGND VPWR VPWR net559 sky130_fd_sc_hd__inv_2
XFILLER_0_129_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16405_ _14568_ VGND VGND VPWR VPWR _01837_ sky130_fd_sc_hd__clkbuf_1
X_32451_ clknet_leaf_248_clk _03873_ VGND VGND VPWR VPWR datamem.data_ram\[27\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14597_ net1898 _13173_ _13181_ VGND VGND VPWR VPWR _13182_ sky130_fd_sc_hd__mux2_1
X_17385_ _04957_ VGND VGND VPWR VPWR _01346_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_223_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19124_ _06441_ _06442_ VGND VGND VPWR VPWR _06443_ sky130_fd_sc_hd__and2_1
X_31402_ clknet_leaf_44_clk _03105_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCE\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16336_ net2816 _14434_ _14525_ VGND VGND VPWR VPWR _14532_ sky130_fd_sc_hd__mux2_1
XFILLER_0_229_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32382_ clknet_leaf_90_clk _03804_ VGND VGND VPWR VPWR datamem.data_ram\[2\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19055_ _06381_ _06382_ VGND VGND VPWR VPWR _06383_ sky130_fd_sc_hd__nor2_1
X_31333_ clknet_leaf_15_clk _03036_ VGND VGND VPWR VPWR rvcpu.dp.plde.RdE\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16267_ _14495_ VGND VGND VPWR VPWR _01902_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15218_ _13314_ _13758_ VGND VGND VPWR VPWR _13759_ sky130_fd_sc_hd__nor2_1
X_18006_ _05373_ VGND VGND VPWR VPWR _05376_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31264_ clknet_leaf_19_clk _02967_ VGND VGND VPWR VPWR rvcpu.dp.plfd.InstrD\[22\]
+ sky130_fd_sc_hd__dfxtp_2
Xclkbuf_1_0__f__10112_ clknet_0__10112_ VGND VGND VPWR VPWR clknet_1_0__leaf__10112_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_23_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16198_ _14450_ VGND VGND VPWR VPWR _01934_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15149_ _13297_ _13506_ VGND VGND VPWR VPWR _13693_ sky130_fd_sc_hd__nand2_1
X_30215_ net569 _01950_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[7\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31195_ clknet_leaf_46_clk _02898_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCPlus4D\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_207_5460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_207_5471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30146_ net508 _01881_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[0\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_19957_ datamem.data_ram\[58\]\[18\] _06692_ _07247_ _07250_ VGND VGND VPWR VPWR
+ _07251_ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18908_ _05240_ _06239_ _06242_ _06248_ VGND VGND VPWR VPWR rvcpu.ALUResultE\[23\]
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_208_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_203_5357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30077_ net439 _01812_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[11\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_203_5368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19888_ datamem.data_ram\[30\]\[17\] _06630_ _06665_ datamem.data_ram\[29\]\[17\]
+ VGND VGND VPWR VPWR _07183_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_203_5379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_5261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_5272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_5283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18839_ _05488_ _06183_ VGND VGND VPWR VPWR _06184_ sky130_fd_sc_hd__xnor2_1
X_23806__390 clknet_1_0__leaf__10206_ VGND VGND VPWR VPWR net516 sky130_fd_sc_hd__inv_2
XFILLER_0_222_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_195_5169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21850_ rvcpu.dp.rf.reg_file_arr\[4\]\[24\] rvcpu.dp.rf.reg_file_arr\[5\]\[24\] rvcpu.dp.rf.reg_file_arr\[6\]\[24\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[24\] _08839_ _08840_ VGND VGND VPWR VPWR _09088_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_171_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_214_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20801_ datamem.data_ram\[54\]\[30\] _06629_ _06783_ datamem.data_ram\[49\]\[30\]
+ _08090_ VGND VGND VPWR VPWR _08091_ sky130_fd_sc_hd__o221a_1
X_21781_ rvcpu.dp.rf.reg_file_arr\[16\]\[21\] rvcpu.dp.rf.reg_file_arr\[17\]\[21\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[21\] rvcpu.dp.rf.reg_file_arr\[19\]\[21\] _08703_
+ _08721_ VGND VGND VPWR VPWR _09022_ sky130_fd_sc_hd__mux4_1
X_30979_ clknet_leaf_160_clk _02714_ VGND VGND VPWR VPWR datamem.data_ram\[39\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23520_ _10168_ VGND VGND VPWR VPWR _01641_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_212_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20732_ _06623_ _08018_ _08021_ _07131_ VGND VGND VPWR VPWR _08022_ sky130_fd_sc_hd__a211o_1
X_32718_ clknet_leaf_284_clk _04140_ VGND VGND VPWR VPWR datamem.data_ram\[17\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_187_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_4290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_186_Right_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32649_ clknet_leaf_243_clk _04071_ VGND VGND VPWR VPWR datamem.data_ram\[19\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_20663_ datamem.data_ram\[58\]\[29\] _06802_ _06812_ datamem.data_ram\[59\]\[29\]
+ _06599_ VGND VGND VPWR VPWR _07954_ sky130_fd_sc_hd__o221a_1
XFILLER_0_133_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_4187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_4198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22402_ rvcpu.dp.rf.reg_file_arr\[24\]\[5\] rvcpu.dp.rf.reg_file_arr\[25\]\[5\] rvcpu.dp.rf.reg_file_arr\[26\]\[5\]
+ rvcpu.dp.rf.reg_file_arr\[27\]\[5\] _09484_ _09431_ VGND VGND VPWR VPWR _09563_
+ sky130_fd_sc_hd__mux4_1
X_26170_ _09479_ _11362_ VGND VGND VPWR VPWR _11422_ sky130_fd_sc_hd__and2_1
XFILLER_0_162_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20594_ datamem.data_ram\[21\]\[13\] _06664_ _07020_ datamem.data_ram\[23\]\[13\]
+ _07884_ VGND VGND VPWR VPWR _07885_ sky130_fd_sc_hd__o221a_1
XFILLER_0_162_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25121_ _10739_ net2364 _10784_ VGND VGND VPWR VPWR _10792_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22333_ _09495_ _09496_ VGND VGND VPWR VPWR _09497_ sky130_fd_sc_hd__nor2_1
XFILLER_0_190_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_4504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_4515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25052_ _10753_ VGND VGND VPWR VPWR _02588_ sky130_fd_sc_hd__clkbuf_1
X_22264_ _08595_ VGND VGND VPWR VPWR _09430_ sky130_fd_sc_hd__buf_4
XFILLER_0_60_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21215_ _08487_ _07597_ _08490_ VGND VGND VPWR VPWR _04425_ sky130_fd_sc_hd__o21ai_1
X_24166__8 clknet_1_1__leaf__10264_ VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__inv_2
XFILLER_0_143_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29860_ net238 _01595_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[18\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_22195_ _09260_ net4221 _09362_ VGND VGND VPWR VPWR _09370_ sky130_fd_sc_hd__mux2_1
X_28811_ _12692_ net3079 _12905_ VGND VGND VPWR VPWR _12908_ sky130_fd_sc_hd__mux2_1
X_21146_ _08430_ _08434_ _07872_ VGND VGND VPWR VPWR _08435_ sky130_fd_sc_hd__a21o_1
XFILLER_0_228_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29791_ net1137 _01526_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[20\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_126_3511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_3522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28742_ _12739_ net2995 net41 VGND VGND VPWR VPWR _12871_ sky130_fd_sc_hd__mux2_1
X_25954_ net1808 _11155_ VGND VGND VPWR VPWR _11299_ sky130_fd_sc_hd__or2_1
X_21077_ _07823_ datamem.data_ram\[43\]\[7\] _07874_ datamem.data_ram\[42\]\[7\] rvcpu.dp.plem.ALUResultM\[3\]
+ VGND VGND VPWR VPWR _08366_ sky130_fd_sc_hd__o221a_1
XFILLER_0_219_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20028_ _07299_ _07321_ VGND VGND VPWR VPWR _07322_ sky130_fd_sc_hd__nand2_1
X_24905_ _10670_ VGND VGND VPWR VPWR _02524_ sky130_fd_sc_hd__clkbuf_1
X_25885_ net1364 _11256_ _11258_ _11259_ VGND VGND VPWR VPWR _02915_ sky130_fd_sc_hd__o211a_1
X_28673_ _12834_ VGND VGND VPWR VPWR _04128_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_122_3419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27624_ _12089_ net2761 net80 VGND VGND VPWR VPWR _12247_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_87_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24836_ _10442_ net3639 _10631_ VGND VGND VPWR VPWR _10633_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27555_ _12210_ VGND VGND VPWR VPWR _03634_ sky130_fd_sc_hd__clkbuf_1
X_24767_ _10593_ VGND VGND VPWR VPWR _02463_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_201_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21979_ _08523_ _09207_ _09209_ _08558_ VGND VGND VPWR VPWR _09210_ sky130_fd_sc_hd__o211a_1
XFILLER_0_197_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27486_ _12173_ VGND VGND VPWR VPWR _03602_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24698_ _10556_ VGND VGND VPWR VPWR _02431_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0__10106_ _10106_ VGND VGND VPWR VPWR clknet_0__10106_ sky130_fd_sc_hd__clkbuf_16
X_29225_ _12601_ _09301_ _09230_ VGND VGND VPWR VPWR _13132_ sky130_fd_sc_hd__a21oi_4
X_26437_ _06478_ _11539_ _11529_ _11199_ _11568_ VGND VGND VPWR VPWR _11569_ sky130_fd_sc_hd__a221o_1
XFILLER_0_181_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_153_Right_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17170_ _04843_ VGND VGND VPWR VPWR _01455_ sky130_fd_sc_hd__clkbuf_1
X_26368_ _11517_ net1512 _11510_ _11518_ VGND VGND VPWR VPWR _03139_ sky130_fd_sc_hd__a31o_1
XFILLER_0_153_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29156_ _09223_ net4244 net64 VGND VGND VPWR VPWR _13095_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16121_ net2166 _13232_ _14396_ VGND VGND VPWR VPWR _14403_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23404__1019 clknet_1_1__leaf__10140_ VGND VGND VPWR VPWR net1145 sky130_fd_sc_hd__inv_2
X_25319_ _10904_ VGND VGND VPWR VPWR _02704_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28107_ _12518_ VGND VGND VPWR VPWR _03878_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26299_ _11482_ VGND VGND VPWR VPWR _03106_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_130_clk clknet_5_31__leaf_clk VGND VGND VPWR VPWR clknet_leaf_130_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_51_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29087_ _10979_ _11123_ _12977_ VGND VGND VPWR VPWR _13058_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_84_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16052_ _14366_ VGND VGND VPWR VPWR _01996_ sky130_fd_sc_hd__clkbuf_1
X_28038_ _12481_ VGND VGND VPWR VPWR _03846_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15003_ _13509_ _13507_ _13550_ VGND VGND VPWR VPWR _13551_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_55_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22959__668 clknet_1_0__leaf__10081_ VGND VGND VPWR VPWR net794 sky130_fd_sc_hd__inv_2
XFILLER_0_103_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30000_ net370 _01735_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[14\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_19811_ _06603_ _07098_ _07100_ _07105_ VGND VGND VPWR VPWR _07106_ sky130_fd_sc_hd__a31o_1
XFILLER_0_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29989_ net359 _01724_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[14\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_24120__626 clknet_1_0__leaf__10260_ VGND VGND VPWR VPWR net752 sky130_fd_sc_hd__inv_2
XFILLER_0_202_1277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19742_ _06823_ VGND VGND VPWR VPWR _07037_ sky130_fd_sc_hd__buf_6
X_16954_ _04728_ VGND VGND VPWR VPWR _01564_ sky130_fd_sc_hd__clkbuf_1
X_15905_ net2336 _13217_ _14286_ VGND VGND VPWR VPWR _14288_ sky130_fd_sc_hd__mux2_1
X_19673_ _06920_ VGND VGND VPWR VPWR _06969_ sky130_fd_sc_hd__buf_4
X_31951_ clknet_leaf_119_clk _03373_ VGND VGND VPWR VPWR datamem.data_ram\[55\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_197_clk clknet_5_29__leaf_clk VGND VGND VPWR VPWR clknet_leaf_197_clk
+ sky130_fd_sc_hd__clkbuf_8
X_16885_ net4381 _14436_ _04684_ VGND VGND VPWR VPWR _04692_ sky130_fd_sc_hd__mux2_1
XFILLER_0_218_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18624_ _05345_ _05784_ VGND VGND VPWR VPWR _05981_ sky130_fd_sc_hd__nor2_1
X_30902_ clknet_leaf_222_clk _02637_ VGND VGND VPWR VPWR datamem.data_ram\[41\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15836_ net2116 _13220_ _14247_ VGND VGND VPWR VPWR _14250_ sky130_fd_sc_hd__mux2_1
X_31882_ clknet_leaf_111_clk _03336_ VGND VGND VPWR VPWR datamem.data_ram\[57\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_220_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_205_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18555_ _05870_ _05914_ _05688_ VGND VGND VPWR VPWR _05915_ sky130_fd_sc_hd__mux2_1
X_30833_ clknet_leaf_152_clk _02568_ VGND VGND VPWR VPWR datamem.data_ram\[44\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_15767_ _14156_ net2625 _14210_ VGND VGND VPWR VPWR _14213_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_190_5044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17506_ _13213_ net2923 _05021_ VGND VGND VPWR VPWR _05022_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_190_5055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14718_ _13273_ VGND VGND VPWR VPWR _03174_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30764_ clknet_leaf_135_clk _02499_ VGND VGND VPWR VPWR datamem.data_ram\[47\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_18486_ _05349_ _05663_ VGND VGND VPWR VPWR _05848_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_190_5066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15698_ _14169_ VGND VGND VPWR VPWR _02169_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_480 _09317_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_491 _09750_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32503_ clknet_leaf_275_clk _03925_ VGND VGND VPWR VPWR datamem.data_ram\[25\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_16_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17437_ _04973_ VGND VGND VPWR VPWR _04985_ sky130_fd_sc_hd__buf_4
XFILLER_0_185_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14649_ _13221_ VGND VGND VPWR VPWR _03191_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_16_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30695_ clknet_leaf_153_clk _02430_ VGND VGND VPWR VPWR datamem.data_ram\[4\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_120_Right_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_16 _06612_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_27 _06633_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32434_ clknet_leaf_238_clk _03856_ VGND VGND VPWR VPWR datamem.data_ram\[27\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_38 _06676_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_49 _06681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17368_ _04948_ VGND VGND VPWR VPWR _01354_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19107_ rvcpu.dp.plde.ImmExtE\[12\] rvcpu.dp.plde.PCE\[12\] VGND VGND VPWR VPWR _06428_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_172_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16319_ _14522_ VGND VGND VPWR VPWR _01877_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_121_clk clknet_5_30__leaf_clk VGND VGND VPWR VPWR clknet_leaf_121_clk
+ sky130_fd_sc_hd__clkbuf_8
X_32365_ clknet_leaf_94_clk _03787_ VGND VGND VPWR VPWR datamem.data_ram\[2\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_17299_ rvcpu.dp.rf.reg_file_arr\[24\]\[22\] _13209_ _04902_ VGND VGND VPWR VPWR
+ _04912_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_209_5500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_209_5511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19038_ rvcpu.dp.plde.ImmExtE\[3\] rvcpu.dp.plde.PCE\[3\] VGND VGND VPWR VPWR _06368_
+ sky130_fd_sc_hd__or2_1
X_31316_ clknet_leaf_28_clk _03019_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCPlus4E\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_209_5522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32296_ clknet_leaf_201_clk _03718_ VGND VGND VPWR VPWR datamem.data_ram\[32\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31247_ clknet_leaf_21_clk _02950_ VGND VGND VPWR VPWR rvcpu.c.ad.opb5 sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_205_5408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_205_5419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21000_ datamem.data_ram\[29\]\[15\] _06660_ _08288_ _08124_ VGND VGND VPWR VPWR
+ _08289_ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31178_ clknet_leaf_216_clk _02881_ VGND VGND VPWR VPWR datamem.data_ram\[5\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2903 datamem.data_ram\[6\]\[16\] VGND VGND VPWR VPWR net4053 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2914 datamem.data_ram\[61\]\[21\] VGND VGND VPWR VPWR net4064 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2925 datamem.data_ram\[7\]\[29\] VGND VGND VPWR VPWR net4075 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2936 datamem.data_ram\[41\]\[9\] VGND VGND VPWR VPWR net4086 sky130_fd_sc_hd__dlygate4sd3_1
X_30129_ net491 _01864_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[10\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2947 datamem.data_ram\[28\]\[15\] VGND VGND VPWR VPWR net4097 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2958 datamem.data_ram\[1\]\[8\] VGND VGND VPWR VPWR net4108 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2969 datamem.data_ram\[52\]\[7\] VGND VGND VPWR VPWR net4119 sky130_fd_sc_hd__dlygate4sd3_1
X_22951_ _10056_ net1392 _10046_ _10077_ VGND VGND VPWR VPWR _01163_ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_188_clk clknet_5_22__leaf_clk VGND VGND VPWR VPWR clknet_leaf_188_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_177_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21902_ _08813_ _09136_ _08579_ VGND VGND VPWR VPWR _09137_ sky130_fd_sc_hd__a21o_1
X_25670_ _11085_ net1696 _11097_ _11103_ VGND VGND VPWR VPWR _02856_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_3_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23878__439 clknet_1_0__leaf__10221_ VGND VGND VPWR VPWR net565 sky130_fd_sc_hd__inv_2
X_22882_ rvcpu.dp.rf.reg_file_arr\[8\]\[30\] rvcpu.dp.rf.reg_file_arr\[10\]\[30\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[30\] rvcpu.dp.rf.reg_file_arr\[11\]\[30\] _09483_
+ _09656_ VGND VGND VPWR VPWR _10018_ sky130_fd_sc_hd__mux4_1
XFILLER_0_218_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24621_ _10513_ VGND VGND VPWR VPWR _02397_ sky130_fd_sc_hd__clkbuf_1
X_21833_ _08842_ _09071_ VGND VGND VPWR VPWR _09072_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_156_4238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27340_ _09309_ VGND VGND VPWR VPWR _12085_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_156_4249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24552_ _09317_ VGND VGND VPWR VPWR _10474_ sky130_fd_sc_hd__clkbuf_2
X_21764_ rvcpu.dp.rf.reg_file_arr\[20\]\[20\] rvcpu.dp.rf.reg_file_arr\[21\]\[20\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[20\] rvcpu.dp.rf.reg_file_arr\[23\]\[20\] _08516_
+ _08518_ VGND VGND VPWR VPWR _09006_ sky130_fd_sc_hd__mux4_2
XFILLER_0_37_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_704 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20715_ datamem.data_ram\[22\]\[5\] _06952_ _06969_ datamem.data_ram\[21\]\[5\] _06810_
+ VGND VGND VPWR VPWR _08006_ sky130_fd_sc_hd__a221o_1
X_27271_ _10818_ net3429 _12043_ VGND VGND VPWR VPWR _12047_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24483_ _09306_ datamem.data_ram\[52\]\[25\] _10430_ VGND VGND VPWR VPWR _10432_
+ sky130_fd_sc_hd__mux2_1
X_21695_ _08523_ _08940_ _08748_ VGND VGND VPWR VPWR _08941_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_149_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29010_ _10069_ _13010_ VGND VGND VPWR VPWR _13016_ sky130_fd_sc_hd__and2_1
X_26222_ net1300 _11371_ _11444_ VGND VGND VPWR VPWR _11449_ sky130_fd_sc_hd__and3_1
XFILLER_0_135_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20646_ datamem.data_ram\[29\]\[29\] _06823_ _06807_ datamem.data_ram\[24\]\[29\]
+ VGND VGND VPWR VPWR _07937_ sky130_fd_sc_hd__o22a_1
XFILLER_0_34_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26153_ _08622_ VGND VGND VPWR VPWR _11413_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_115_3245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_112_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_112_clk
+ sky130_fd_sc_hd__clkbuf_8
X_20577_ _07867_ VGND VGND VPWR VPWR _07868_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_115_3256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25104_ _10075_ VGND VGND VPWR VPWR _10783_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_46_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_225_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22316_ _09390_ VGND VGND VPWR VPWR _09481_ sky130_fd_sc_hd__buf_2
X_26084_ rvcpu.dp.plfd.InstrD\[6\] _11374_ _06572_ VGND VGND VPWR VPWR _11375_ sky130_fd_sc_hd__and3b_1
XFILLER_0_21_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_186_4957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_186_4968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29912_ net282 _01647_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[16\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_25035_ _10468_ net3280 net90 VGND VGND VPWR VPWR _10744_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22247_ _08589_ VGND VGND VPWR VPWR _09413_ sky130_fd_sc_hd__clkbuf_4
X_29843_ net221 _01578_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[18\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_22178_ _09360_ VGND VGND VPWR VPWR _01107_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_218_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21129_ _07839_ _08417_ VGND VGND VPWR VPWR _08418_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_50_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29774_ net1120 _01509_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[20\]\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_89_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26986_ _11877_ VGND VGND VPWR VPWR _03398_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_89_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_3964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28725_ _12756_ net3255 _12859_ VGND VGND VPWR VPWR _12862_ sky130_fd_sc_hd__mux2_1
X_25937_ _11289_ VGND VGND VPWR VPWR _11290_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_145_3986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_179_clk clknet_5_19__leaf_clk VGND VGND VPWR VPWR clknet_leaf_179_clk
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_222_Right_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_214_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24193__33 clknet_1_1__leaf__10266_ VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__inv_2
XFILLER_0_92_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16670_ _04578_ VGND VGND VPWR VPWR _01706_ sky130_fd_sc_hd__clkbuf_1
X_28656_ _12825_ VGND VGND VPWR VPWR _04120_ sky130_fd_sc_hd__clkbuf_1
X_25868_ _11246_ VGND VGND VPWR VPWR _02911_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15621_ net4253 _13257_ _14114_ VGND VGND VPWR VPWR _14119_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27607_ _12151_ net2586 net81 VGND VGND VPWR VPWR _12238_ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24819_ _10623_ VGND VGND VPWR VPWR _02485_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28587_ _12788_ VGND VGND VPWR VPWR _04088_ sky130_fd_sc_hd__clkbuf_1
X_25799_ rvcpu.dp.pcreg.q\[16\] _11188_ VGND VGND VPWR VPWR _11191_ sky130_fd_sc_hd__and2_1
XFILLER_0_124_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18340_ _05704_ VGND VGND VPWR VPWR _05705_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15552_ _13467_ _13462_ _13878_ VGND VGND VPWR VPWR _14076_ sky130_fd_sc_hd__a21oi_1
X_27538_ _12201_ VGND VGND VPWR VPWR _03626_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_104_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15483_ _13542_ _13824_ _14011_ _13994_ _13600_ VGND VGND VPWR VPWR _14012_ sky130_fd_sc_hd__a32o_1
X_18271_ rvcpu.dp.plde.RD1E\[27\] _05564_ _05538_ VGND VGND VPWR VPWR _05636_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_13_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27469_ _12089_ net3470 net83 VGND VGND VPWR VPWR _12164_ sky130_fd_sc_hd__mux2_1
XFILLER_0_194_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29208_ _10042_ _10947_ VGND VGND VPWR VPWR _13123_ sky130_fd_sc_hd__nor2_2
X_17222_ _14141_ net2221 _04865_ VGND VGND VPWR VPWR _04871_ sky130_fd_sc_hd__mux2_1
X_30480_ net158 _02215_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[19\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29139_ _09266_ net3032 net39 VGND VGND VPWR VPWR _13086_ sky130_fd_sc_hd__mux2_1
X_17153_ _04834_ VGND VGND VPWR VPWR _01463_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_103_clk clknet_5_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_103_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_52_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16104_ net2211 _13207_ _14385_ VGND VGND VPWR VPWR _14394_ sky130_fd_sc_hd__mux2_1
X_32150_ clknet_leaf_230_clk _03572_ VGND VGND VPWR VPWR datamem.data_ram\[38\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_17084_ _14139_ net4425 _04793_ VGND VGND VPWR VPWR _04798_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold809 rvcpu.dp.rf.reg_file_arr\[0\]\[1\] VGND VGND VPWR VPWR net1959 sky130_fd_sc_hd__dlygate4sd3_1
X_31101_ clknet_leaf_108_clk _02836_ VGND VGND VPWR VPWR datamem.data_ram\[19\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16035_ _14357_ VGND VGND VPWR VPWR _02004_ sky130_fd_sc_hd__clkbuf_1
X_32081_ clknet_leaf_63_clk _03503_ VGND VGND VPWR VPWR datamem.data_ram\[47\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31032_ clknet_leaf_102_clk _02767_ VGND VGND VPWR VPWR datamem.data_ram\[12\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_229_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17986_ _05354_ _05355_ VGND VGND VPWR VPWR _05356_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_200_5305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1509 rvcpu.dp.rf.reg_file_arr\[21\]\[0\] VGND VGND VPWR VPWR net2659 sky130_fd_sc_hd__dlygate4sd3_1
X_19725_ _06784_ VGND VGND VPWR VPWR _07020_ sky130_fd_sc_hd__buf_6
XFILLER_0_100_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16937_ _13179_ _14234_ VGND VGND VPWR VPWR _04719_ sky130_fd_sc_hd__nor2_2
X_32983_ clknet_leaf_174_clk _04405_ VGND VGND VPWR VPWR datamem.data_ram\[63\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31934_ clknet_leaf_113_clk _03356_ VGND VGND VPWR VPWR datamem.data_ram\[60\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_19656_ _06951_ VGND VGND VPWR VPWR _06952_ sky130_fd_sc_hd__buf_4
X_23265__911 clknet_1_1__leaf__10128_ VGND VGND VPWR VPWR net1037 sky130_fd_sc_hd__inv_2
XFILLER_0_79_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_192_5106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16868_ _04682_ VGND VGND VPWR VPWR _01604_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_205_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18607_ _05349_ _05664_ _05851_ VGND VGND VPWR VPWR _05965_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_177_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15819_ net2019 _13195_ _14236_ VGND VGND VPWR VPWR _14241_ sky130_fd_sc_hd__mux2_1
X_31865_ clknet_leaf_122_clk _03319_ VGND VGND VPWR VPWR datamem.data_ram\[63\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_19587_ datamem.data_ram\[46\]\[8\] _06743_ _06661_ datamem.data_ram\[45\]\[8\] _06882_
+ VGND VGND VPWR VPWR _06883_ sky130_fd_sc_hd__o221a_1
X_16799_ net2723 _14486_ _04611_ VGND VGND VPWR VPWR _04646_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18538_ _05704_ _05896_ _05898_ _05692_ VGND VGND VPWR VPWR _05899_ sky130_fd_sc_hd__a211o_1
X_30816_ clknet_leaf_259_clk _02551_ VGND VGND VPWR VPWR datamem.data_ram\[45\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_31796_ clknet_leaf_214_clk _03250_ VGND VGND VPWR VPWR datamem.data_ram\[2\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30747_ clknet_leaf_135_clk _02482_ VGND VGND VPWR VPWR datamem.data_ram\[48\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_18469_ _05313_ _05320_ _05506_ _05334_ _05579_ _05663_ VGND VGND VPWR VPWR _05832_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_157_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_4113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20500_ _07021_ VGND VGND VPWR VPWR _07791_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_151_4124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21480_ rvcpu.dp.rf.reg_file_arr\[0\]\[5\] rvcpu.dp.rf.reg_file_arr\[1\]\[5\] rvcpu.dp.rf.reg_file_arr\[2\]\[5\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[5\] _08566_ _08569_ VGND VGND VPWR VPWR _08737_ sky130_fd_sc_hd__mux4_1
X_30678_ clknet_leaf_96_clk _02413_ VGND VGND VPWR VPWR datamem.data_ram\[4\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32417_ clknet_leaf_76_clk _03839_ VGND VGND VPWR VPWR datamem.data_ram\[28\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20431_ datamem.data_ram\[15\]\[12\] _06784_ _07722_ _06601_ VGND VGND VPWR VPWR
+ _07723_ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23150_ clknet_1_0__leaf__10079_ VGND VGND VPWR VPWR _10108_ sky130_fd_sc_hd__buf_1
XFILLER_0_71_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload230 clknet_leaf_109_clk VGND VGND VPWR VPWR clkload230/Y sky130_fd_sc_hd__clkinv_1
X_32348_ clknet_leaf_169_clk _03770_ VGND VGND VPWR VPWR datamem.data_ram\[30\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20362_ datamem.data_ram\[0\]\[28\] _06695_ _06730_ datamem.data_ram\[3\]\[28\] _06678_
+ VGND VGND VPWR VPWR _07654_ sky130_fd_sc_hd__o221a_1
Xclkload241 clknet_leaf_123_clk VGND VGND VPWR VPWR clkload241/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_0_130_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload252 clknet_leaf_190_clk VGND VGND VPWR VPWR clkload252/Y sky130_fd_sc_hd__inv_6
X_22101_ rvcpu.dp.plem.WriteDataM\[3\] _08488_ _09293_ VGND VGND VPWR VPWR _09312_
+ sky130_fd_sc_hd__and3_1
Xclkload263 clknet_leaf_196_clk VGND VGND VPWR VPWR clkload263/Y sky130_fd_sc_hd__clkinv_8
XTAP_TAPCELL_ROW_228_5964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload274 clknet_leaf_129_clk VGND VGND VPWR VPWR clkload274/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_3_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_228_5975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_110_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32279_ clknet_leaf_89_clk _03701_ VGND VGND VPWR VPWR datamem.data_ram\[33\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_20293_ datamem.data_ram\[13\]\[19\] _06662_ _06646_ datamem.data_ram\[8\]\[19\]
+ VGND VGND VPWR VPWR _07586_ sky130_fd_sc_hd__o22a_1
Xclkload285 clknet_1_0__leaf__10224_ VGND VGND VPWR VPWR clkload285/X sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_110_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_4064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload296 clknet_1_0__leaf__10220_ VGND VGND VPWR VPWR clkload296/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_149_4075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22032_ _09255_ VGND VGND VPWR VPWR _09256_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_140_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_181_4832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_181_4843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2700 datamem.data_ram\[19\]\[13\] VGND VGND VPWR VPWR net3850 sky130_fd_sc_hd__dlygate4sd3_1
X_26840_ _11679_ _11786_ VGND VGND VPWR VPWR _11788_ sky130_fd_sc_hd__and2_1
Xhold2711 datamem.data_ram\[11\]\[21\] VGND VGND VPWR VPWR net3861 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2722 rvcpu.dp.rf.reg_file_arr\[25\]\[4\] VGND VGND VPWR VPWR net3872 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_71_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2733 rvcpu.dp.rf.reg_file_arr\[5\]\[29\] VGND VGND VPWR VPWR net3883 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2744 rvcpu.dp.rf.reg_file_arr\[23\]\[6\] VGND VGND VPWR VPWR net3894 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2755 datamem.data_ram\[35\]\[24\] VGND VGND VPWR VPWR net3905 sky130_fd_sc_hd__dlygate4sd3_1
X_26771_ _11735_ net1856 _11737_ _11745_ VGND VGND VPWR VPWR _03315_ sky130_fd_sc_hd__a31o_1
Xhold2766 datamem.data_ram\[55\]\[9\] VGND VGND VPWR VPWR net3916 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2777 datamem.data_ram\[49\]\[21\] VGND VGND VPWR VPWR net3927 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2788 rvcpu.dp.rf.reg_file_arr\[30\]\[31\] VGND VGND VPWR VPWR net3938 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2799 datamem.data_ram\[53\]\[19\] VGND VGND VPWR VPWR net3949 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28510_ _12741_ net3701 net43 VGND VGND VPWR VPWR _12742_ sky130_fd_sc_hd__mux2_1
X_23403__1018 clknet_1_0__leaf__10140_ VGND VGND VPWR VPWR net1144 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_108_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22934_ _10064_ _10053_ VGND VGND VPWR VPWR _10065_ sky130_fd_sc_hd__and2_1
X_25722_ _10814_ net3020 _11133_ VGND VGND VPWR VPWR _11135_ sky130_fd_sc_hd__mux2_1
X_29490_ net852 _01225_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[2\]\[29\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_84_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_3850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_140_3861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28441_ _12701_ VGND VGND VPWR VPWR _04029_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_210_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25653_ _10064_ _11094_ _11095_ net1327 VGND VGND VPWR VPWR _02847_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_179_4783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22865_ _09481_ _10001_ VGND VGND VPWR VPWR _10002_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_179_4794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23127__804 clknet_1_0__leaf__10105_ VGND VGND VPWR VPWR net930 sky130_fd_sc_hd__inv_2
XFILLER_0_39_805 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24604_ _10504_ VGND VGND VPWR VPWR _02389_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21816_ _08672_ _09047_ _09051_ _09055_ VGND VGND VPWR VPWR _09056_ sky130_fd_sc_hd__and4_1
X_25584_ _08124_ _07177_ VGND VGND VPWR VPWR _11054_ sky130_fd_sc_hd__nor2_1
X_28372_ _12661_ VGND VGND VPWR VPWR _04000_ sky130_fd_sc_hd__clkbuf_1
X_22796_ rvcpu.dp.rf.reg_file_arr\[16\]\[26\] rvcpu.dp.rf.reg_file_arr\[17\]\[26\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[26\] rvcpu.dp.rf.reg_file_arr\[19\]\[26\] _09445_
+ _09447_ VGND VGND VPWR VPWR _09936_ sky130_fd_sc_hd__mux4_1
Xwire82 _12215_ VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__buf_4
XFILLER_0_167_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27323_ _10048_ _12076_ _12077_ net1406 VGND VGND VPWR VPWR _03535_ sky130_fd_sc_hd__a22o_1
XFILLER_0_183_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24535_ _10398_ net4419 _10456_ VGND VGND VPWR VPWR _10463_ sky130_fd_sc_hd__mux2_1
X_21747_ rvcpu.dp.rf.reg_file_arr\[28\]\[19\] rvcpu.dp.rf.reg_file_arr\[30\]\[19\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[19\] rvcpu.dp.rf.reg_file_arr\[31\]\[19\] _08559_
+ _08636_ VGND VGND VPWR VPWR _08990_ sky130_fd_sc_hd__mux4_1
XFILLER_0_4_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_3307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27254_ _07791_ _10043_ _10600_ VGND VGND VPWR VPWR _12041_ sky130_fd_sc_hd__nor3_1
XFILLER_0_136_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24466_ _09306_ net3911 _10421_ VGND VGND VPWR VPWR _10423_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21678_ _08795_ _08918_ _08920_ _08924_ _08808_ VGND VGND VPWR VPWR _08925_ sky130_fd_sc_hd__a311o_1
XFILLER_0_188_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_184_1011 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26205_ _11361_ _11379_ VGND VGND VPWR VPWR _11441_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27185_ _11991_ net1661 _11995_ _12000_ VGND VGND VPWR VPWR _03474_ sky130_fd_sc_hd__a31o_1
X_20629_ _07871_ _07893_ _07919_ VGND VGND VPWR VPWR _07920_ sky130_fd_sc_hd__a21oi_4
X_24397_ _09273_ net3954 _10376_ VGND VGND VPWR VPWR _10378_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_184_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26136_ net1844 _11397_ VGND VGND VPWR VPWR _11404_ sky130_fd_sc_hd__and2_1
XFILLER_0_62_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26067_ _11363_ VGND VGND VPWR VPWR _02993_ sky130_fd_sc_hd__buf_2
XFILLER_0_104_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25018_ _10732_ VGND VGND VPWR VPWR _02575_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_218_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23746__336 clknet_1_1__leaf__10200_ VGND VGND VPWR VPWR net462 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_37_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17840_ _13225_ rvcpu.dp.plde.RD2E\[17\] _05195_ VGND VGND VPWR VPWR _05221_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29826_ net204 _01561_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[1\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17771_ rvcpu.dp.plem.RdM\[3\] rvcpu.dp.plde.Rs2E\[3\] VGND VGND VPWR VPWR _05169_
+ sky130_fd_sc_hd__nor2_1
X_29757_ net1103 _01492_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[21\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_14983_ _13301_ _13434_ VGND VGND VPWR VPWR _13531_ sky130_fd_sc_hd__nor2_2
X_26969_ _11863_ net2049 _11865_ _11868_ VGND VGND VPWR VPWR _03390_ sky130_fd_sc_hd__a31o_1
X_19510_ _06805_ VGND VGND VPWR VPWR _06806_ sky130_fd_sc_hd__buf_6
X_16722_ _04605_ VGND VGND VPWR VPWR _01681_ sky130_fd_sc_hd__clkbuf_1
X_28708_ _12692_ net2713 _12850_ VGND VGND VPWR VPWR _12853_ sky130_fd_sc_hd__mux2_1
XFILLER_0_191_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29688_ net1034 _01423_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[23\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19441_ _06730_ VGND VGND VPWR VPWR _06737_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_202_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16653_ _14185_ net4105 _04562_ VGND VGND VPWR VPWR _04569_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_18_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28639_ _12816_ VGND VGND VPWR VPWR _04112_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_18_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_215_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15604_ net2589 _13232_ _14103_ VGND VGND VPWR VPWR _14110_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31650_ clknet_leaf_24_clk net1221 VGND VGND VPWR VPWR rvcpu.dp.plmw.lAuiPCW\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_19372_ _06667_ VGND VGND VPWR VPWR _06668_ sky130_fd_sc_hd__buf_4
X_16584_ _14185_ net3355 _04525_ VGND VGND VPWR VPWR _04532_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_201_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18323_ _05579_ VGND VGND VPWR VPWR _05688_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30601_ clknet_leaf_219_clk _02336_ VGND VGND VPWR VPWR datamem.data_ram\[53\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_15535_ _13398_ _13546_ _13872_ VGND VGND VPWR VPWR _14061_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_151_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_201_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31581_ clknet_leaf_71_clk datamem.rd_data_mem\[31\] VGND VGND VPWR VPWR rvcpu.dp.plmw.ReadDataW\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18254_ _05573_ _05618_ _05481_ VGND VGND VPWR VPWR _05619_ sky130_fd_sc_hd__a21oi_2
X_30532_ clknet_leaf_175_clk _02267_ VGND VGND VPWR VPWR datamem.data_ram\[56\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_15466_ _13350_ _13995_ VGND VGND VPWR VPWR _13996_ sky130_fd_sc_hd__nand2_1
XFILLER_0_167_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17205_ _04861_ VGND VGND VPWR VPWR _01438_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23295__937 clknet_1_0__leaf__10132_ VGND VGND VPWR VPWR net1063 sky130_fd_sc_hd__inv_2
X_18185_ _05531_ _05537_ _05543_ _05549_ VGND VGND VPWR VPWR _05550_ sky130_fd_sc_hd__and4_1
X_30463_ net141 _02198_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[19\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_15397_ _13378_ _13929_ _13590_ _13410_ VGND VGND VPWR VPWR _13930_ sky130_fd_sc_hd__a211o_1
XFILLER_0_163_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32202_ clknet_leaf_88_clk _03624_ VGND VGND VPWR VPWR datamem.data_ram\[36\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17136_ _14191_ net3097 _04815_ VGND VGND VPWR VPWR _04825_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold606 datamem.data_ram\[22\]\[6\] VGND VGND VPWR VPWR net1756 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30394_ net732 _02129_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[31\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_208_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold617 datamem.data_ram\[10\]\[7\] VGND VGND VPWR VPWR net1767 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24126__632 clknet_1_0__leaf__10260_ VGND VGND VPWR VPWR net758 sky130_fd_sc_hd__inv_2
Xhold628 datamem.data_ram\[26\]\[0\] VGND VGND VPWR VPWR net1778 sky130_fd_sc_hd__dlygate4sd3_1
X_32133_ clknet_leaf_234_clk _03555_ VGND VGND VPWR VPWR datamem.data_ram\[10\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold639 datamem.data_ram\[58\]\[0\] VGND VGND VPWR VPWR net1789 sky130_fd_sc_hd__dlygate4sd3_1
X_17067_ _04788_ VGND VGND VPWR VPWR _01503_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_204_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16018_ _14271_ _14347_ VGND VGND VPWR VPWR _14348_ sky130_fd_sc_hd__nor2_2
X_32064_ clknet_leaf_133_clk _03486_ VGND VGND VPWR VPWR datamem.data_ram\[48\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_209_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_223_5850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31015_ clknet_leaf_191_clk _02750_ VGND VGND VPWR VPWR datamem.data_ram\[42\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_5_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2007 datamem.data_ram\[53\]\[24\] VGND VGND VPWR VPWR net3157 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2018 rvcpu.dp.rf.reg_file_arr\[6\]\[17\] VGND VGND VPWR VPWR net3168 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2029 datamem.data_ram\[47\]\[25\] VGND VGND VPWR VPWR net3179 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1306 rvcpu.dp.rf.reg_file_arr\[18\]\[20\] VGND VGND VPWR VPWR net2456 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1317 datamem.data_ram\[36\]\[17\] VGND VGND VPWR VPWR net2467 sky130_fd_sc_hd__dlygate4sd3_1
X_17969_ _05294_ VGND VGND VPWR VPWR _05340_ sky130_fd_sc_hd__clkbuf_4
Xhold1328 datamem.data_ram\[45\]\[31\] VGND VGND VPWR VPWR net2478 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1339 rvcpu.dp.rf.reg_file_arr\[18\]\[15\] VGND VGND VPWR VPWR net2489 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19708_ datamem.data_ram\[23\]\[0\] _06926_ _06948_ datamem.data_ram\[17\]\[0\] VGND
+ VGND VPWR VPWR _07004_ sky130_fd_sc_hd__a22o_1
X_20980_ _08261_ _08268_ _07903_ VGND VGND VPWR VPWR _08269_ sky130_fd_sc_hd__a21o_1
X_32966_ clknet_leaf_207_clk _04388_ VGND VGND VPWR VPWR datamem.data_ram\[63\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_56 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31917_ _04429_ net120 VGND VGND VPWR VPWR datamem.rd_data_mem\[22\] sky130_fd_sc_hd__dlxtn_1
X_24172__14 clknet_1_0__leaf__10264_ VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__inv_2
X_19639_ _06933_ _06934_ VGND VGND VPWR VPWR _06935_ sky130_fd_sc_hd__nor2_8
XFILLER_0_178_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32897_ clknet_leaf_228_clk _04319_ VGND VGND VPWR VPWR datamem.data_ram\[0\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22650_ rvcpu.dp.rf.reg_file_arr\[16\]\[18\] rvcpu.dp.rf.reg_file_arr\[17\]\[18\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[18\] rvcpu.dp.rf.reg_file_arr\[19\]\[18\] _09384_
+ _09430_ VGND VGND VPWR VPWR _09798_ sky130_fd_sc_hd__mux4_1
XFILLER_0_94_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31848_ clknet_leaf_111_clk _03302_ VGND VGND VPWR VPWR datamem.data_ram\[61\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_193_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21601_ _08742_ _08851_ VGND VGND VPWR VPWR _08852_ sky130_fd_sc_hd__or2_1
XFILLER_0_165_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_217_5698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22581_ _09442_ _09728_ _09730_ _09732_ VGND VGND VPWR VPWR _09733_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_174_4680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31779_ clknet_leaf_262_clk _03233_ VGND VGND VPWR VPWR datamem.data_ram\[6\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24320_ _10335_ VGND VGND VPWR VPWR _02274_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21532_ _08511_ _08785_ VGND VGND VPWR VPWR _08786_ sky130_fd_sc_hd__nor2_1
XFILLER_0_146_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_4566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_170_4577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24251_ _07122_ VGND VGND VPWR VPWR _10297_ sky130_fd_sc_hd__buf_8
X_21463_ _08712_ _08716_ _08720_ _08625_ VGND VGND VPWR VPWR _01032_ sky130_fd_sc_hd__o31a_1
XFILLER_0_172_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23202_ _09256_ net2706 _10115_ VGND VGND VPWR VPWR _10122_ sky130_fd_sc_hd__mux2_1
X_20414_ datamem.data_ram\[63\]\[12\] _06705_ _07704_ _07705_ VGND VGND VPWR VPWR
+ _07706_ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21394_ rvcpu.dp.rf.reg_file_arr\[16\]\[2\] rvcpu.dp.rf.reg_file_arr\[17\]\[2\] rvcpu.dp.rf.reg_file_arr\[18\]\[2\]
+ rvcpu.dp.rf.reg_file_arr\[19\]\[2\] _08628_ _08629_ VGND VGND VPWR VPWR _08654_
+ sky130_fd_sc_hd__mux4_1
X_20345_ _07635_ datamem.data_ram\[59\]\[4\] _07636_ _06776_ VGND VGND VPWR VPWR _07637_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_4_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28990_ _13004_ VGND VGND VPWR VPWR _04275_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_73_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27941_ _12359_ net2327 _12421_ VGND VGND VPWR VPWR _12423_ sky130_fd_sc_hd__mux2_1
X_23064_ _09267_ net3658 _10093_ VGND VGND VPWR VPWR _10094_ sky130_fd_sc_hd__mux2_1
X_20276_ datamem.data_ram\[47\]\[19\] _06725_ _06765_ datamem.data_ram\[44\]\[19\]
+ VGND VGND VPWR VPWR _07569_ sky130_fd_sc_hd__o22a_1
XFILLER_0_12_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold3220 rvcpu.dp.rf.reg_file_arr\[21\]\[11\] VGND VGND VPWR VPWR net4370 sky130_fd_sc_hd__dlygate4sd3_1
X_22015_ rvcpu.dp.plem.WriteDataM\[19\] _09221_ VGND VGND VPWR VPWR _09242_ sky130_fd_sc_hd__and2_1
Xhold3231 rvcpu.dp.rf.reg_file_arr\[18\]\[24\] VGND VGND VPWR VPWR net4381 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3242 datamem.data_ram\[22\]\[23\] VGND VGND VPWR VPWR net4392 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_216_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold3253 rvcpu.dp.rf.reg_file_arr\[14\]\[11\] VGND VGND VPWR VPWR net4403 sky130_fd_sc_hd__dlygate4sd3_1
X_27872_ _12147_ net2997 net77 VGND VGND VPWR VPWR _12385_ sky130_fd_sc_hd__mux2_1
Xhold3264 datamem.data_ram\[5\]\[12\] VGND VGND VPWR VPWR net4414 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2530 datamem.data_ram\[12\]\[8\] VGND VGND VPWR VPWR net3680 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3275 rvcpu.dp.rf.reg_file_arr\[21\]\[27\] VGND VGND VPWR VPWR net4425 sky130_fd_sc_hd__dlygate4sd3_1
X_29611_ net965 _01346_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[25\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_26823_ _11767_ net1649 _11773_ _11777_ VGND VGND VPWR VPWR _03335_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_142_3901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3286 datamem.data_ram\[28\]\[20\] VGND VGND VPWR VPWR net4436 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2541 datamem.data_ram\[12\]\[12\] VGND VGND VPWR VPWR net3691 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3297 rvcpu.dp.plfd.InstrD\[10\] VGND VGND VPWR VPWR net4447 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2552 datamem.data_ram\[46\]\[12\] VGND VGND VPWR VPWR net3702 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2563 datamem.data_ram\[7\]\[23\] VGND VGND VPWR VPWR net3713 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2574 datamem.data_ram\[42\]\[17\] VGND VGND VPWR VPWR net3724 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1840 datamem.data_ram\[19\]\[20\] VGND VGND VPWR VPWR net2990 sky130_fd_sc_hd__dlygate4sd3_1
X_29542_ net896 _01277_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[27\]\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_32_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2585 datamem.data_ram\[27\]\[30\] VGND VGND VPWR VPWR net3735 sky130_fd_sc_hd__dlygate4sd3_1
X_26754_ _11104_ VGND VGND VPWR VPWR _11735_ sky130_fd_sc_hd__buf_2
XFILLER_0_216_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2596 datamem.data_ram\[50\]\[17\] VGND VGND VPWR VPWR net3746 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1851 rvcpu.dp.rf.reg_file_arr\[2\]\[22\] VGND VGND VPWR VPWR net3001 sky130_fd_sc_hd__dlygate4sd3_1
X_23966_ _09260_ net3787 _10229_ VGND VGND VPWR VPWR _10237_ sky130_fd_sc_hd__mux2_1
Xhold1862 datamem.data_ram\[35\]\[26\] VGND VGND VPWR VPWR net3012 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1873 datamem.data_ram\[47\]\[16\] VGND VGND VPWR VPWR net3023 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1884 datamem.data_ram\[26\]\[13\] VGND VGND VPWR VPWR net3034 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1895 rvcpu.dp.rf.reg_file_arr\[20\]\[24\] VGND VGND VPWR VPWR net3045 sky130_fd_sc_hd__dlygate4sd3_1
X_25705_ _10814_ net3880 _11124_ VGND VGND VPWR VPWR _11126_ sky130_fd_sc_hd__mux2_1
X_22917_ _10050_ VGND VGND VPWR VPWR _10051_ sky130_fd_sc_hd__buf_6
XFILLER_0_168_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29473_ net835 _01208_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[2\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_26685_ _11683_ net1697 _11693_ _11696_ VGND VGND VPWR VPWR _03278_ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28424_ _09305_ VGND VGND VPWR VPWR _12690_ sky130_fd_sc_hd__clkbuf_2
X_25636_ _11086_ _11079_ VGND VGND VPWR VPWR _11087_ sky130_fd_sc_hd__and2_1
X_22848_ _09461_ _09983_ _09985_ _09489_ VGND VGND VPWR VPWR _09986_ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_607 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28355_ _12652_ VGND VGND VPWR VPWR _03992_ sky130_fd_sc_hd__clkbuf_1
X_25567_ _10408_ _11042_ VGND VGND VPWR VPWR _11044_ sky130_fd_sc_hd__and2_1
XFILLER_0_149_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22779_ rvcpu.dp.rf.reg_file_arr\[20\]\[25\] rvcpu.dp.rf.reg_file_arr\[21\]\[25\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[25\] rvcpu.dp.rf.reg_file_arr\[23\]\[25\] _09434_
+ _09558_ VGND VGND VPWR VPWR _09920_ sky130_fd_sc_hd__mux4_1
X_27306_ _11968_ _12066_ VGND VGND VPWR VPWR _12068_ sky130_fd_sc_hd__and2_1
X_15320_ _13548_ _13847_ _13599_ VGND VGND VPWR VPWR _13857_ sky130_fd_sc_hd__a21o_1
XFILLER_0_148_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24518_ _10453_ VGND VGND VPWR VPWR _02354_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28286_ _12615_ VGND VGND VPWR VPWR _03960_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_136_3749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25498_ _10820_ net3397 _10999_ VGND VGND VPWR VPWR _11004_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15251_ _13329_ _13744_ _13483_ rvcpu.dp.pcreg.q\[8\] VGND VGND VPWR VPWR _13791_
+ sky130_fd_sc_hd__a211o_1
X_27237_ _11965_ _12031_ VGND VGND VPWR VPWR _12032_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24449_ _10055_ VGND VGND VPWR VPWR _10412_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_163_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15182_ _13554_ _13716_ _13724_ VGND VGND VPWR VPWR _13725_ sky130_fd_sc_hd__or3b_1
X_27168_ _11976_ _11984_ VGND VGND VPWR VPWR _11990_ sky130_fd_sc_hd__and2_1
X_23451__101 clknet_1_0__leaf__10156_ VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__inv_2
X_26119_ net1671 _11386_ VGND VGND VPWR VPWR _11395_ sky130_fd_sc_hd__and2_1
XFILLER_0_151_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19990_ datamem.data_ram\[4\]\[2\] _06953_ _06946_ datamem.data_ram\[1\]\[2\] VGND
+ VGND VPWR VPWR _07284_ sky130_fd_sc_hd__a22o_1
XFILLER_0_160_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27099_ _10066_ VGND VGND VPWR VPWR _11946_ sky130_fd_sc_hd__clkbuf_4
X_23980__515 clknet_1_1__leaf__10239_ VGND VGND VPWR VPWR net641 sky130_fd_sc_hd__inv_2
X_18941_ _05549_ _06278_ VGND VGND VPWR VPWR _06279_ sky130_fd_sc_hd__xor2_1
XFILLER_0_219_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18872_ _05694_ _06095_ VGND VGND VPWR VPWR _06215_ sky130_fd_sc_hd__nand2_1
XFILLER_0_197_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17823_ rvcpu.dp.plem.ALUResultM\[25\] _05209_ _05178_ VGND VGND VPWR VPWR _05210_
+ sky130_fd_sc_hd__mux2_1
X_29809_ net1147 _01544_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[1\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3 rvcpu.dp.plde.PCPlus4E\[19\] VGND VGND VPWR VPWR net1153 sky130_fd_sc_hd__dlygate4sd3_1
X_26513__1 clknet_1_1__leaf__10080_ VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__inv_2
X_32820_ clknet_leaf_233_clk _04242_ VGND VGND VPWR VPWR datamem.data_ram\[12\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17754_ _05152_ VGND VGND VPWR VPWR _01164_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_221_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14966_ _13511_ _13512_ _13514_ VGND VGND VPWR VPWR _13515_ sky130_fd_sc_hd__o21a_1
XFILLER_0_178_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16705_ _04596_ VGND VGND VPWR VPWR _01689_ sky130_fd_sc_hd__clkbuf_1
X_32751_ clknet_leaf_184_clk _04173_ VGND VGND VPWR VPWR datamem.data_ram\[15\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17685_ net2904 _13277_ _05081_ VGND VGND VPWR VPWR _05116_ sky130_fd_sc_hd__mux2_1
X_14897_ _13343_ _13447_ VGND VGND VPWR VPWR _13448_ sky130_fd_sc_hd__nand2_1
XFILLER_0_162_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31702_ clknet_leaf_43_clk _03160_ VGND VGND VPWR VPWR rvcpu.dp.pcreg.q\[20\] sky130_fd_sc_hd__dfxtp_1
X_19424_ datamem.data_ram\[38\]\[16\] _06719_ _06687_ datamem.data_ram\[36\]\[16\]
+ VGND VGND VPWR VPWR _06720_ sky130_fd_sc_hd__o22a_1
X_16636_ _14168_ net2841 _04551_ VGND VGND VPWR VPWR _04560_ sky130_fd_sc_hd__mux2_1
X_32682_ clknet_leaf_87_clk _04104_ VGND VGND VPWR VPWR datamem.data_ram\[18\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31633_ clknet_leaf_48_clk net1244 VGND VGND VPWR VPWR rvcpu.dp.plmw.lAuiPCW\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_19355_ _06650_ VGND VGND VPWR VPWR _06651_ sky130_fd_sc_hd__buf_6
XFILLER_0_186_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16567_ _14168_ net3057 _04514_ VGND VGND VPWR VPWR _04523_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18306_ _05670_ VGND VGND VPWR VPWR _05671_ sky130_fd_sc_hd__clkbuf_4
X_15518_ _13327_ _13771_ _14044_ VGND VGND VPWR VPWR _14045_ sky130_fd_sc_hd__and3_1
XFILLER_0_70_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_190_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31564_ clknet_leaf_63_clk datamem.rd_data_mem\[14\] VGND VGND VPWR VPWR rvcpu.dp.plmw.ReadDataW\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_19286_ _06581_ VGND VGND VPWR VPWR _06582_ sky130_fd_sc_hd__clkbuf_4
X_16498_ _04486_ VGND VGND VPWR VPWR _01794_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23915__472 clknet_1_0__leaf__10225_ VGND VGND VPWR VPWR net598 sky130_fd_sc_hd__inv_2
XFILLER_0_155_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_212_5573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18237_ _05410_ _05600_ _05419_ _05601_ VGND VGND VPWR VPWR _05602_ sky130_fd_sc_hd__nor4b_1
X_30515_ clknet_leaf_195_clk _02250_ VGND VGND VPWR VPWR datamem.data_ram\[56\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_212_5584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15449_ _13469_ _13961_ _13968_ _13979_ VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__o211ai_2
XTAP_TAPCELL_ROW_212_5595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31495_ clknet_leaf_44_clk rvcpu.dp.lAuiPCE\[21\] VGND VGND VPWR VPWR rvcpu.dp.plem.lAuiPCM\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18168_ rvcpu.dp.plde.RD1E\[24\] _05291_ _05532_ VGND VGND VPWR VPWR _05533_ sky130_fd_sc_hd__o21a_1
X_23614__233 clknet_1_0__leaf__10179_ VGND VGND VPWR VPWR net359 sky130_fd_sc_hd__inv_2
X_30446_ net784 _02181_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[29\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_23402__1017 clknet_1_0__leaf__10140_ VGND VGND VPWR VPWR net1143 sky130_fd_sc_hd__inv_2
Xmax_cap100 _10725_ VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__buf_4
XFILLER_0_111_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold403 datamem.data_ram\[57\]\[5\] VGND VGND VPWR VPWR net1553 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap111 _09300_ VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__clkbuf_2
Xhold414 datamem.data_ram\[19\]\[0\] VGND VGND VPWR VPWR net1564 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap122 rvcpu.dp.plem.ALUResultM\[2\] VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__buf_12
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17119_ _04816_ VGND VGND VPWR VPWR _01479_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_225_5901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold425 datamem.data_ram\[59\]\[6\] VGND VGND VPWR VPWR net1575 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold436 datamem.data_ram\[55\]\[2\] VGND VGND VPWR VPWR net1586 sky130_fd_sc_hd__dlygate4sd3_1
X_18099_ _05465_ _05466_ VGND VGND VPWR VPWR _05467_ sky130_fd_sc_hd__nor2_2
XFILLER_0_13_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30377_ net723 _02112_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[3\]\[28\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_146_4001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold447 rvcpu.dp.plfd.PCPlus4D\[2\] VGND VGND VPWR VPWR net1597 sky130_fd_sc_hd__dlygate4sd3_1
Xhold458 datamem.data_ram\[60\]\[2\] VGND VGND VPWR VPWR net1608 sky130_fd_sc_hd__dlygate4sd3_1
X_32116_ clknet_leaf_99_clk _03538_ VGND VGND VPWR VPWR datamem.data_ram\[0\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_20130_ datamem.data_ram\[8\]\[27\] _06696_ _06686_ datamem.data_ram\[12\]\[27\]
+ VGND VGND VPWR VPWR _07423_ sky130_fd_sc_hd__o22a_1
Xhold469 datamem.data_ram\[37\]\[7\] VGND VGND VPWR VPWR net1619 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_229_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_221_5809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_1267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32047_ clknet_leaf_132_clk _03469_ VGND VGND VPWR VPWR datamem.data_ram\[49\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_20061_ datamem.data_ram\[59\]\[26\] _06631_ VGND VGND VPWR VPWR _07355_ sky130_fd_sc_hd__or2_1
XFILLER_0_209_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26509__61 clknet_1_0__leaf__11602_ VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__inv_2
Xhold1103 datamem.data_ram\[11\]\[15\] VGND VGND VPWR VPWR net2253 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1114 rvcpu.dp.rf.reg_file_arr\[9\]\[2\] VGND VGND VPWR VPWR net2264 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1125 rvcpu.dp.rf.reg_file_arr\[7\]\[1\] VGND VGND VPWR VPWR net2275 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1136 datamem.data_ram\[11\]\[30\] VGND VGND VPWR VPWR net2286 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1147 rvcpu.dp.rf.reg_file_arr\[21\]\[16\] VGND VGND VPWR VPWR net2297 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1158 datamem.data_ram\[43\]\[22\] VGND VGND VPWR VPWR net2308 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1169 datamem.data_ram\[8\]\[20\] VGND VGND VPWR VPWR net2319 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20963_ datamem.data_ram\[57\]\[15\] _06653_ _08251_ _06598_ VGND VGND VPWR VPWR
+ _08252_ sky130_fd_sc_hd__o211a_1
XANTENNA_309 _14160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32949_ clknet_leaf_215_clk _04371_ VGND VGND VPWR VPWR datamem.data_ram\[6\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_219_5749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_176_4720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_92_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_92_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_176_4731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22702_ _09627_ _09845_ _09847_ _09795_ VGND VGND VPWR VPWR _09848_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_66_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26470_ _11576_ _11241_ _11540_ _06545_ _11591_ VGND VGND VPWR VPWR _11592_ sky130_fd_sc_hd__a221o_1
XFILLER_0_36_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20894_ datamem.data_ram\[2\]\[22\] datamem.data_ram\[3\]\[22\] _07837_ VGND VGND
+ VPWR VPWR _08184_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_172_4617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_4628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25421_ _10966_ VGND VGND VPWR VPWR _02744_ sky130_fd_sc_hd__clkbuf_1
X_22633_ rvcpu.dp.rf.reg_file_arr\[28\]\[17\] rvcpu.dp.rf.reg_file_arr\[30\]\[17\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[17\] rvcpu.dp.rf.reg_file_arr\[31\]\[17\] _09446_
+ _09402_ VGND VGND VPWR VPWR _09782_ sky130_fd_sc_hd__mux4_1
XFILLER_0_222_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25352_ _10408_ _10923_ VGND VGND VPWR VPWR _10925_ sky130_fd_sc_hd__and2_1
X_28140_ _12445_ net2091 _12528_ VGND VGND VPWR VPWR _12536_ sky130_fd_sc_hd__mux2_1
X_23243__891 clknet_1_0__leaf__10126_ VGND VGND VPWR VPWR net1017 sky130_fd_sc_hd__inv_2
X_22564_ rvcpu.dp.rf.reg_file_arr\[4\]\[13\] rvcpu.dp.rf.reg_file_arr\[5\]\[13\] rvcpu.dp.rf.reg_file_arr\[6\]\[13\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[13\] _09604_ _09716_ VGND VGND VPWR VPWR _09717_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_91_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24303_ _07125_ VGND VGND VPWR VPWR _10325_ sky130_fd_sc_hd__buf_6
XFILLER_0_17_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21515_ rvcpu.dp.rf.reg_file_arr\[0\]\[7\] rvcpu.dp.rf.reg_file_arr\[1\]\[7\] rvcpu.dp.rf.reg_file_arr\[2\]\[7\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[7\] _08550_ _08554_ VGND VGND VPWR VPWR _08770_ sky130_fd_sc_hd__mux4_1
X_28071_ _12499_ VGND VGND VPWR VPWR _03861_ sky130_fd_sc_hd__clkbuf_1
X_25283_ _10735_ net2902 _10878_ VGND VGND VPWR VPWR _10884_ sky130_fd_sc_hd__mux2_1
X_22495_ _09643_ _09647_ _09651_ _09491_ VGND VGND VPWR VPWR _01133_ sky130_fd_sc_hd__o31a_1
XFILLER_0_161_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27022_ _10325_ _11112_ _11898_ VGND VGND VPWR VPWR _11899_ sky130_fd_sc_hd__and3_1
X_24234_ _10268_ _09269_ _10269_ VGND VGND VPWR VPWR _10288_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_75_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21446_ rvcpu.dp.rf.reg_file_arr\[16\]\[4\] rvcpu.dp.rf.reg_file_arr\[17\]\[4\] rvcpu.dp.rf.reg_file_arr\[18\]\[4\]
+ rvcpu.dp.rf.reg_file_arr\[19\]\[4\] _08703_ _08629_ VGND VGND VPWR VPWR _08704_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_224_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_3635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_3646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23589__210 clknet_1_1__leaf__10177_ VGND VGND VPWR VPWR net336 sky130_fd_sc_hd__inv_2
XFILLER_0_82_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21377_ rvcpu.dp.rf.reg_file_arr\[28\]\[1\] rvcpu.dp.rf.reg_file_arr\[30\]\[1\] rvcpu.dp.rf.reg_file_arr\[29\]\[1\]
+ rvcpu.dp.rf.reg_file_arr\[31\]\[1\] _08635_ _08637_ VGND VGND VPWR VPWR _08638_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_9_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20328_ datamem.data_ram\[17\]\[4\] _06997_ _07617_ _07619_ VGND VGND VPWR VPWR _07620_
+ sky130_fd_sc_hd__a211o_1
X_28973_ _06587_ VGND VGND VPWR VPWR _12995_ sky130_fd_sc_hd__clkbuf_4
X_24096_ clknet_1_0__leaf__10244_ VGND VGND VPWR VPWR _10258_ sky130_fd_sc_hd__buf_1
Xhold970 datamem.data_ram\[45\]\[14\] VGND VGND VPWR VPWR net2120 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold981 rvcpu.dp.rf.reg_file_arr\[19\]\[14\] VGND VGND VPWR VPWR net2131 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_34_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27924_ _12128_ net4442 _12412_ VGND VGND VPWR VPWR _12414_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_34_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold992 rvcpu.dp.rf.reg_file_arr\[10\]\[3\] VGND VGND VPWR VPWR net2142 sky130_fd_sc_hd__dlygate4sd3_1
X_20259_ _06988_ _07529_ _07551_ VGND VGND VPWR VPWR _07552_ sky130_fd_sc_hd__and3_1
Xhold3050 datamem.data_ram\[29\]\[29\] VGND VGND VPWR VPWR net4200 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3061 rvcpu.dp.rf.reg_file_arr\[21\]\[9\] VGND VGND VPWR VPWR net4211 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold3072 datamem.data_ram\[58\]\[19\] VGND VGND VPWR VPWR net4222 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27855_ _12130_ net2921 _12373_ VGND VGND VPWR VPWR _12376_ sky130_fd_sc_hd__mux2_1
Xhold3083 rvcpu.dp.rf.reg_file_arr\[21\]\[20\] VGND VGND VPWR VPWR net4233 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3094 datamem.data_ram\[7\]\[16\] VGND VGND VPWR VPWR net4244 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2360 datamem.data_ram\[63\]\[16\] VGND VGND VPWR VPWR net3510 sky130_fd_sc_hd__dlygate4sd3_1
X_26806_ _11752_ VGND VGND VPWR VPWR _11767_ sky130_fd_sc_hd__buf_2
XFILLER_0_204_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14820_ _13314_ _13291_ VGND VGND VPWR VPWR _13373_ sky130_fd_sc_hd__nand2_1
Xhold2371 datamem.data_ram\[38\]\[8\] VGND VGND VPWR VPWR net3521 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2382 rvcpu.dp.rf.reg_file_arr\[27\]\[4\] VGND VGND VPWR VPWR net3532 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2393 datamem.data_ram\[46\]\[24\] VGND VGND VPWR VPWR net3543 sky130_fd_sc_hd__dlygate4sd3_1
X_27786_ _12095_ net2872 _12326_ VGND VGND VPWR VPWR _12334_ sky130_fd_sc_hd__mux2_1
X_24998_ _10448_ net3244 _10715_ VGND VGND VPWR VPWR _10720_ sky130_fd_sc_hd__mux2_1
Xhold1670 datamem.data_ram\[44\]\[22\] VGND VGND VPWR VPWR net2820 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_153_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29525_ clknet_leaf_261_clk _01260_ VGND VGND VPWR VPWR datamem.data_ram\[5\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_26737_ _11725_ _11603_ VGND VGND VPWR VPWR _11726_ sky130_fd_sc_hd__nor2_1
X_14751_ _13303_ VGND VGND VPWR VPWR _13304_ sky130_fd_sc_hd__clkbuf_4
Xhold1681 datamem.data_ram\[43\]\[18\] VGND VGND VPWR VPWR net2831 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1692 datamem.data_ram\[21\]\[12\] VGND VGND VPWR VPWR net2842 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_83_clk clknet_5_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_83_clk sky130_fd_sc_hd__clkbuf_8
X_17470_ _05002_ VGND VGND VPWR VPWR _01306_ sky130_fd_sc_hd__clkbuf_1
X_29456_ net818 _01191_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[30\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_26668_ _11683_ net1747 _11675_ _11685_ VGND VGND VPWR VPWR _03272_ sky130_fd_sc_hd__a31o_1
XFILLER_0_54_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14682_ _13246_ VGND VGND VPWR VPWR _03183_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16421_ net3122 _14451_ _14572_ VGND VGND VPWR VPWR _14577_ sky130_fd_sc_hd__mux2_1
X_28407_ _12680_ VGND VGND VPWR VPWR _04016_ sky130_fd_sc_hd__clkbuf_1
X_25619_ _10739_ net3130 net53 VGND VGND VPWR VPWR _11074_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_903 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29387_ clknet_leaf_174_clk _01122_ VGND VGND VPWR VPWR datamem.data_ram\[60\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_26599_ _11089_ _11640_ VGND VGND VPWR VPWR _11647_ sky130_fd_sc_hd__and2_1
XFILLER_0_132_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_184_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19140_ _06455_ _06456_ VGND VGND VPWR VPWR _06457_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_17_Left_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23025__727 clknet_1_0__leaf__10088_ VGND VGND VPWR VPWR net853 sky130_fd_sc_hd__inv_2
X_28338_ _12643_ VGND VGND VPWR VPWR _03984_ sky130_fd_sc_hd__clkbuf_1
X_16352_ _14540_ VGND VGND VPWR VPWR _01862_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0__10199_ _10199_ VGND VGND VPWR VPWR clknet_0__10199_ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_60_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_229_6001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15303_ _13419_ _13293_ _13482_ _13505_ VGND VGND VPWR VPWR _13841_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_229_6012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19071_ _06381_ _06388_ _06390_ _06386_ VGND VGND VPWR VPWR _06397_ sky130_fd_sc_hd__o31a_1
XFILLER_0_165_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_229_6023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28269_ _12361_ net3892 _12603_ VGND VGND VPWR VPWR _12606_ sky130_fd_sc_hd__mux2_1
X_16283_ net2881 _14449_ _14500_ VGND VGND VPWR VPWR _14504_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23105__784 clknet_1_1__leaf__10103_ VGND VGND VPWR VPWR net910 sky130_fd_sc_hd__inv_2
XFILLER_0_125_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18022_ _05391_ net115 _05173_ _05172_ rvcpu.dp.plde.ALUSrcE VGND VGND VPWR VPWR
+ _05392_ sky130_fd_sc_hd__a221o_1
X_30300_ net646 _02035_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[5\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_15234_ _13772_ _13774_ VGND VGND VPWR VPWR _13775_ sky130_fd_sc_hd__nand2_1
X_31280_ clknet_leaf_127_clk _02983_ VGND VGND VPWR VPWR datamem.data_ram\[24\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30231_ net585 _01966_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[7\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_15165_ _13509_ _13507_ _13565_ _13506_ VGND VGND VPWR VPWR _13709_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_2_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15096_ _13403_ _13523_ _13639_ _13640_ VGND VGND VPWR VPWR _13641_ sky130_fd_sc_hd__a211o_1
X_19973_ datamem.data_ram\[28\]\[18\] _06619_ _07265_ _07266_ VGND VGND VPWR VPWR
+ _07267_ sky130_fd_sc_hd__o211a_1
XFILLER_0_26_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30162_ net524 _01897_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[0\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_26_Left_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18924_ _05525_ _05537_ _05535_ VGND VGND VPWR VPWR _06263_ sky130_fd_sc_hd__a21o_1
XFILLER_0_66_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_226_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30093_ net455 _01828_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[11\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_600 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18855_ _05481_ _05728_ _06197_ _06198_ VGND VGND VPWR VPWR _06199_ sky130_fd_sc_hd__a211o_1
XFILLER_0_98_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17806_ _05198_ VGND VGND VPWR VPWR rvcpu.dp.SrcBFW_Mux.y\[31\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_59_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18786_ _05513_ _05616_ VGND VGND VPWR VPWR _06134_ sky130_fd_sc_hd__or2_1
X_15998_ net2136 _13254_ _14333_ VGND VGND VPWR VPWR _14337_ sky130_fd_sc_hd__mux2_1
XFILLER_0_222_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_167_Right_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32803_ clknet_leaf_165_clk _04225_ VGND VGND VPWR VPWR datamem.data_ram\[13\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_17737_ _13254_ net2525 _05140_ VGND VGND VPWR VPWR _05144_ sky130_fd_sc_hd__mux2_1
X_14949_ _13370_ _13373_ _13447_ VGND VGND VPWR VPWR _13498_ sky130_fd_sc_hd__or3_1
X_23186__856 clknet_1_0__leaf__10112_ VGND VGND VPWR VPWR net982 sky130_fd_sc_hd__inv_2
XFILLER_0_222_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30995_ clknet_leaf_99_clk _02730_ VGND VGND VPWR VPWR datamem.data_ram\[13\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_74_clk clknet_5_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_74_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32734_ clknet_leaf_83_clk _04156_ VGND VGND VPWR VPWR datamem.data_ram\[16\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_17668_ _05107_ VGND VGND VPWR VPWR _01205_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19407_ _06702_ VGND VGND VPWR VPWR _06703_ sky130_fd_sc_hd__buf_6
XFILLER_0_15_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_35_Left_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16619_ _04539_ VGND VGND VPWR VPWR _04551_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_214_5624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32665_ clknet_leaf_251_clk _04087_ VGND VGND VPWR VPWR datamem.data_ram\[19\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_214_5635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17599_ _13251_ net3496 _05068_ VGND VGND VPWR VPWR _05071_ sky130_fd_sc_hd__mux2_1
X_23458__107 clknet_1_0__leaf__10157_ VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__inv_2
XFILLER_0_174_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31616_ clknet_leaf_13_clk net1260 VGND VGND VPWR VPWR rvcpu.dp.plmw.RdW\[2\] sky130_fd_sc_hd__dfxtp_1
X_19338_ _06633_ VGND VGND VPWR VPWR _06634_ sky130_fd_sc_hd__buf_8
XFILLER_0_116_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32596_ clknet_leaf_252_clk _04018_ VGND VGND VPWR VPWR datamem.data_ram\[21\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19269_ rvcpu.c.ad.funct7b5 _06568_ rvcpu.c.ad.opb5 rvcpu.dp.plfd.InstrD\[12\] rvcpu.dp.plfd.InstrD\[13\]
+ VGND VGND VPWR VPWR _06569_ sky130_fd_sc_hd__a311o_1
X_31547_ clknet_leaf_14_clk net1154 VGND VGND VPWR VPWR rvcpu.dp.plem.RegWriteM sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21300_ rvcpu.dp.rf.reg_file_arr\[8\]\[0\] rvcpu.dp.rf.reg_file_arr\[10\]\[0\] rvcpu.dp.rf.reg_file_arr\[9\]\[0\]
+ rvcpu.dp.rf.reg_file_arr\[11\]\[0\] _08560_ _08561_ VGND VGND VPWR VPWR _08562_
+ sky130_fd_sc_hd__mux4_1
X_22280_ _09401_ VGND VGND VPWR VPWR _09445_ sky130_fd_sc_hd__buf_4
XFILLER_0_5_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31478_ clknet_leaf_65_clk rvcpu.dp.lAuiPCE\[4\] VGND VGND VPWR VPWR rvcpu.dp.plem.lAuiPCM\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold200 datamem.data_ram\[40\]\[5\] VGND VGND VPWR VPWR net1350 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21231_ datamem.data_ram\[52\]\[31\] datamem.data_ram\[52\]\[23\] datamem.data_ram\[53\]\[15\]
+ datamem.data_ram\[52\]\[15\] VGND VGND VPWR VPWR _08494_ sky130_fd_sc_hd__or4_1
Xhold211 datamem.data_ram\[42\]\[7\] VGND VGND VPWR VPWR net1361 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30429_ net767 _02164_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[29\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold222 datamem.data_ram\[17\]\[6\] VGND VGND VPWR VPWR net1372 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold233 datamem.data_ram\[6\]\[6\] VGND VGND VPWR VPWR net1383 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold244 datamem.data_ram\[13\]\[4\] VGND VGND VPWR VPWR net1394 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_44_Left_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold255 datamem.data_ram\[20\]\[3\] VGND VGND VPWR VPWR net1405 sky130_fd_sc_hd__dlygate4sd3_1
X_21162_ datamem.data_ram\[6\]\[23\] datamem.data_ram\[7\]\[23\] _07911_ VGND VGND
+ VPWR VPWR _08451_ sky130_fd_sc_hd__mux2_1
Xhold266 datamem.data_ram\[6\]\[3\] VGND VGND VPWR VPWR net1416 sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 datamem.data_ram\[56\]\[3\] VGND VGND VPWR VPWR net1427 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_165_4454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold288 datamem.data_ram\[29\]\[5\] VGND VGND VPWR VPWR net1438 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_165_4465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20113_ datamem.data_ram\[26\]\[10\] _06689_ _06645_ datamem.data_ram\[24\]\[10\]
+ VGND VGND VPWR VPWR _07407_ sky130_fd_sc_hd__o22a_1
Xhold299 datamem.data_ram\[12\]\[6\] VGND VGND VPWR VPWR net1449 sky130_fd_sc_hd__dlygate4sd3_1
X_25970_ net31 _11289_ VGND VGND VPWR VPWR _11308_ sky130_fd_sc_hd__or2_1
X_21093_ datamem.data_ram\[0\]\[7\] _06935_ _08381_ _07636_ _06598_ VGND VGND VPWR
+ VPWR _08382_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24024__555 clknet_1_1__leaf__10243_ VGND VGND VPWR VPWR net681 sky130_fd_sc_hd__inv_2
XFILLER_0_0_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24921_ _10465_ net3330 net91 VGND VGND VPWR VPWR _10679_ sky130_fd_sc_hd__mux2_1
X_20044_ datamem.data_ram\[2\]\[26\] _06691_ _07334_ _07337_ VGND VGND VPWR VPWR _07338_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_225_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27640_ _12255_ VGND VGND VPWR VPWR _03674_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24852_ _10385_ net3693 net93 VGND VGND VPWR VPWR _10642_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_3461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_134_Right_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_124_3472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27571_ _12087_ net3890 net82 VGND VGND VPWR VPWR _12219_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21995_ _07159_ VGND VGND VPWR VPWR _09225_ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_124_3483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24783_ _10468_ net3179 net94 VGND VGND VPWR VPWR _10604_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_65_clk clknet_5_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_65_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_106 _07023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_117 _07191_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29310_ clknet_leaf_290_clk _01045_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD1E\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_64_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_128 _07808_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26522_ _10061_ _11604_ _11605_ net1343 VGND VGND VPWR VPWR _03206_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_53_Left_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20946_ _07829_ _08235_ VGND VGND VPWR VPWR _08236_ sky130_fd_sc_hd__or2_1
XANTENNA_139 _07833_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29241_ _13140_ VGND VGND VPWR VPWR _04390_ sky130_fd_sc_hd__clkbuf_1
X_26453_ net1668 _11573_ _11580_ _11570_ VGND VGND VPWR VPWR _03162_ sky130_fd_sc_hd__o211a_1
XFILLER_0_193_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20877_ datamem.data_ram\[42\]\[14\] datamem.data_ram\[43\]\[14\] _07828_ VGND VGND
+ VPWR VPWR _08167_ sky130_fd_sc_hd__mux2_1
XFILLER_0_187_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25404_ _10416_ _10950_ VGND VGND VPWR VPWR _10957_ sky130_fd_sc_hd__and2_1
XFILLER_0_119_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_193_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29172_ _09225_ _10114_ _09230_ VGND VGND VPWR VPWR _13103_ sky130_fd_sc_hd__a21oi_2
X_22616_ _09390_ _09765_ VGND VGND VPWR VPWR _09766_ sky130_fd_sc_hd__or2_1
X_26384_ _13665_ _11268_ _11528_ _11530_ _10041_ VGND VGND VPWR VPWR _03143_ sky130_fd_sc_hd__o221a_1
XFILLER_0_153_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_193_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28123_ _12371_ net2932 _12519_ VGND VGND VPWR VPWR _12527_ sky130_fd_sc_hd__mux2_1
X_25335_ _10913_ VGND VGND VPWR VPWR _02711_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22547_ rvcpu.dp.rf.reg_file_arr\[12\]\[12\] rvcpu.dp.rf.reg_file_arr\[13\]\[12\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[12\] rvcpu.dp.rf.reg_file_arr\[15\]\[12\] _09552_
+ _09382_ VGND VGND VPWR VPWR _09701_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_98_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28054_ _12490_ VGND VGND VPWR VPWR _03853_ sky130_fd_sc_hd__clkbuf_1
X_25266_ _10538_ net1500 _10867_ _10874_ VGND VGND VPWR VPWR _02681_ sky130_fd_sc_hd__a31o_1
X_22478_ _09633_ _09634_ _09449_ VGND VGND VPWR VPWR _09635_ sky130_fd_sc_hd__mux2_2
XFILLER_0_49_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27005_ _11863_ net1723 _11885_ _11888_ VGND VGND VPWR VPWR _03406_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_94_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24217_ _10268_ _09229_ _10269_ VGND VGND VPWR VPWR _10279_ sky130_fd_sc_hd__a21oi_4
XPHY_EDGE_ROW_62_Left_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21429_ rvcpu.dp.rf.reg_file_arr\[4\]\[3\] rvcpu.dp.rf.reg_file_arr\[5\]\[3\] rvcpu.dp.rf.reg_file_arr\[6\]\[3\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[3\] _08687_ _08649_ VGND VGND VPWR VPWR _08688_ sky130_fd_sc_hd__mux4_1
X_25197_ _10836_ VGND VGND VPWR VPWR _02650_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_198_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24079_ _10251_ VGND VGND VPWR VPWR _02117_ sky130_fd_sc_hd__clkbuf_1
X_16970_ net2903 _14453_ _04731_ VGND VGND VPWR VPWR _04737_ sky130_fd_sc_hd__mux2_1
X_28956_ _12747_ net4261 _12978_ VGND VGND VPWR VPWR _12985_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27907_ _12145_ net3447 net47 VGND VGND VPWR VPWR _12405_ sky130_fd_sc_hd__mux2_1
X_15921_ net2405 _13241_ _14286_ VGND VGND VPWR VPWR _14296_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28887_ _12764_ net3889 _12941_ VGND VGND VPWR VPWR _12948_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18640_ _05996_ VGND VGND VPWR VPWR rvcpu.ALUResultE\[7\] sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_21_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27838_ _09317_ VGND VGND VPWR VPWR _12365_ sky130_fd_sc_hd__buf_2
X_15852_ _14235_ VGND VGND VPWR VPWR _14258_ sky130_fd_sc_hd__buf_4
XFILLER_0_217_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_216_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2190 datamem.data_ram\[36\]\[29\] VGND VGND VPWR VPWR net3340 sky130_fd_sc_hd__dlygate4sd3_1
X_14803_ rvcpu.dp.pcreg.q\[8\] _13313_ VGND VGND VPWR VPWR _13356_ sky130_fd_sc_hd__or2_1
XFILLER_0_203_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18571_ _05930_ VGND VGND VPWR VPWR rvcpu.ALUResultE\[4\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_118_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_803 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15783_ _14198_ VGND VGND VPWR VPWR _14221_ sky130_fd_sc_hd__buf_4
X_27769_ _12324_ VGND VGND VPWR VPWR _03734_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_101_Right_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_56_clk clknet_5_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_56_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29508_ net870 _01243_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[28\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_17522_ _13238_ net3536 _05021_ VGND VGND VPWR VPWR _05030_ sky130_fd_sc_hd__mux2_1
X_14734_ _13286_ VGND VGND VPWR VPWR _13287_ sky130_fd_sc_hd__buf_4
XFILLER_0_169_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30780_ clknet_leaf_194_clk _02515_ VGND VGND VPWR VPWR datamem.data_ram\[46\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_212_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17453_ _04993_ VGND VGND VPWR VPWR _01314_ sky130_fd_sc_hd__clkbuf_1
X_29439_ net801 _01174_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[30\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14665_ _13233_ VGND VGND VPWR VPWR _03187_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_211_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16404_ net2094 _14434_ _14561_ VGND VGND VPWR VPWR _14568_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32450_ clknet_leaf_286_clk _03872_ VGND VGND VPWR VPWR datamem.data_ram\[27\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17384_ _14166_ net3677 _04949_ VGND VGND VPWR VPWR _04957_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14596_ _13180_ VGND VGND VPWR VPWR _13181_ sky130_fd_sc_hd__buf_4
X_19123_ rvcpu.dp.plde.ImmExtE\[14\] rvcpu.dp.plde.PCE\[14\] VGND VGND VPWR VPWR _06442_
+ sky130_fd_sc_hd__or2_1
X_31401_ clknet_leaf_43_clk _03104_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCE\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_229_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16335_ _14531_ VGND VGND VPWR VPWR _01870_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32381_ clknet_leaf_166_clk _03803_ VGND VGND VPWR VPWR datamem.data_ram\[2\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_19054_ rvcpu.dp.plde.ImmExtE\[5\] rvcpu.dp.plde.PCE\[5\] VGND VGND VPWR VPWR _06382_
+ sky130_fd_sc_hd__and2_1
X_31332_ clknet_leaf_16_clk _03035_ VGND VGND VPWR VPWR rvcpu.dp.plde.RdE\[3\] sky130_fd_sc_hd__dfxtp_1
X_23986__521 clknet_1_1__leaf__10239_ VGND VGND VPWR VPWR net647 sky130_fd_sc_hd__inv_2
XFILLER_0_152_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16266_ net2238 _14432_ _14489_ VGND VGND VPWR VPWR _14495_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_207_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18005_ _05321_ rvcpu.dp.SrcBFW_Mux.y\[3\] _05369_ VGND VGND VPWR VPWR _05375_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_2_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15217_ _13343_ _13300_ VGND VGND VPWR VPWR _13758_ sky130_fd_sc_hd__nand2_2
XFILLER_0_164_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31263_ clknet_leaf_20_clk _02966_ VGND VGND VPWR VPWR rvcpu.dp.plfd.InstrD\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16197_ net2149 _14449_ _14443_ VGND VGND VPWR VPWR _14450_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__10111_ clknet_0__10111_ VGND VGND VPWR VPWR clknet_1_0__leaf__10111_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_23_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30214_ net568 _01949_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[7\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_15148_ _13297_ _13419_ VGND VGND VPWR VPWR _13692_ sky130_fd_sc_hd__nand2_1
XFILLER_0_140_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31194_ clknet_leaf_46_clk _02897_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCPlus4D\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_207_5461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30145_ net507 _01880_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[0\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_207_5472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15079_ _13450_ _13489_ _13484_ VGND VGND VPWR VPWR _13625_ sky130_fd_sc_hd__a21boi_1
X_19956_ datamem.data_ram\[62\]\[18\] _06628_ _06601_ _07249_ VGND VGND VPWR VPWR
+ _07250_ sky130_fd_sc_hd__o211a_1
X_18907_ _05703_ _06243_ _06246_ _06247_ VGND VGND VPWR VPWR _06248_ sky130_fd_sc_hd__a211o_1
X_30076_ net438 _01811_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[12\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_203_5358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19887_ _06688_ VGND VGND VPWR VPWR _07182_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_203_5369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_4340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_199_5262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_199_5273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18838_ _05497_ _06168_ _05571_ VGND VGND VPWR VPWR _06183_ sky130_fd_sc_hd__o21a_1
XFILLER_0_101_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_223_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_222_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18769_ _05335_ _06108_ _06118_ VGND VGND VPWR VPWR _06119_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_47_clk clknet_5_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_47_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_195_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20800_ datamem.data_ram\[51\]\[30\] _07849_ _08089_ _07851_ VGND VGND VPWR VPWR
+ _08090_ sky130_fd_sc_hd__a211o_1
XFILLER_0_222_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23309__950 clknet_1_1__leaf__10133_ VGND VGND VPWR VPWR net1076 sky130_fd_sc_hd__inv_2
X_21780_ _09021_ VGND VGND VPWR VPWR _01048_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_194_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30978_ clknet_leaf_91_clk _02713_ VGND VGND VPWR VPWR datamem.data_ram\[39\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20731_ _06615_ _08019_ _08020_ _07845_ VGND VGND VPWR VPWR _08021_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_158_4280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32717_ clknet_leaf_287_clk _04139_ VGND VGND VPWR VPWR datamem.data_ram\[17\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_158_4291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32648_ clknet_leaf_152_clk _04070_ VGND VGND VPWR VPWR datamem.data_ram\[1\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_20662_ datamem.data_ram\[61\]\[29\] _06661_ _06811_ datamem.data_ram\[56\]\[29\]
+ VGND VGND VPWR VPWR _07953_ sky130_fd_sc_hd__o22a_1
X_22401_ _09495_ _09561_ VGND VGND VPWR VPWR _09562_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_154_4188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_906 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22982__689 clknet_1_0__leaf__10083_ VGND VGND VPWR VPWR net815 sky130_fd_sc_hd__inv_2
XFILLER_0_163_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_4199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32579_ clknet_leaf_240_clk _04001_ VGND VGND VPWR VPWR datamem.data_ram\[21\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_20593_ datamem.data_ram\[22\]\[13\] _06628_ _07230_ datamem.data_ram\[20\]\[13\]
+ _07883_ VGND VGND VPWR VPWR _07884_ sky130_fd_sc_hd__o221a_1
XFILLER_0_2_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25120_ _10791_ VGND VGND VPWR VPWR _02618_ sky130_fd_sc_hd__clkbuf_1
X_22332_ rvcpu.dp.rf.reg_file_arr\[28\]\[2\] rvcpu.dp.rf.reg_file_arr\[30\]\[2\] rvcpu.dp.rf.reg_file_arr\[29\]\[2\]
+ rvcpu.dp.rf.reg_file_arr\[31\]\[2\] _09443_ _09453_ VGND VGND VPWR VPWR _09496_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_144_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_182_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_167_4505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25051_ _10751_ net3070 _10752_ VGND VGND VPWR VPWR _10753_ sky130_fd_sc_hd__mux2_1
X_22263_ _09399_ VGND VGND VPWR VPWR _09429_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21214_ _08487_ _07276_ _08490_ VGND VGND VPWR VPWR _04424_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_143_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22194_ _09369_ VGND VGND VPWR VPWR _01114_ sky130_fd_sc_hd__clkbuf_1
X_23355__992 clknet_1_0__leaf__10137_ VGND VGND VPWR VPWR net1118 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_203_Right_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28810_ _12907_ VGND VGND VPWR VPWR _04192_ sky130_fd_sc_hd__clkbuf_1
X_21145_ _07831_ _08431_ _08433_ VGND VGND VPWR VPWR _08434_ sky130_fd_sc_hd__o21a_1
X_29790_ net1136 _01525_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[20\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_126_3512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28741_ _12870_ VGND VGND VPWR VPWR _04160_ sky130_fd_sc_hd__clkbuf_1
X_25953_ net1823 _11290_ _11286_ _11298_ VGND VGND VPWR VPWR _02944_ sky130_fd_sc_hd__o211a_1
X_21076_ datamem.data_ram\[40\]\[7\] datamem.data_ram\[41\]\[7\] _07825_ VGND VGND
+ VPWR VPWR _08365_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_126_3523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20027_ _06715_ _07304_ _07309_ _07320_ VGND VGND VPWR VPWR _07321_ sky130_fd_sc_hd__a31o_1
X_24904_ _10385_ net4041 _10669_ VGND VGND VPWR VPWR _10670_ sky130_fd_sc_hd__mux2_1
X_28672_ _12754_ net2891 _12832_ VGND VGND VPWR VPWR _12834_ sky130_fd_sc_hd__mux2_1
X_25884_ rvcpu.dp.plfd.PCD\[1\] _11143_ VGND VGND VPWR VPWR _11259_ sky130_fd_sc_hd__or2_1
X_27623_ _12246_ VGND VGND VPWR VPWR _03666_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_225_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24835_ _10632_ VGND VGND VPWR VPWR _02492_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_38_clk clknet_5_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_38_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_87_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27554_ _12149_ net3988 net98 VGND VGND VPWR VPWR _12210_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24766_ _10472_ net3975 _10589_ VGND VGND VPWR VPWR _10593_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_200_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21978_ _08540_ _09208_ VGND VGND VPWR VPWR _09209_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23855__418 clknet_1_1__leaf__10219_ VGND VGND VPWR VPWR net544 sky130_fd_sc_hd__inv_2
X_20929_ datamem.data_ram\[36\]\[22\] datamem.data_ram\[37\]\[22\] _07827_ VGND VGND
+ VPWR VPWR _08219_ sky130_fd_sc_hd__mux2_1
X_27485_ _12132_ net2879 _12169_ VGND VGND VPWR VPWR _12173_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24697_ _10446_ net4178 _10552_ VGND VGND VPWR VPWR _10556_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0__10105_ _10105_ VGND VGND VPWR VPWR clknet_0__10105_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_96_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29224_ _11533_ net1417 _13122_ _13131_ VGND VGND VPWR VPWR _04382_ sky130_fd_sc_hd__a31o_1
X_26436_ _11545_ rvcpu.ALUResultE\[18\] VGND VGND VPWR VPWR _11568_ sky130_fd_sc_hd__and2_1
XFILLER_0_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23648_ _10190_ VGND VGND VPWR VPWR _01747_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29155_ _12601_ _10114_ _12977_ VGND VGND VPWR VPWR _13094_ sky130_fd_sc_hd__a21oi_4
X_26367_ _11089_ _11511_ VGND VGND VPWR VPWR _11518_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_70_Left_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16120_ _14402_ VGND VGND VPWR VPWR _01964_ sky130_fd_sc_hd__clkbuf_1
X_28106_ _12462_ net3056 _12510_ VGND VGND VPWR VPWR _12518_ sky130_fd_sc_hd__mux2_1
X_25318_ _10820_ net2591 _10899_ VGND VGND VPWR VPWR _10904_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29086_ _13057_ VGND VGND VPWR VPWR _04318_ sky130_fd_sc_hd__clkbuf_1
X_26298_ net1295 _11478_ VGND VGND VPWR VPWR _11482_ sky130_fd_sc_hd__and2_1
XFILLER_0_228_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_59_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28037_ _12445_ net2248 _12473_ VGND VGND VPWR VPWR _12481_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16051_ net2351 _13229_ _14360_ VGND VGND VPWR VPWR _14366_ sky130_fd_sc_hd__mux2_1
X_25249_ _10864_ VGND VGND VPWR VPWR _02674_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15002_ _13320_ _13510_ VGND VGND VPWR VPWR _13550_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19810_ _06680_ _07102_ _07104_ VGND VGND VPWR VPWR _07105_ sky130_fd_sc_hd__and3_1
XFILLER_0_103_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29988_ net358 _01723_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[14\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19741_ datamem.data_ram\[38\]\[25\] _06719_ _06687_ datamem.data_ram\[36\]\[25\]
+ VGND VGND VPWR VPWR _07036_ sky130_fd_sc_hd__o22a_1
X_16953_ net2251 _14436_ _04720_ VGND VGND VPWR VPWR _04728_ sky130_fd_sc_hd__mux2_1
XFILLER_0_202_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28939_ _12975_ VGND VGND VPWR VPWR _04253_ sky130_fd_sc_hd__clkbuf_1
X_15904_ _14287_ VGND VGND VPWR VPWR _02073_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_218_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19672_ datamem.data_ram\[51\]\[0\] _06966_ _06927_ datamem.data_ram\[55\]\[0\] _06967_
+ VGND VGND VPWR VPWR _06968_ sky130_fd_sc_hd__a221o_1
X_31950_ clknet_leaf_92_clk _03372_ VGND VGND VPWR VPWR datamem.data_ram\[32\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_23567__190 clknet_1_1__leaf__10175_ VGND VGND VPWR VPWR net316 sky130_fd_sc_hd__inv_2
XFILLER_0_217_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16884_ _04691_ VGND VGND VPWR VPWR _01597_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_194_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18623_ _05346_ _05405_ _05979_ VGND VGND VPWR VPWR _05980_ sky130_fd_sc_hd__o21a_1
X_30901_ clknet_leaf_222_clk _02636_ VGND VGND VPWR VPWR datamem.data_ram\[41\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15835_ _14249_ VGND VGND VPWR VPWR _02104_ sky130_fd_sc_hd__clkbuf_1
X_31881_ clknet_leaf_123_clk _03335_ VGND VGND VPWR VPWR datamem.data_ram\[57\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_29_clk clknet_5_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_29_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_204_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30832_ clknet_leaf_149_clk _02567_ VGND VGND VPWR VPWR datamem.data_ram\[44\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_18554_ _05365_ _05376_ _05662_ VGND VGND VPWR VPWR _05914_ sky130_fd_sc_hd__mux2_1
XFILLER_0_220_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15766_ _14212_ VGND VGND VPWR VPWR _02144_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17505_ _05009_ VGND VGND VPWR VPWR _05021_ sky130_fd_sc_hd__buf_4
X_14717_ net2264 _13272_ _13245_ VGND VGND VPWR VPWR _13273_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_190_5045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30763_ clknet_leaf_134_clk _02498_ VGND VGND VPWR VPWR datamem.data_ram\[47\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_18485_ _05441_ _05421_ _05769_ VGND VGND VPWR VPWR _05847_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_190_5056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15697_ _14168_ net2686 _14152_ VGND VGND VPWR VPWR _14169_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_190_5067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_470 _08954_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_699 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32502_ clknet_leaf_250_clk _03924_ VGND VGND VPWR VPWR datamem.data_ram\[25\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_481 _09317_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_492 _09750_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17436_ _04984_ VGND VGND VPWR VPWR _01322_ sky130_fd_sc_hd__clkbuf_1
X_14648_ net1981 _13220_ _13214_ VGND VGND VPWR VPWR _13221_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24053__581 clknet_1_0__leaf__10246_ VGND VGND VPWR VPWR net707 sky130_fd_sc_hd__inv_2
X_30694_ clknet_leaf_155_clk _02429_ VGND VGND VPWR VPWR datamem.data_ram\[4\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_17 _06612_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32433_ clknet_leaf_231_clk _03855_ VGND VGND VPWR VPWR datamem.data_ram\[27\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_28 _06634_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_39 _06677_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17367_ _14149_ net3553 _04938_ VGND VGND VPWR VPWR _04948_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19106_ rvcpu.dp.plde.ImmExtE\[12\] rvcpu.dp.plde.PCE\[12\] VGND VGND VPWR VPWR _06427_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_67_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16318_ net1959 _14484_ _14488_ VGND VGND VPWR VPWR _14522_ sky130_fd_sc_hd__mux2_1
X_32364_ clknet_leaf_94_clk _03786_ VGND VGND VPWR VPWR datamem.data_ram\[2\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_17298_ _04911_ VGND VGND VPWR VPWR _01395_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_209_5501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19037_ rvcpu.dp.plde.ImmExtE\[3\] rvcpu.dp.plde.PCE\[3\] VGND VGND VPWR VPWR _06367_
+ sky130_fd_sc_hd__nand2_1
X_31315_ clknet_leaf_29_clk _03018_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCPlus4E\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_209_5512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16249_ net3077 _14484_ _14421_ VGND VGND VPWR VPWR _14485_ sky130_fd_sc_hd__mux2_1
XFILLER_0_179_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32295_ clknet_leaf_193_clk _03717_ VGND VGND VPWR VPWR datamem.data_ram\[32\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_209_5523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_600 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31246_ clknet_leaf_21_clk _02949_ VGND VGND VPWR VPWR rvcpu.dp.plfd.InstrD\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_205_5409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31177_ clknet_leaf_235_clk _02880_ VGND VGND VPWR VPWR datamem.data_ram\[5\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2904 datamem.data_ram\[46\]\[19\] VGND VGND VPWR VPWR net4054 sky130_fd_sc_hd__dlygate4sd3_1
X_30128_ net490 _01863_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[10\]\[19\] sky130_fd_sc_hd__dfxtp_1
Xhold2915 rvcpu.dp.rf.reg_file_arr\[21\]\[13\] VGND VGND VPWR VPWR net4065 sky130_fd_sc_hd__dlygate4sd3_1
X_19939_ datamem.data_ram\[38\]\[18\] _06629_ _07231_ _07232_ VGND VGND VPWR VPWR
+ _07233_ sky130_fd_sc_hd__o211a_1
Xhold2926 datamem.data_ram\[6\]\[26\] VGND VGND VPWR VPWR net4076 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2937 datamem.data_ram\[21\]\[16\] VGND VGND VPWR VPWR net4087 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2948 datamem.data_ram\[10\]\[25\] VGND VGND VPWR VPWR net4098 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2959 rvcpu.dp.rf.reg_file_arr\[28\]\[2\] VGND VGND VPWR VPWR net4109 sky130_fd_sc_hd__dlygate4sd3_1
X_24095__604 clknet_1_0__leaf__10248_ VGND VGND VPWR VPWR net730 sky130_fd_sc_hd__inv_2
X_22950_ _10076_ _10053_ VGND VGND VPWR VPWR _10077_ sky130_fd_sc_hd__and2_1
XFILLER_0_138_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30059_ net421 _01794_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[12\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21901_ rvcpu.dp.rf.reg_file_arr\[4\]\[27\] rvcpu.dp.rf.reg_file_arr\[5\]\[27\] rvcpu.dp.rf.reg_file_arr\[6\]\[27\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[27\] _08628_ _08856_ VGND VGND VPWR VPWR _09136_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_179_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22881_ _09429_ _10014_ _10016_ VGND VGND VPWR VPWR _10017_ sky130_fd_sc_hd__a21o_1
XFILLER_0_222_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_218_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24620_ _10442_ net3746 _10511_ VGND VGND VPWR VPWR _10513_ sky130_fd_sc_hd__mux2_1
X_21832_ rvcpu.dp.rf.reg_file_arr\[0\]\[23\] rvcpu.dp.rf.reg_file_arr\[1\]\[23\] rvcpu.dp.rf.reg_file_arr\[2\]\[23\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[23\] _08550_ _08554_ VGND VGND VPWR VPWR _09071_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_211_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_179_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_214_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_156_4228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_4239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24551_ _10473_ VGND VGND VPWR VPWR _02367_ sky130_fd_sc_hd__clkbuf_1
X_21763_ _08514_ _09004_ VGND VGND VPWR VPWR _09005_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26494__47 clknet_1_1__leaf__11601_ VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__inv_2
X_20714_ datamem.data_ram\[18\]\[5\] _06932_ _06958_ datamem.data_ram\[17\]\[5\] VGND
+ VGND VPWR VPWR _08005_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27270_ _12046_ VGND VGND VPWR VPWR _03513_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_191_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24482_ _10431_ VGND VGND VPWR VPWR _02340_ sky130_fd_sc_hd__clkbuf_1
X_21694_ rvcpu.dp.rf.reg_file_arr\[28\]\[16\] rvcpu.dp.rf.reg_file_arr\[30\]\[16\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[16\] rvcpu.dp.rf.reg_file_arr\[31\]\[16\] _08568_
+ _08683_ VGND VGND VPWR VPWR _08940_ sky130_fd_sc_hd__mux4_1
XFILLER_0_110_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26221_ _11448_ VGND VGND VPWR VPWR _03062_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_3360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20645_ datamem.data_ram\[31\]\[29\] _06671_ _06806_ datamem.data_ram\[28\]\[29\]
+ VGND VGND VPWR VPWR _07936_ sky130_fd_sc_hd__o22a_1
X_23433_ clknet_1_0__leaf__10152_ VGND VGND VPWR VPWR _10155_ sky130_fd_sc_hd__buf_1
XFILLER_0_11_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_866 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_1248 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26152_ _11412_ VGND VGND VPWR VPWR _03028_ sky130_fd_sc_hd__clkbuf_1
X_20576_ _07866_ VGND VGND VPWR VPWR _07867_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_115_3246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_3257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25103_ _10073_ _10779_ _10781_ net1592 VGND VGND VPWR VPWR _02610_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_410 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22315_ rvcpu.dp.rf.reg_file_arr\[12\]\[1\] rvcpu.dp.rf.reg_file_arr\[13\]\[1\] rvcpu.dp.rf.reg_file_arr\[14\]\[1\]
+ rvcpu.dp.rf.reg_file_arr\[15\]\[1\] _09478_ _09479_ VGND VGND VPWR VPWR _09480_
+ sky130_fd_sc_hd__mux4_1
X_26083_ rvcpu.c.ad.opb5 VGND VGND VPWR VPWR _11374_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_186_4958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_186_4969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29911_ net281 _01646_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[16\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_25034_ _10743_ VGND VGND VPWR VPWR _02580_ sky130_fd_sc_hd__clkbuf_1
X_22246_ _09411_ VGND VGND VPWR VPWR _09412_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_132_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_225_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29842_ net220 _01577_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[18\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_22177_ _09330_ net2212 _09352_ VGND VGND VPWR VPWR _09360_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21128_ datamem.data_ram\[38\]\[23\] datamem.data_ram\[39\]\[23\] _07912_ VGND VGND
+ VPWR VPWR _08417_ sky130_fd_sc_hd__mux2_1
X_29773_ net1119 _01508_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[20\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_26985_ _10754_ net3083 _11875_ VGND VGND VPWR VPWR _11877_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28724_ _12861_ VGND VGND VPWR VPWR _04152_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_145_3965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25936_ _11288_ VGND VGND VPWR VPWR _11289_ sky130_fd_sc_hd__clkbuf_2
X_21059_ datamem.data_ram\[46\]\[31\] datamem.data_ram\[47\]\[31\] _07825_ VGND VGND
+ VPWR VPWR _08348_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_145_3976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28655_ _12690_ net3612 _12823_ VGND VGND VPWR VPWR _12825_ sky130_fd_sc_hd__mux2_1
X_25867_ _11206_ _11207_ _11245_ VGND VGND VPWR VPWR _11246_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_775 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15620_ _14118_ VGND VGND VPWR VPWR _02196_ sky130_fd_sc_hd__clkbuf_1
X_27606_ _12237_ VGND VGND VPWR VPWR _03658_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24818_ _10388_ net3580 _10621_ VGND VGND VPWR VPWR _10623_ sky130_fd_sc_hd__mux2_1
XFILLER_0_214_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28586_ _12737_ net4142 _12786_ VGND VGND VPWR VPWR _12788_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25798_ net1728 _11181_ _11177_ _11190_ VGND VGND VPWR VPWR _02897_ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15551_ _13760_ _13420_ _14074_ _13458_ VGND VGND VPWR VPWR _14075_ sky130_fd_sc_hd__a31o_1
X_27537_ _12132_ net2322 _12197_ VGND VGND VPWR VPWR _12201_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24749_ _10392_ net3450 _10580_ VGND VGND VPWR VPWR _10584_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_104_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_210_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18270_ _05632_ _05528_ _05634_ VGND VGND VPWR VPWR _05635_ sky130_fd_sc_hd__o21a_1
XFILLER_0_96_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15482_ _13297_ _13322_ _13586_ VGND VGND VPWR VPWR _14011_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_13_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27468_ _12163_ VGND VGND VPWR VPWR _03594_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29207_ _13121_ VGND VGND VPWR VPWR _13122_ sky130_fd_sc_hd__buf_2
XFILLER_0_37_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17221_ _04870_ VGND VGND VPWR VPWR _01431_ sky130_fd_sc_hd__clkbuf_1
X_26419_ _06432_ _11539_ _11529_ _11180_ _11556_ VGND VGND VPWR VPWR _11557_ sky130_fd_sc_hd__a221o_1
XFILLER_0_140_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27399_ _12119_ VGND VGND VPWR VPWR _03569_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_182_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17152_ _14139_ net4410 _04829_ VGND VGND VPWR VPWR _04834_ sky130_fd_sc_hd__mux2_1
X_29138_ _10979_ _10092_ _12977_ VGND VGND VPWR VPWR _13085_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_108_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16103_ _14393_ VGND VGND VPWR VPWR _01972_ sky130_fd_sc_hd__clkbuf_1
X_29069_ _13048_ VGND VGND VPWR VPWR _04310_ sky130_fd_sc_hd__clkbuf_1
X_17083_ _04797_ VGND VGND VPWR VPWR _01496_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31100_ clknet_leaf_280_clk _02835_ VGND VGND VPWR VPWR datamem.data_ram\[9\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16034_ net2547 _13204_ _14349_ VGND VGND VPWR VPWR _14357_ sky130_fd_sc_hd__mux2_1
X_32080_ clknet_leaf_93_clk _03502_ VGND VGND VPWR VPWR datamem.data_ram\[33\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_1034 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31031_ clknet_leaf_54_clk _02766_ VGND VGND VPWR VPWR datamem.data_ram\[12\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17985_ _05349_ _05353_ VGND VGND VPWR VPWR _05355_ sky130_fd_sc_hd__nor2_1
XFILLER_0_165_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_200_5306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16936_ _04718_ VGND VGND VPWR VPWR _01572_ sky130_fd_sc_hd__clkbuf_1
X_19724_ _06865_ VGND VGND VPWR VPWR _07019_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_196_5210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23723__315 clknet_1_0__leaf__10198_ VGND VGND VPWR VPWR net441 sky130_fd_sc_hd__inv_2
X_32982_ clknet_leaf_269_clk _04404_ VGND VGND VPWR VPWR datamem.data_ram\[63\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_19655_ _06950_ VGND VGND VPWR VPWR _06951_ sky130_fd_sc_hd__buf_4
X_31933_ clknet_leaf_113_clk _03355_ VGND VGND VPWR VPWR datamem.data_ram\[60\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_16867_ net2564 _14486_ _04647_ VGND VGND VPWR VPWR _04682_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_192_5107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18606_ _05750_ _05963_ VGND VGND VPWR VPWR _05964_ sky130_fd_sc_hd__nor2_1
X_15818_ _14240_ VGND VGND VPWR VPWR _02112_ sky130_fd_sc_hd__clkbuf_1
X_31864_ clknet_leaf_111_clk _03318_ VGND VGND VPWR VPWR datamem.data_ram\[63\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_19586_ datamem.data_ram\[42\]\[8\] _06689_ _06644_ datamem.data_ram\[40\]\[8\] VGND
+ VGND VPWR VPWR _06882_ sky130_fd_sc_hd__o22a_1
X_16798_ _04645_ VGND VGND VPWR VPWR _01645_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_204_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_9_Left_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18537_ _05704_ _05897_ VGND VGND VPWR VPWR _05898_ sky130_fd_sc_hd__nor2_1
X_30815_ clknet_leaf_264_clk _02550_ VGND VGND VPWR VPWR datamem.data_ram\[45\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_15749_ _14203_ VGND VGND VPWR VPWR _02152_ sky130_fd_sc_hd__clkbuf_1
X_31795_ clknet_leaf_235_clk _03249_ VGND VGND VPWR VPWR datamem.data_ram\[2\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30746_ clknet_leaf_136_clk _02481_ VGND VGND VPWR VPWR datamem.data_ram\[48\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_18468_ _05327_ _05446_ _05412_ _05441_ _05683_ _05688_ VGND VGND VPWR VPWR _05831_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_8_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_151_4114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17419_ _14133_ net4034 _04974_ VGND VGND VPWR VPWR _04976_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_151_4125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30677_ clknet_leaf_96_clk _02412_ VGND VGND VPWR VPWR datamem.data_ram\[4\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_18399_ _05705_ _05762_ VGND VGND VPWR VPWR _05763_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20430_ datamem.data_ram\[14\]\[12\] _07085_ _06618_ datamem.data_ram\[12\]\[12\]
+ _07721_ VGND VGND VPWR VPWR _07722_ sky130_fd_sc_hd__o221a_1
X_32416_ clknet_leaf_182_clk _03838_ VGND VGND VPWR VPWR datamem.data_ram\[28\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32347_ clknet_leaf_80_clk _03769_ VGND VGND VPWR VPWR datamem.data_ram\[30\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload220 clknet_leaf_176_clk VGND VGND VPWR VPWR clkload220/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20361_ datamem.data_ram\[7\]\[28\] _06725_ _07243_ datamem.data_ram\[1\]\[28\] VGND
+ VGND VPWR VPWR _07653_ sky130_fd_sc_hd__o22a_1
Xclkload231 clknet_leaf_110_clk VGND VGND VPWR VPWR clkload231/Y sky130_fd_sc_hd__clkinv_1
Xclkbuf_leaf_9_clk clknet_5_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_8
Xclkload242 clknet_leaf_124_clk VGND VGND VPWR VPWR clkload242/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_0_3_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22100_ _09311_ VGND VGND VPWR VPWR _01078_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_5_15__f_clk clknet_2_1_0_clk VGND VGND VPWR VPWR clknet_5_15__leaf_clk sky130_fd_sc_hd__clkbuf_16
Xclkload253 clknet_leaf_191_clk VGND VGND VPWR VPWR clkload253/Y sky130_fd_sc_hd__clkinv_4
Xclkload264 clknet_leaf_197_clk VGND VGND VPWR VPWR clkload264/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_228_5965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload275 clknet_leaf_130_clk VGND VGND VPWR VPWR clkload275/Y sky130_fd_sc_hd__clkinv_1
X_32278_ clknet_leaf_90_clk _03700_ VGND VGND VPWR VPWR datamem.data_ram\[33\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_20292_ datamem.data_ram\[14\]\[19\] _06764_ _06700_ datamem.data_ram\[9\]\[19\]
+ VGND VGND VPWR VPWR _07585_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_110_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_228_5976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload286 clknet_1_1__leaf__10243_ VGND VGND VPWR VPWR clkload286/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_110_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_4065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload297 clknet_1_1__leaf__10219_ VGND VGND VPWR VPWR clkload297/Y sky130_fd_sc_hd__clkinvlp_4
X_22031_ rvcpu.dp.plem.WriteDataM\[6\] _09215_ _09219_ _09254_ VGND VGND VPWR VPWR
+ _09255_ sky130_fd_sc_hd__a31o_4
XTAP_TAPCELL_ROW_149_4076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31229_ clknet_leaf_43_clk _02932_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCD\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_220_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_181_4833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24103__611 clknet_1_0__leaf__10258_ VGND VGND VPWR VPWR net737 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_181_4844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2701 rvcpu.dp.rf.reg_file_arr\[30\]\[19\] VGND VGND VPWR VPWR net3851 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2712 datamem.data_ram\[39\]\[14\] VGND VGND VPWR VPWR net3862 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2723 rvcpu.dp.rf.reg_file_arr\[4\]\[24\] VGND VGND VPWR VPWR net3873 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2734 rvcpu.dp.rf.reg_file_arr\[29\]\[21\] VGND VGND VPWR VPWR net3884 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2745 rvcpu.dp.rf.reg_file_arr\[8\]\[17\] VGND VGND VPWR VPWR net3895 sky130_fd_sc_hd__dlygate4sd3_1
X_26770_ _11689_ _11738_ VGND VGND VPWR VPWR _11745_ sky130_fd_sc_hd__and2_1
Xhold2756 rvcpu.dp.rf.reg_file_arr\[30\]\[20\] VGND VGND VPWR VPWR net3906 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_199_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2767 rvcpu.dp.rf.reg_file_arr\[12\]\[28\] VGND VGND VPWR VPWR net3917 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2778 rvcpu.dp.rf.reg_file_arr\[19\]\[8\] VGND VGND VPWR VPWR net3928 sky130_fd_sc_hd__dlygate4sd3_1
X_23663__262 clknet_1_0__leaf__10191_ VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__inv_2
Xhold2789 datamem.data_ram\[56\]\[16\] VGND VGND VPWR VPWR net3939 sky130_fd_sc_hd__dlygate4sd3_1
X_25721_ _11134_ VGND VGND VPWR VPWR _02876_ sky130_fd_sc_hd__clkbuf_1
X_22933_ _10063_ VGND VGND VPWR VPWR _10064_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_84_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28440_ _12700_ net3993 _12688_ VGND VGND VPWR VPWR _12701_ sky130_fd_sc_hd__mux2_1
X_25652_ _10061_ _11094_ _11095_ net1320 VGND VGND VPWR VPWR _02846_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_140_3851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_210_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_616 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_140_3862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22864_ rvcpu.dp.rf.reg_file_arr\[12\]\[29\] rvcpu.dp.rf.reg_file_arr\[13\]\[29\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[29\] rvcpu.dp.rf.reg_file_arr\[15\]\[29\] _09462_
+ _09465_ VGND VGND VPWR VPWR _10001_ sky130_fd_sc_hd__mux4_1
XFILLER_0_74_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_179_4784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_179_4795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24603_ _10468_ net3073 _10502_ VGND VGND VPWR VPWR _10504_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21815_ _08817_ _09052_ _09054_ _08700_ VGND VGND VPWR VPWR _09055_ sky130_fd_sc_hd__a211o_1
X_28371_ _12359_ net3497 _12659_ VGND VGND VPWR VPWR _12661_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25583_ _11052_ VGND VGND VPWR VPWR _11053_ sky130_fd_sc_hd__buf_2
XFILLER_0_149_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22795_ _09927_ _09931_ _09935_ _09491_ VGND VGND VPWR VPWR _01149_ sky130_fd_sc_hd__o31a_1
X_27322_ _10780_ _12076_ VGND VGND VPWR VPWR _12077_ sky130_fd_sc_hd__nor2_2
XFILLER_0_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire94 _10602_ VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__buf_4
X_24534_ _10462_ VGND VGND VPWR VPWR _02361_ sky130_fd_sc_hd__clkbuf_1
X_21746_ _08798_ _08988_ VGND VGND VPWR VPWR _08989_ sky130_fd_sc_hd__or2_1
XFILLER_0_93_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27253_ _12036_ net1534 _12030_ _12040_ VGND VGND VPWR VPWR _03502_ sky130_fd_sc_hd__a31o_1
XFILLER_0_148_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24465_ _10422_ VGND VGND VPWR VPWR _02332_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21677_ _08798_ _08921_ _08923_ _08806_ VGND VGND VPWR VPWR _08924_ sky130_fd_sc_hd__o211a_1
XFILLER_0_19_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_184_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26204_ _11440_ VGND VGND VPWR VPWR _03053_ sky130_fd_sc_hd__buf_1
XFILLER_0_164_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27184_ _11972_ _11996_ VGND VGND VPWR VPWR _12000_ sky130_fd_sc_hd__and2_1
XFILLER_0_149_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20628_ _07898_ _07904_ _07918_ VGND VGND VPWR VPWR _07919_ sky130_fd_sc_hd__and3_1
XFILLER_0_190_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24396_ _10377_ VGND VGND VPWR VPWR _02308_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_78_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26135_ _11403_ VGND VGND VPWR VPWR _03020_ sky130_fd_sc_hd__clkbuf_1
X_20559_ _07823_ datamem.data_ram\[10\]\[21\] datamem.data_ram\[11\]\[21\] _07849_
+ VGND VGND VPWR VPWR _07850_ sky130_fd_sc_hd__a22o_1
X_23347_ clknet_1_0__leaf__10130_ VGND VGND VPWR VPWR _10137_ sky130_fd_sc_hd__buf_1
XFILLER_0_85_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26066_ rvcpu.dp.plfd.InstrD\[6\] _11361_ _11362_ VGND VGND VPWR VPWR _11363_ sky130_fd_sc_hd__and3b_1
X_25017_ _10731_ net4198 net100 VGND VGND VPWR VPWR _10732_ sky130_fd_sc_hd__mux2_1
X_22229_ _09394_ VGND VGND VPWR VPWR _09395_ sky130_fd_sc_hd__buf_4
XFILLER_0_30_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29825_ net203 _01560_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[1\]\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_37_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17770_ rvcpu.dp.plem.RdM\[3\] rvcpu.dp.plde.Rs2E\[3\] VGND VGND VPWR VPWR _05168_
+ sky130_fd_sc_hd__and2_1
X_14982_ _13423_ _13525_ _13527_ _13529_ VGND VGND VPWR VPWR _13530_ sky130_fd_sc_hd__o211a_1
X_26968_ _11825_ _11866_ VGND VGND VPWR VPWR _11868_ sky130_fd_sc_hd__and2_1
X_29756_ net1102 _01491_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[21\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_16721_ _14185_ net2965 _04598_ VGND VGND VPWR VPWR _04605_ sky130_fd_sc_hd__mux2_1
X_25919_ _11142_ VGND VGND VPWR VPWR _11279_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_191_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28707_ _12852_ VGND VGND VPWR VPWR _04144_ sky130_fd_sc_hd__clkbuf_1
X_29687_ net1033 _01422_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[23\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_26899_ _11822_ _11823_ VGND VGND VPWR VPWR _11824_ sky130_fd_sc_hd__and2_1
XFILLER_0_156_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19440_ datamem.data_ram\[32\]\[16\] _06698_ _06720_ _06735_ VGND VGND VPWR VPWR
+ _06736_ sky130_fd_sc_hd__o211a_1
X_16652_ _04568_ VGND VGND VPWR VPWR _01714_ sky130_fd_sc_hd__clkbuf_1
X_28638_ _12737_ net1979 net71 VGND VGND VPWR VPWR _12816_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15603_ _14109_ VGND VGND VPWR VPWR _02204_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_187_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19371_ _06666_ _06623_ VGND VGND VPWR VPWR _06667_ sky130_fd_sc_hd__nand2_8
X_28569_ _12754_ net2977 _12777_ VGND VGND VPWR VPWR _12779_ sky130_fd_sc_hd__mux2_1
X_16583_ _04531_ VGND VGND VPWR VPWR _01754_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_215_73 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18322_ _05373_ _05663_ _05686_ VGND VGND VPWR VPWR _05687_ sky130_fd_sc_hd__o21a_1
X_30600_ clknet_leaf_219_clk _02335_ VGND VGND VPWR VPWR datamem.data_ram\[53\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_215_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15534_ _13564_ _14059_ _13442_ VGND VGND VPWR VPWR _14060_ sky130_fd_sc_hd__a21o_1
XFILLER_0_174_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31580_ clknet_leaf_75_clk datamem.rd_data_mem\[30\] VGND VGND VPWR VPWR rvcpu.dp.plmw.ReadDataW\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18253_ _05574_ _05485_ _05616_ _05617_ VGND VGND VPWR VPWR _05618_ sky130_fd_sc_hd__o22a_1
X_30531_ clknet_leaf_180_clk _02266_ VGND VGND VPWR VPWR datamem.data_ram\[56\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_15465_ _13893_ _13994_ VGND VGND VPWR VPWR _13995_ sky130_fd_sc_hd__nand2_1
XFILLER_0_166_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_568 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17204_ _14191_ net2187 _04851_ VGND VGND VPWR VPWR _04861_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18184_ _05547_ _05548_ VGND VGND VPWR VPWR _05549_ sky130_fd_sc_hd__nor2_2
X_30462_ net140 _02197_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[19\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_15396_ _13434_ _13574_ VGND VGND VPWR VPWR _13929_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32201_ clknet_leaf_169_clk _03623_ VGND VGND VPWR VPWR datamem.data_ram\[36\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17135_ _04824_ VGND VGND VPWR VPWR _01471_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30393_ net731 _02128_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[31\]\[4\] sky130_fd_sc_hd__dfxtp_1
Xhold607 datamem.data_ram\[9\]\[5\] VGND VGND VPWR VPWR net1757 sky130_fd_sc_hd__dlygate4sd3_1
Xhold618 datamem.data_ram\[25\]\[2\] VGND VGND VPWR VPWR net1768 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32132_ clknet_leaf_233_clk _03554_ VGND VGND VPWR VPWR datamem.data_ram\[10\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold629 datamem.data_ram\[62\]\[3\] VGND VGND VPWR VPWR net1779 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17066_ net1961 _14480_ _04779_ VGND VGND VPWR VPWR _04788_ sky130_fd_sc_hd__mux2_1
X_23532__159 clknet_1_0__leaf__10171_ VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__inv_2
XFILLER_0_64_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16017_ rvcpu.dp.plmw.RegWriteW _14346_ rvcpu.dp.plmw.RdW\[1\] VGND VGND VPWR VPWR
+ _14347_ sky130_fd_sc_hd__nand3_4
X_32063_ clknet_leaf_133_clk _03485_ VGND VGND VPWR VPWR datamem.data_ram\[48\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31014_ clknet_leaf_155_clk _02749_ VGND VGND VPWR VPWR datamem.data_ram\[42\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_223_5840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_223_5851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2008 datamem.data_ram\[7\]\[8\] VGND VGND VPWR VPWR net3158 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2019 datamem.data_ram\[10\]\[30\] VGND VGND VPWR VPWR net3169 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_225_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_260_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_260_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold1307 rvcpu.dp.rf.reg_file_arr\[11\]\[9\] VGND VGND VPWR VPWR net2457 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1318 rvcpu.dp.rf.reg_file_arr\[29\]\[7\] VGND VGND VPWR VPWR net2468 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17968_ _05293_ VGND VGND VPWR VPWR _05339_ sky130_fd_sc_hd__buf_2
Xhold1329 rvcpu.dp.plfd.InstrD\[24\] VGND VGND VPWR VPWR net2479 sky130_fd_sc_hd__dlygate4sd3_1
X_19707_ datamem.data_ram\[1\]\[0\] _06997_ _06999_ _07002_ VGND VGND VPWR VPWR _07003_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_139_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16919_ net1874 _14470_ _04706_ VGND VGND VPWR VPWR _04710_ sky130_fd_sc_hd__mux2_1
XFILLER_0_212_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32965_ clknet_leaf_218_clk _04387_ VGND VGND VPWR VPWR datamem.data_ram\[63\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_17899_ _05268_ VGND VGND VPWR VPWR _05272_ sky130_fd_sc_hd__buf_2
XFILLER_0_205_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31916_ _04428_ net120 VGND VGND VPWR VPWR datamem.rd_data_mem\[21\] sky130_fd_sc_hd__dlxtn_1
X_19638_ _06606_ _06614_ VGND VGND VPWR VPWR _06934_ sky130_fd_sc_hd__nand2_8
XFILLER_0_36_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_215_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32896_ clknet_leaf_165_clk _04318_ VGND VGND VPWR VPWR datamem.data_ram\[10\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31847_ clknet_leaf_124_clk _03301_ VGND VGND VPWR VPWR datamem.data_ram\[61\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19569_ _06724_ VGND VGND VPWR VPWR _06865_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_177_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21600_ rvcpu.dp.rf.reg_file_arr\[24\]\[11\] rvcpu.dp.rf.reg_file_arr\[25\]\[11\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[11\] rvcpu.dp.rf.reg_file_arr\[27\]\[11\] _08548_
+ _08526_ VGND VGND VPWR VPWR _08851_ sky130_fd_sc_hd__mux4_1
XFILLER_0_34_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22580_ _09422_ _09731_ _09472_ VGND VGND VPWR VPWR _09732_ sky130_fd_sc_hd__o21ai_1
X_31778_ clknet_leaf_255_clk _03232_ VGND VGND VPWR VPWR datamem.data_ram\[6\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_217_5699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_4670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_174_4681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21531_ _08627_ _08780_ _08782_ _08784_ VGND VGND VPWR VPWR _08785_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_35_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30729_ clknet_leaf_219_clk _02464_ VGND VGND VPWR VPWR datamem.data_ram\[48\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23693__288 clknet_1_1__leaf__10195_ VGND VGND VPWR VPWR net414 sky130_fd_sc_hd__inv_2
XFILLER_0_1_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_4567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_185_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_4578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24250_ _10296_ VGND VGND VPWR VPWR _02243_ sky130_fd_sc_hd__clkbuf_1
X_21462_ _08565_ _08717_ _08719_ _08652_ VGND VGND VPWR VPWR _08720_ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23201_ _10121_ VGND VGND VPWR VPWR _01369_ sky130_fd_sc_hd__clkbuf_1
X_20413_ datamem.data_ram\[58\]\[12\] _06609_ _06617_ datamem.data_ram\[60\]\[12\]
+ _06598_ VGND VGND VPWR VPWR _07705_ sky130_fd_sc_hd__o221a_1
X_21393_ _08643_ _08647_ _08653_ _08625_ VGND VGND VPWR VPWR _01029_ sky130_fd_sc_hd__o31a_1
XFILLER_0_4_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20344_ _06607_ VGND VGND VPWR VPWR _07636_ sky130_fd_sc_hd__buf_6
XFILLER_0_144_1040 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23063_ _09299_ _10092_ _09361_ VGND VGND VPWR VPWR _10093_ sky130_fd_sc_hd__a21oi_4
X_27940_ _12422_ VGND VGND VPWR VPWR _03807_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_73_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20275_ datamem.data_ram\[46\]\[19\] _06764_ _06700_ datamem.data_ram\[41\]\[19\]
+ VGND VGND VPWR VPWR _07568_ sky130_fd_sc_hd__o22a_1
XFILLER_0_222_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3210 rvcpu.dp.rf.reg_file_arr\[2\]\[28\] VGND VGND VPWR VPWR net4360 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3221 datamem.data_ram\[61\]\[18\] VGND VGND VPWR VPWR net4371 sky130_fd_sc_hd__dlygate4sd3_1
X_22014_ _09241_ VGND VGND VPWR VPWR _01062_ sky130_fd_sc_hd__clkbuf_1
Xhold3232 rvcpu.dp.rf.reg_file_arr\[29\]\[24\] VGND VGND VPWR VPWR net4382 sky130_fd_sc_hd__dlygate4sd3_1
X_27871_ _12384_ VGND VGND VPWR VPWR _03776_ sky130_fd_sc_hd__clkbuf_1
Xhold3243 rvcpu.dp.rf.reg_file_arr\[16\]\[2\] VGND VGND VPWR VPWR net4393 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3254 datamem.data_ram\[28\]\[27\] VGND VGND VPWR VPWR net4404 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2520 datamem.data_ram\[53\]\[16\] VGND VGND VPWR VPWR net3670 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3265 datamem.data_ram\[2\]\[20\] VGND VGND VPWR VPWR net4415 sky130_fd_sc_hd__dlygate4sd3_1
X_26822_ _11681_ _11774_ VGND VGND VPWR VPWR _11777_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_251_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_251_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold2531 datamem.data_ram\[26\]\[10\] VGND VGND VPWR VPWR net3681 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3276 rvcpu.dp.rf.reg_file_arr\[24\]\[15\] VGND VGND VPWR VPWR net4426 sky130_fd_sc_hd__dlygate4sd3_1
X_29610_ net964 _01345_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[25\]\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_142_3902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3287 rvcpu.dp.rf.reg_file_arr\[24\]\[9\] VGND VGND VPWR VPWR net4437 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2542 datamem.data_ram\[48\]\[25\] VGND VGND VPWR VPWR net3692 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3298 rvcpu.dp.plfd.InstrD\[9\] VGND VGND VPWR VPWR net4448 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2553 datamem.data_ram\[41\]\[19\] VGND VGND VPWR VPWR net3703 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2564 datamem.data_ram\[39\]\[29\] VGND VGND VPWR VPWR net3714 sky130_fd_sc_hd__dlygate4sd3_1
X_29541_ net895 _01276_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[27\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_32_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1830 datamem.data_ram\[15\]\[28\] VGND VGND VPWR VPWR net2980 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2575 datamem.data_ram\[59\]\[24\] VGND VGND VPWR VPWR net3725 sky130_fd_sc_hd__dlygate4sd3_1
X_26753_ _11734_ VGND VGND VPWR VPWR _03308_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_32_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1841 datamem.data_ram\[31\]\[11\] VGND VGND VPWR VPWR net2991 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2586 datamem.data_ram\[21\]\[14\] VGND VGND VPWR VPWR net3736 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23965_ _10236_ VGND VGND VPWR VPWR _02018_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_32_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2597 rvcpu.dp.rf.reg_file_arr\[10\]\[11\] VGND VGND VPWR VPWR net3747 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1852 datamem.data_ram\[58\]\[28\] VGND VGND VPWR VPWR net3002 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1863 rvcpu.dp.rf.reg_file_arr\[6\]\[14\] VGND VGND VPWR VPWR net3013 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1874 datamem.data_ram\[44\]\[19\] VGND VGND VPWR VPWR net3024 sky130_fd_sc_hd__dlygate4sd3_1
X_25704_ _11125_ VGND VGND VPWR VPWR _02868_ sky130_fd_sc_hd__clkbuf_1
X_22916_ _09217_ _09262_ _09220_ VGND VGND VPWR VPWR _10050_ sky130_fd_sc_hd__a21o_2
Xhold1885 rvcpu.dp.rf.reg_file_arr\[28\]\[12\] VGND VGND VPWR VPWR net3035 sky130_fd_sc_hd__dlygate4sd3_1
X_29472_ net834 _01207_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[2\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26684_ _11679_ _11694_ VGND VGND VPWR VPWR _11696_ sky130_fd_sc_hd__and2_1
Xhold1896 rvcpu.dp.rf.reg_file_arr\[17\]\[8\] VGND VGND VPWR VPWR net3046 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28423_ _12689_ VGND VGND VPWR VPWR _04023_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25635_ _10063_ VGND VGND VPWR VPWR _11086_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_195_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22847_ _09469_ _09984_ VGND VGND VPWR VPWR _09985_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28354_ _12450_ net3607 net95 VGND VGND VPWR VPWR _12652_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25566_ _11018_ net1485 _11041_ _11043_ VGND VGND VPWR VPWR _02812_ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22778_ rvcpu.dp.rf.reg_file_arr\[16\]\[25\] rvcpu.dp.rf.reg_file_arr\[17\]\[25\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[25\] rvcpu.dp.rf.reg_file_arr\[19\]\[25\] _09445_
+ _09447_ VGND VGND VPWR VPWR _09919_ sky130_fd_sc_hd__mux4_1
XFILLER_0_94_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27305_ _12061_ net1789 _12065_ _12067_ VGND VGND VPWR VPWR _03527_ sky130_fd_sc_hd__a31o_1
XFILLER_0_183_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24517_ _10452_ net4441 _10440_ VGND VGND VPWR VPWR _10453_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28285_ _12433_ net3240 _12613_ VGND VGND VPWR VPWR _12615_ sky130_fd_sc_hd__mux2_1
X_21729_ _08725_ _08972_ VGND VGND VPWR VPWR _08973_ sky130_fd_sc_hd__nor2_1
X_25497_ _11003_ VGND VGND VPWR VPWR _02783_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15250_ _13638_ _13789_ VGND VGND VPWR VPWR _13790_ sky130_fd_sc_hd__nand2_1
X_27236_ _10268_ _10921_ _10922_ VGND VGND VPWR VPWR _12031_ sky130_fd_sc_hd__and3_1
XFILLER_0_164_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24448_ _10056_ datamem.data_ram\[53\]\[2\] _10404_ _10411_ VGND VGND VPWR VPWR _02326_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23220__870 clknet_1_0__leaf__10124_ VGND VGND VPWR VPWR net996 sky130_fd_sc_hd__inv_2
X_15181_ _13719_ _13720_ _13723_ _13412_ VGND VGND VPWR VPWR _13724_ sky130_fd_sc_hd__a31o_1
X_27167_ _11974_ net1496 _11983_ _11989_ VGND VGND VPWR VPWR _03467_ sky130_fd_sc_hd__a31o_1
XFILLER_0_152_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24379_ _10368_ VGND VGND VPWR VPWR _02300_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26118_ _11394_ VGND VGND VPWR VPWR _03012_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27098_ _11938_ net1786 _11940_ _11945_ VGND VGND VPWR VPWR _03442_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_39_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26049_ _11104_ VGND VGND VPWR VPWR _11353_ sky130_fd_sc_hd__clkbuf_4
X_18940_ _05525_ _05531_ _05537_ _05552_ VGND VGND VPWR VPWR _06278_ sky130_fd_sc_hd__a31o_1
XFILLER_0_63_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_1232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_148_Right_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18871_ _05619_ _06213_ _06055_ VGND VGND VPWR VPWR _06214_ sky130_fd_sc_hd__o21a_1
XFILLER_0_218_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_242_clk clknet_5_17__leaf_clk VGND VGND VPWR VPWR clknet_leaf_242_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_219_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17822_ _13200_ rvcpu.dp.plde.RD2E\[25\] _05196_ VGND VGND VPWR VPWR _05209_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29808_ net1146 _01543_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[1\]\[3\] sky130_fd_sc_hd__dfxtp_1
Xhold4 rvcpu.dp.plde.RegWriteE VGND VGND VPWR VPWR net1154 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_176_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14965_ _13311_ _13513_ VGND VGND VPWR VPWR _13514_ sky130_fd_sc_hd__nor2_4
X_29739_ net1085 _01474_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[21\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_17753_ _13278_ net3451 _05117_ VGND VGND VPWR VPWR _05152_ sky130_fd_sc_hd__mux2_1
XFILLER_0_221_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24156__659 clknet_1_1__leaf__10263_ VGND VGND VPWR VPWR net785 sky130_fd_sc_hd__inv_2
X_16704_ _14168_ net3629 _04587_ VGND VGND VPWR VPWR _04596_ sky130_fd_sc_hd__mux2_1
X_32750_ clknet_leaf_237_clk _04172_ VGND VGND VPWR VPWR datamem.data_ram\[15\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_17684_ _05115_ VGND VGND VPWR VPWR _01197_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_226_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14896_ _13446_ VGND VGND VPWR VPWR _13447_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_187_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31701_ clknet_leaf_43_clk _03159_ VGND VGND VPWR VPWR rvcpu.dp.pcreg.q\[19\] sky130_fd_sc_hd__dfxtp_1
X_19423_ _06718_ VGND VGND VPWR VPWR _06719_ sky130_fd_sc_hd__buf_8
X_16635_ _04559_ VGND VGND VPWR VPWR _01722_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32681_ clknet_leaf_80_clk _04103_ VGND VGND VPWR VPWR datamem.data_ram\[18\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31632_ clknet_leaf_52_clk net1228 VGND VGND VPWR VPWR rvcpu.dp.plmw.lAuiPCW\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19354_ _05185_ net1 VGND VGND VPWR VPWR _06650_ sky130_fd_sc_hd__nor2_2
X_16566_ _04522_ VGND VGND VPWR VPWR _01762_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_186_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15517_ _13659_ _14043_ VGND VGND VPWR VPWR _14044_ sky130_fd_sc_hd__or2b_1
X_18305_ _05669_ VGND VGND VPWR VPWR _05670_ sky130_fd_sc_hd__clkbuf_4
X_31563_ clknet_leaf_74_clk datamem.rd_data_mem\[13\] VGND VGND VPWR VPWR rvcpu.dp.plmw.ReadDataW\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19285_ rvcpu.dp.plem.funct3M\[0\] rvcpu.dp.plem.funct3M\[2\] rvcpu.dp.plem.funct3M\[1\]
+ VGND VGND VPWR VPWR _06581_ sky130_fd_sc_hd__or3b_1
XPHY_EDGE_ROW_99_Left_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16497_ net3688 _14457_ _04478_ VGND VGND VPWR VPWR _04486_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18236_ _05427_ _05431_ VGND VGND VPWR VPWR _05601_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30514_ clknet_leaf_205_clk _02249_ VGND VGND VPWR VPWR datamem.data_ram\[56\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15448_ _13969_ _13972_ _13521_ _13978_ VGND VGND VPWR VPWR _13979_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_212_5574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31494_ clknet_leaf_44_clk rvcpu.dp.lAuiPCE\[20\] VGND VGND VPWR VPWR rvcpu.dp.plem.lAuiPCM\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_212_5585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18167_ rvcpu.dp.plem.ALUResultM\[24\] _05293_ _05294_ _13203_ VGND VGND VPWR VPWR
+ _05532_ sky130_fd_sc_hd__o22a_1
XFILLER_0_4_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30445_ net783 _02180_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[29\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_15379_ _13308_ _13767_ _13357_ _13654_ VGND VGND VPWR VPWR _13913_ sky130_fd_sc_hd__or4_1
XFILLER_0_4_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold404 datamem.data_ram\[5\]\[5\] VGND VGND VPWR VPWR net1554 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17118_ _14172_ net4370 _04815_ VGND VGND VPWR VPWR _04816_ sky130_fd_sc_hd__mux2_1
Xhold415 datamem.data_ram\[33\]\[0\] VGND VGND VPWR VPWR net1565 sky130_fd_sc_hd__dlygate4sd3_1
X_18098_ _05463_ _05464_ VGND VGND VPWR VPWR _05466_ sky130_fd_sc_hd__and2_1
X_30376_ net722 _02111_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[3\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_225_5902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold426 datamem.data_ram\[50\]\[7\] VGND VGND VPWR VPWR net1576 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold437 datamem.data_ram\[29\]\[3\] VGND VGND VPWR VPWR net1587 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold448 datamem.data_ram\[55\]\[1\] VGND VGND VPWR VPWR net1598 sky130_fd_sc_hd__dlygate4sd3_1
X_32115_ clknet_leaf_97_clk _03537_ VGND VGND VPWR VPWR datamem.data_ram\[0\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_146_4002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold459 datamem.data_ram\[55\]\[7\] VGND VGND VPWR VPWR net1609 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17049_ _04756_ VGND VGND VPWR VPWR _04779_ sky130_fd_sc_hd__buf_4
X_23729__321 clknet_1_1__leaf__10198_ VGND VGND VPWR VPWR net447 sky130_fd_sc_hd__inv_2
XFILLER_0_99_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32046_ clknet_leaf_131_clk _03468_ VGND VGND VPWR VPWR datamem.data_ram\[49\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_115_Right_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20060_ datamem.data_ram\[62\]\[26\] _06743_ _06704_ datamem.data_ram\[63\]\[26\]
+ _06598_ VGND VGND VPWR VPWR _07354_ sky130_fd_sc_hd__o221a_1
XFILLER_0_209_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_221_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_233_clk clknet_5_20__leaf_clk VGND VGND VPWR VPWR clknet_leaf_233_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold1104 rvcpu.dp.rf.reg_file_arr\[8\]\[28\] VGND VGND VPWR VPWR net2254 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1115 rvcpu.dp.rf.reg_file_arr\[16\]\[13\] VGND VGND VPWR VPWR net2265 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1126 datamem.data_ram\[12\]\[22\] VGND VGND VPWR VPWR net2276 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1137 rvcpu.dp.rf.reg_file_arr\[10\]\[23\] VGND VGND VPWR VPWR net2287 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1148 rvcpu.dp.rf.reg_file_arr\[10\]\[19\] VGND VGND VPWR VPWR net2298 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_105_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1159 datamem.data_ram\[12\]\[21\] VGND VGND VPWR VPWR net2309 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_176_4710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20962_ datamem.data_ram\[59\]\[15\] _06631_ _08250_ _06922_ VGND VGND VPWR VPWR
+ _08251_ sky130_fd_sc_hd__o22a_1
X_32948_ clknet_leaf_215_clk _04370_ VGND VGND VPWR VPWR datamem.data_ram\[6\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_176_4721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22701_ _09481_ _09846_ VGND VGND VPWR VPWR _09847_ sky130_fd_sc_hd__and2_1
XFILLER_0_178_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_923 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32879_ clknet_leaf_56_clk _04301_ VGND VGND VPWR VPWR datamem.data_ram\[10\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_20893_ _05391_ _06586_ _08123_ _08182_ _07120_ VGND VGND VPWR VPWR _08183_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_66_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25420_ _10760_ net3501 _10961_ VGND VGND VPWR VPWR _10966_ sky130_fd_sc_hd__mux2_1
X_23163__835 clknet_1_1__leaf__10110_ VGND VGND VPWR VPWR net961 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_172_4618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22632_ _09516_ _09780_ VGND VGND VPWR VPWR _09781_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_172_4629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23701__295 clknet_1_0__leaf__10196_ VGND VGND VPWR VPWR net421 sky130_fd_sc_hd__inv_2
XFILLER_0_76_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23775__363 clknet_1_0__leaf__10202_ VGND VGND VPWR VPWR net489 sky130_fd_sc_hd__inv_2
XFILLER_0_48_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25351_ _10876_ net1393 _10920_ _10924_ VGND VGND VPWR VPWR _02716_ sky130_fd_sc_hd__a31o_1
XFILLER_0_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22563_ _09400_ VGND VGND VPWR VPWR _09716_ sky130_fd_sc_hd__buf_4
XFILLER_0_10_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24302_ _10324_ VGND VGND VPWR VPWR _02267_ sky130_fd_sc_hd__clkbuf_1
X_28070_ _12369_ net3735 _12492_ VGND VGND VPWR VPWR _12499_ sky130_fd_sc_hd__mux2_1
X_21514_ rvcpu.dp.rf.reg_file_arr\[4\]\[7\] rvcpu.dp.rf.reg_file_arr\[5\]\[7\] rvcpu.dp.rf.reg_file_arr\[6\]\[7\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[7\] _08551_ _08555_ VGND VGND VPWR VPWR _08769_ sky130_fd_sc_hd__mux4_1
XFILLER_0_134_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25282_ _10883_ VGND VGND VPWR VPWR _02688_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22494_ _09476_ _09648_ _09650_ _09474_ VGND VGND VPWR VPWR _09651_ sky130_fd_sc_hd__o211a_1
X_27021_ _10051_ VGND VGND VPWR VPWR _11898_ sky130_fd_sc_hd__buf_2
XFILLER_0_44_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_185_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24233_ _10287_ VGND VGND VPWR VPWR _02235_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_75_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21445_ _08535_ VGND VGND VPWR VPWR _08703_ sky130_fd_sc_hd__buf_4
XFILLER_0_72_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_131_3636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_3647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21376_ _08636_ VGND VGND VPWR VPWR _08637_ sky130_fd_sc_hd__buf_4
XFILLER_0_222_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20327_ datamem.data_ram\[16\]\[4\] _07138_ _06977_ datamem.data_ram\[20\]\[4\] _07618_
+ VGND VGND VPWR VPWR _07619_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28972_ _12727_ net1769 _12988_ _12994_ VGND VGND VPWR VPWR _04267_ sky130_fd_sc_hd__a31o_1
XFILLER_0_102_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold960 rvcpu.dp.rf.reg_file_arr\[3\]\[11\] VGND VGND VPWR VPWR net2110 sky130_fd_sc_hd__dlygate4sd3_1
Xhold971 datamem.data_ram\[58\]\[15\] VGND VGND VPWR VPWR net2121 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold982 datamem.data_ram\[2\]\[13\] VGND VGND VPWR VPWR net2132 sky130_fd_sc_hd__dlygate4sd3_1
X_20258_ _07071_ _07534_ _07539_ _07550_ VGND VGND VPWR VPWR _07551_ sky130_fd_sc_hd__a31o_1
X_27923_ _12413_ VGND VGND VPWR VPWR _03799_ sky130_fd_sc_hd__clkbuf_1
Xhold993 datamem.data_ram\[39\]\[23\] VGND VGND VPWR VPWR net2143 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_34_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3040 datamem.data_ram\[14\]\[12\] VGND VGND VPWR VPWR net4190 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3051 rvcpu.dp.rf.reg_file_arr\[9\]\[14\] VGND VGND VPWR VPWR net4201 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_224_clk clknet_5_21__leaf_clk VGND VGND VPWR VPWR clknet_leaf_224_clk
+ sky130_fd_sc_hd__clkbuf_8
X_27854_ _12375_ VGND VGND VPWR VPWR _03768_ sky130_fd_sc_hd__clkbuf_1
Xhold3062 datamem.data_ram\[42\]\[28\] VGND VGND VPWR VPWR net4212 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20189_ _07476_ _07481_ _06596_ VGND VGND VPWR VPWR _07482_ sky130_fd_sc_hd__o21a_1
Xhold3073 rvcpu.dp.rf.reg_file_arr\[2\]\[29\] VGND VGND VPWR VPWR net4223 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold3084 rvcpu.dp.rf.reg_file_arr\[23\]\[18\] VGND VGND VPWR VPWR net4234 sky130_fd_sc_hd__dlygate4sd3_1
X_23431__83 clknet_1_1__leaf__10154_ VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__inv_2
XFILLER_0_216_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2350 datamem.data_ram\[6\]\[21\] VGND VGND VPWR VPWR net3500 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3095 rvcpu.dp.plfd.InstrD\[2\] VGND VGND VPWR VPWR net4245 sky130_fd_sc_hd__dlygate4sd3_1
X_26805_ _11753_ net1427 _11761_ _11766_ VGND VGND VPWR VPWR _03328_ sky130_fd_sc_hd__a31o_1
Xhold2361 rvcpu.dp.rf.reg_file_arr\[15\]\[24\] VGND VGND VPWR VPWR net3511 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2372 datamem.data_ram\[51\]\[17\] VGND VGND VPWR VPWR net3522 sky130_fd_sc_hd__dlygate4sd3_1
X_27785_ _12333_ VGND VGND VPWR VPWR _03741_ sky130_fd_sc_hd__clkbuf_1
X_24997_ _10719_ VGND VGND VPWR VPWR _02567_ sky130_fd_sc_hd__clkbuf_1
Xhold2383 rvcpu.dp.rf.reg_file_arr\[22\]\[1\] VGND VGND VPWR VPWR net3533 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2394 datamem.data_ram\[7\]\[18\] VGND VGND VPWR VPWR net3544 sky130_fd_sc_hd__dlygate4sd3_1
X_23481__128 clknet_1_1__leaf__10159_ VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__inv_2
XFILLER_0_99_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1660 rvcpu.dp.rf.reg_file_arr\[1\]\[15\] VGND VGND VPWR VPWR net2810 sky130_fd_sc_hd__dlygate4sd3_1
X_14750_ _13284_ VGND VGND VPWR VPWR _13303_ sky130_fd_sc_hd__buf_4
X_26736_ _09227_ VGND VGND VPWR VPWR _11725_ sky130_fd_sc_hd__buf_2
Xhold1671 datamem.data_ram\[36\]\[16\] VGND VGND VPWR VPWR net2821 sky130_fd_sc_hd__dlygate4sd3_1
X_29524_ net886 _01259_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[28\]\[31\] sky130_fd_sc_hd__dfxtp_1
Xhold1682 datamem.data_ram\[44\]\[29\] VGND VGND VPWR VPWR net2832 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1693 datamem.data_ram\[24\]\[20\] VGND VGND VPWR VPWR net2843 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29455_ net817 _01190_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[30\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26667_ _11684_ _11677_ VGND VGND VPWR VPWR _11685_ sky130_fd_sc_hd__and2_1
XFILLER_0_196_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14681_ net2194 _13244_ _13245_ VGND VGND VPWR VPWR _13246_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_917 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16420_ _14576_ VGND VGND VPWR VPWR _01830_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0__10267_ _10267_ VGND VGND VPWR VPWR clknet_0__10267_ sky130_fd_sc_hd__clkbuf_16
X_28406_ _12450_ net2752 _12678_ VGND VGND VPWR VPWR _12680_ sky130_fd_sc_hd__mux2_1
X_25618_ _11073_ VGND VGND VPWR VPWR _02834_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_196_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_184_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29386_ clknet_leaf_269_clk _01121_ VGND VGND VPWR VPWR datamem.data_ram\[60\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_26598_ _11618_ net1771 _11639_ _11646_ VGND VGND VPWR VPWR _03241_ sky130_fd_sc_hd__a31o_1
XFILLER_0_67_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28337_ _12433_ net3529 _12641_ VGND VGND VPWR VPWR _12643_ sky130_fd_sc_hd__mux2_1
X_16351_ net2202 _14449_ _14536_ VGND VGND VPWR VPWR _14540_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25549_ _10756_ net4172 _11030_ VGND VGND VPWR VPWR _11033_ sky130_fd_sc_hd__mux2_1
Xclkbuf_0__10198_ _10198_ VGND VGND VPWR VPWR clknet_0__10198_ sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15302_ _13385_ _13836_ _13837_ _13374_ _13839_ VGND VGND VPWR VPWR _13840_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_229_6002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19070_ _06394_ _06395_ VGND VGND VPWR VPWR _06396_ sky130_fd_sc_hd__nand2_1
XFILLER_0_183_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16282_ _14503_ VGND VGND VPWR VPWR _01895_ sky130_fd_sc_hd__clkbuf_1
X_28268_ _12605_ VGND VGND VPWR VPWR _03952_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_229_6013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_217_Right_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_229_6024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18021_ rvcpu.dp.plem.ALUResultM\[0\] VGND VGND VPWR VPWR _05391_ sky130_fd_sc_hd__inv_2
XFILLER_0_212_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27219_ _11968_ _12019_ VGND VGND VPWR VPWR _12021_ sky130_fd_sc_hd__and2_1
X_15233_ _13378_ _13773_ _13442_ VGND VGND VPWR VPWR _13774_ sky130_fd_sc_hd__or3_1
XFILLER_0_180_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28199_ _12567_ VGND VGND VPWR VPWR _03921_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30230_ net584 _01965_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[7\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_15164_ _13674_ _13707_ VGND VGND VPWR VPWR _13708_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30161_ net523 _01896_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[0\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_15095_ _13304_ _13589_ VGND VGND VPWR VPWR _13640_ sky130_fd_sc_hd__and2_1
X_19972_ datamem.data_ram\[26\]\[18\] _06690_ _06633_ datamem.data_ram\[27\]\[18\]
+ _06600_ VGND VGND VPWR VPWR _07266_ sky130_fd_sc_hd__o221a_1
XFILLER_0_50_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18923_ _05239_ _06249_ _06250_ _06254_ _06262_ VGND VGND VPWR VPWR rvcpu.ALUResultE\[24\]
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_157_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30092_ net454 _01827_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[11\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_219_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_215_clk clknet_5_20__leaf_clk VGND VGND VPWR VPWR clknet_leaf_215_clk
+ sky130_fd_sc_hd__clkbuf_8
X_23945__499 clknet_1_1__leaf__10228_ VGND VGND VPWR VPWR net625 sky130_fd_sc_hd__inv_2
XFILLER_0_206_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18854_ _05480_ _05785_ _06108_ _05479_ VGND VGND VPWR VPWR _06198_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_59_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17805_ rvcpu.dp.plem.ALUResultM\[31\] _05197_ _05178_ VGND VGND VPWR VPWR _05198_
+ sky130_fd_sc_hd__mux2_1
X_18785_ _05454_ _05513_ _05886_ VGND VGND VPWR VPWR _06133_ sky130_fd_sc_hd__a21o_1
X_15997_ _14336_ VGND VGND VPWR VPWR _02029_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_207_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32802_ clknet_leaf_156_clk _04224_ VGND VGND VPWR VPWR datamem.data_ram\[13\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_14948_ _13493_ _13495_ _13496_ VGND VGND VPWR VPWR _13497_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_167_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17736_ _05143_ VGND VGND VPWR VPWR _01173_ sky130_fd_sc_hd__clkbuf_1
X_30994_ clknet_leaf_102_clk _02729_ VGND VGND VPWR VPWR datamem.data_ram\[13\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32733_ clknet_leaf_78_clk _04155_ VGND VGND VPWR VPWR datamem.data_ram\[16\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_14879_ _13430_ VGND VGND VPWR VPWR _13431_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_212_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17667_ net4070 _13250_ _05104_ VGND VGND VPWR VPWR _05107_ sky130_fd_sc_hd__mux2_1
X_19406_ _06662_ VGND VGND VPWR VPWR _06702_ sky130_fd_sc_hd__buf_6
XFILLER_0_187_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16618_ _04550_ VGND VGND VPWR VPWR _01730_ sky130_fd_sc_hd__clkbuf_1
X_23227__876 clknet_1_0__leaf__10125_ VGND VGND VPWR VPWR net1002 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_214_5625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32664_ clknet_leaf_171_clk _04086_ VGND VGND VPWR VPWR datamem.data_ram\[19\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_17598_ _05070_ VGND VGND VPWR VPWR _01238_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_214_5636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19337_ _06632_ VGND VGND VPWR VPWR _06633_ sky130_fd_sc_hd__buf_6
X_31615_ clknet_leaf_14_clk net1256 VGND VGND VPWR VPWR rvcpu.dp.plmw.RdW\[1\] sky130_fd_sc_hd__dfxtp_4
X_16549_ _04513_ VGND VGND VPWR VPWR _01770_ sky130_fd_sc_hd__clkbuf_1
X_32595_ clknet_leaf_251_clk _04017_ VGND VGND VPWR VPWR datamem.data_ram\[21\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19268_ rvcpu.dp.plfd.InstrD\[14\] VGND VGND VPWR VPWR _06568_ sky130_fd_sc_hd__inv_2
X_31546_ clknet_leaf_17_clk net1259 VGND VGND VPWR VPWR rvcpu.dp.plem.RdM\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18219_ _05374_ _05377_ VGND VGND VPWR VPWR _05584_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31477_ clknet_leaf_65_clk rvcpu.dp.lAuiPCE\[3\] VGND VGND VPWR VPWR rvcpu.dp.plem.lAuiPCM\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_19199_ _06507_ _06508_ VGND VGND VPWR VPWR _06509_ sky130_fd_sc_hd__or2b_1
XFILLER_0_26_683 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21230_ datamem.data_ram\[52\]\[29\] datamem.data_ram\[52\]\[21\] datamem.data_ram\[53\]\[13\]
+ datamem.data_ram\[52\]\[13\] VGND VGND VPWR VPWR _08493_ sky130_fd_sc_hd__or4_1
XFILLER_0_206_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30428_ net766 _02163_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[29\]\[7\] sky130_fd_sc_hd__dfxtp_1
Xhold201 datamem.data_ram\[34\]\[6\] VGND VGND VPWR VPWR net1351 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold212 rvcpu.dp.pcreg.q\[16\] VGND VGND VPWR VPWR net1362 sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 datamem.data_ram\[14\]\[7\] VGND VGND VPWR VPWR net1373 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold234 datamem.data_ram\[2\]\[7\] VGND VGND VPWR VPWR net1384 sky130_fd_sc_hd__dlygate4sd3_1
X_21161_ datamem.data_ram\[4\]\[23\] datamem.data_ram\[5\]\[23\] _07911_ VGND VGND
+ VPWR VPWR _08450_ sky130_fd_sc_hd__mux2_1
Xhold245 datamem.data_ram\[59\]\[5\] VGND VGND VPWR VPWR net1395 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30359_ net705 _02094_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[3\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold256 datamem.data_ram\[0\]\[0\] VGND VGND VPWR VPWR net1406 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold267 datamem.data_ram\[6\]\[7\] VGND VGND VPWR VPWR net1417 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_165_4444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold278 datamem.data_ram\[21\]\[5\] VGND VGND VPWR VPWR net1428 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_165_4455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20112_ datamem.data_ram\[29\]\[10\] _06723_ _06686_ datamem.data_ram\[28\]\[10\]
+ VGND VGND VPWR VPWR _07406_ sky130_fd_sc_hd__o22a_1
Xhold289 datamem.data_ram\[59\]\[4\] VGND VGND VPWR VPWR net1439 sky130_fd_sc_hd__dlygate4sd3_1
X_21092_ datamem.data_ram\[2\]\[7\] datamem.data_ram\[3\]\[7\] _07912_ VGND VGND VPWR
+ VPWR _08381_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_165_4466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_206_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_206_clk
+ sky130_fd_sc_hd__clkbuf_8
X_32029_ clknet_leaf_128_clk _03451_ VGND VGND VPWR VPWR datamem.data_ram\[26\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_24920_ _10113_ _10601_ _10611_ VGND VGND VPWR VPWR _10678_ sky130_fd_sc_hd__a21oi_1
X_20043_ datamem.data_ram\[5\]\[26\] _06722_ _07335_ _07336_ VGND VGND VPWR VPWR _07337_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24851_ _10598_ _10640_ _10611_ VGND VGND VPWR VPWR _10641_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_226_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_124_3462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27570_ _12218_ VGND VGND VPWR VPWR _03641_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_124_3473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24782_ _10603_ VGND VGND VPWR VPWR _02468_ sky130_fd_sc_hd__clkbuf_1
X_21994_ _09223_ VGND VGND VPWR VPWR _09224_ sky130_fd_sc_hd__clkbuf_2
XANTENNA_107 _07023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_197_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26521_ _10058_ _11604_ _11605_ net1434 VGND VGND VPWR VPWR _03205_ sky130_fd_sc_hd__a22o_1
XANTENNA_118 _07191_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_178_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23733_ clknet_1_1__leaf__10192_ VGND VGND VPWR VPWR _10199_ sky130_fd_sc_hd__buf_1
XANTENNA_129 _07808_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_200_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20945_ datamem.data_ram\[62\]\[22\] _07860_ _07863_ datamem.data_ram\[60\]\[22\]
+ _08234_ VGND VGND VPWR VPWR _08235_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23699__294 clknet_1_0__leaf__10195_ VGND VGND VPWR VPWR net420 sky130_fd_sc_hd__inv_2
X_29240_ _09329_ net2453 _13132_ VGND VGND VPWR VPWR _13140_ sky130_fd_sc_hd__mux2_1
X_26452_ _11576_ _11215_ _11540_ _06505_ _11579_ VGND VGND VPWR VPWR _11580_ sky130_fd_sc_hd__a221o_1
XFILLER_0_163_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20876_ _05347_ _08159_ _08163_ _08165_ _08124_ VGND VGND VPWR VPWR _08166_ sky130_fd_sc_hd__a221o_1
XFILLER_0_166_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25403_ _10954_ net1638 _10949_ _10956_ VGND VGND VPWR VPWR _02736_ sky130_fd_sc_hd__a31o_1
XFILLER_0_138_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_193_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29171_ _13102_ VGND VGND VPWR VPWR _04358_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_27_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22615_ rvcpu.dp.rf.reg_file_arr\[24\]\[16\] rvcpu.dp.rf.reg_file_arr\[25\]\[16\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[16\] rvcpu.dp.rf.reg_file_arr\[27\]\[16\] _09392_
+ _09394_ VGND VGND VPWR VPWR _09765_ sky130_fd_sc_hd__mux4_1
X_26383_ _11150_ _11529_ VGND VGND VPWR VPWR _11530_ sky130_fd_sc_hd__and2_1
XFILLER_0_113_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28122_ _12526_ VGND VGND VPWR VPWR _03885_ sky130_fd_sc_hd__clkbuf_1
X_25334_ _10758_ net2768 _10909_ VGND VGND VPWR VPWR _10913_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22546_ rvcpu.dp.rf.reg_file_arr\[8\]\[12\] rvcpu.dp.rf.reg_file_arr\[10\]\[12\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[12\] rvcpu.dp.rf.reg_file_arr\[11\]\[12\] _09608_
+ _09532_ VGND VGND VPWR VPWR _09700_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_98_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_98_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28053_ _12460_ net2266 net96 VGND VGND VPWR VPWR _12490_ sky130_fd_sc_hd__mux2_1
X_25265_ _10416_ _10868_ VGND VGND VPWR VPWR _10874_ sky130_fd_sc_hd__and2_1
X_22477_ rvcpu.dp.rf.reg_file_arr\[20\]\[9\] rvcpu.dp.rf.reg_file_arr\[21\]\[9\] rvcpu.dp.rf.reg_file_arr\[22\]\[9\]
+ rvcpu.dp.rf.reg_file_arr\[23\]\[9\] _09434_ _09558_ VGND VGND VPWR VPWR _09634_
+ sky130_fd_sc_hd__mux4_1
X_27004_ _11825_ _11886_ VGND VGND VPWR VPWR _11888_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_94_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24216_ _10278_ VGND VGND VPWR VPWR _02227_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21428_ _08535_ VGND VGND VPWR VPWR _08687_ sky130_fd_sc_hd__buf_6
X_25196_ _10737_ net2595 _10829_ VGND VGND VPWR VPWR _10836_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_80_Right_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21359_ rvcpu.dp.plde.JumpE rvcpu.dp.plde.JalrE VGND VGND VPWR VPWR _08621_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_57_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24078_ _09273_ net4151 _10249_ VGND VGND VPWR VPWR _10251_ sky130_fd_sc_hd__mux2_1
X_28955_ _12984_ VGND VGND VPWR VPWR _04260_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold790 datamem.data_ram\[17\]\[30\] VGND VGND VPWR VPWR net1940 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23332__971 clknet_1_0__leaf__10135_ VGND VGND VPWR VPWR net1097 sky130_fd_sc_hd__inv_2
XFILLER_0_120_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27906_ _12404_ VGND VGND VPWR VPWR _03791_ sky130_fd_sc_hd__clkbuf_1
X_15920_ _14295_ VGND VGND VPWR VPWR _02065_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_53_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28886_ _12947_ VGND VGND VPWR VPWR _04228_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15851_ _14257_ VGND VGND VPWR VPWR _02096_ sky130_fd_sc_hd__clkbuf_1
X_27837_ _12364_ VGND VGND VPWR VPWR _03762_ sky130_fd_sc_hd__clkbuf_1
Xhold2180 datamem.data_ram\[45\]\[24\] VGND VGND VPWR VPWR net3330 sky130_fd_sc_hd__dlygate4sd3_1
X_14802_ _13344_ _13351_ _13354_ VGND VGND VPWR VPWR _13355_ sky130_fd_sc_hd__a21oi_1
Xhold2191 datamem.data_ram\[60\]\[26\] VGND VGND VPWR VPWR net3341 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_189_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18570_ _05910_ _05911_ _05929_ VGND VGND VPWR VPWR _05930_ sky130_fd_sc_hd__a21bo_1
X_15782_ _14220_ VGND VGND VPWR VPWR _02136_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27768_ _12157_ net4177 _12316_ VGND VGND VPWR VPWR _12324_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_207_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1490 datamem.data_ram\[35\]\[29\] VGND VGND VPWR VPWR net2640 sky130_fd_sc_hd__dlygate4sd3_1
X_14733_ rvcpu.dp.pcreg.q\[4\] VGND VGND VPWR VPWR _13286_ sky130_fd_sc_hd__buf_2
X_29507_ net869 _01242_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[28\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_17521_ _05029_ VGND VGND VPWR VPWR _01282_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_207_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26719_ _11715_ VGND VGND VPWR VPWR _03293_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27699_ _12287_ VGND VGND VPWR VPWR _03701_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17452_ _14166_ net3973 _04985_ VGND VGND VPWR VPWR _04993_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14664_ net1882 _13232_ _13214_ VGND VGND VPWR VPWR _13233_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1__f__10219_ clknet_0__10219_ VGND VGND VPWR VPWR clknet_1_1__leaf__10219_
+ sky130_fd_sc_hd__clkbuf_16
X_29438_ net800 _01173_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[30\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_200_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16403_ _14567_ VGND VGND VPWR VPWR _01838_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_223_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17383_ _04956_ VGND VGND VPWR VPWR _01347_ sky130_fd_sc_hd__clkbuf_1
X_14595_ _13177_ _13179_ VGND VGND VPWR VPWR _13180_ sky130_fd_sc_hd__nor2_2
X_29369_ clknet_leaf_205_clk _01104_ VGND VGND VPWR VPWR datamem.data_ram\[60\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19122_ rvcpu.dp.plde.ImmExtE\[14\] rvcpu.dp.plde.PCE\[14\] VGND VGND VPWR VPWR _06441_
+ sky130_fd_sc_hd__nand2_1
X_31400_ clknet_leaf_46_clk _03103_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCE\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16334_ net4110 _14432_ _14525_ VGND VGND VPWR VPWR _14531_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32380_ clknet_leaf_162_clk _03802_ VGND VGND VPWR VPWR datamem.data_ram\[2\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19053_ rvcpu.dp.plde.ImmExtE\[5\] rvcpu.dp.plde.PCE\[5\] VGND VGND VPWR VPWR _06381_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31331_ clknet_leaf_15_clk _03034_ VGND VGND VPWR VPWR rvcpu.dp.plde.RdE\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_644 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16265_ _14494_ VGND VGND VPWR VPWR _01903_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_11_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15216_ _13739_ _13743_ _13753_ _13757_ VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__o211a_1
X_18004_ _05370_ _05373_ VGND VGND VPWR VPWR _05374_ sky130_fd_sc_hd__nand2_1
X_31262_ clknet_leaf_19_clk _02965_ VGND VGND VPWR VPWR rvcpu.dp.plfd.InstrD\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16196_ _13222_ VGND VGND VPWR VPWR _14449_ sky130_fd_sc_hd__buf_4
Xclkbuf_1_0__f__10110_ clknet_0__10110_ VGND VGND VPWR VPWR clknet_1_0__leaf__10110_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_168_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30213_ net567 _01948_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[7\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_15147_ _13375_ _13689_ _13690_ VGND VGND VPWR VPWR _13691_ sky130_fd_sc_hd__a21oi_1
X_31193_ clknet_leaf_51_clk _02896_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCPlus4D\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30144_ net506 _01879_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[0\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_207_5462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15078_ _13410_ _13420_ _13623_ _13466_ VGND VGND VPWR VPWR _13624_ sky130_fd_sc_hd__a2bb2o_1
X_19955_ datamem.data_ram\[56\]\[18\] _06646_ _06765_ datamem.data_ram\[60\]\[18\]
+ _07248_ VGND VGND VPWR VPWR _07249_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_207_5473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18906_ _06136_ _05988_ VGND VGND VPWR VPWR _06247_ sky130_fd_sc_hd__nor2_1
X_30075_ net437 _01810_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[12\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_19886_ datamem.data_ram\[26\]\[17\] _06613_ _07077_ datamem.data_ram\[27\]\[17\]
+ _07180_ VGND VGND VPWR VPWR _07181_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_203_5359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_4330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_5263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_4341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_5274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18837_ _05239_ _06166_ _06167_ _06182_ VGND VGND VPWR VPWR rvcpu.ALUResultE\[18\]
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_222_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18768_ _05749_ _06111_ _06115_ _05702_ _06117_ VGND VGND VPWR VPWR _06118_ sky130_fd_sc_hd__a221o_1
XFILLER_0_222_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_214_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17719_ _05134_ VGND VGND VPWR VPWR _01181_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_222_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18699_ _06037_ _06038_ _06042_ _06052_ VGND VGND VPWR VPWR rvcpu.ALUResultE\[10\]
+ sky130_fd_sc_hd__a211o_2
X_30977_ clknet_leaf_166_clk _02712_ VGND VGND VPWR VPWR datamem.data_ram\[39\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_203_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20730_ datamem.data_ram\[24\]\[6\] datamem.data_ram\[25\]\[6\] datamem.data_ram\[26\]\[6\]
+ datamem.data_ram\[27\]\[6\] _07836_ _07822_ VGND VGND VPWR VPWR _08020_ sky130_fd_sc_hd__mux4_1
X_32716_ clknet_leaf_253_clk _04138_ VGND VGND VPWR VPWR datamem.data_ram\[17\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_158_4281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_4292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32647_ clknet_leaf_157_clk _04069_ VGND VGND VPWR VPWR datamem.data_ram\[1\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20661_ datamem.data_ram\[62\]\[29\] _06627_ _06805_ datamem.data_ram\[60\]\[29\]
+ VGND VGND VPWR VPWR _07952_ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22400_ rvcpu.dp.rf.reg_file_arr\[28\]\[5\] rvcpu.dp.rf.reg_file_arr\[30\]\[5\] rvcpu.dp.rf.reg_file_arr\[29\]\[5\]
+ rvcpu.dp.rf.reg_file_arr\[31\]\[5\] _09443_ _09453_ VGND VGND VPWR VPWR _09561_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_163_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_4189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23380_ clknet_1_1__leaf__10130_ VGND VGND VPWR VPWR _10140_ sky130_fd_sc_hd__buf_1
X_20592_ _07839_ _07880_ _07882_ _07867_ VGND VGND VPWR VPWR _07883_ sky130_fd_sc_hd__a211o_1
XFILLER_0_34_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32578_ clknet_leaf_265_clk _04000_ VGND VGND VPWR VPWR datamem.data_ram\[21\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22331_ _09398_ VGND VGND VPWR VPWR _09495_ sky130_fd_sc_hd__clkbuf_4
X_31529_ clknet_leaf_28_clk net1199 VGND VGND VPWR VPWR rvcpu.dp.plem.PCPlus4M\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_1290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_4506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25050_ _10741_ _10630_ _10705_ VGND VGND VPWR VPWR _10752_ sky130_fd_sc_hd__a21oi_4
X_22262_ _09415_ _09420_ _09427_ VGND VGND VPWR VPWR _09428_ sky130_fd_sc_hd__a21o_1
XFILLER_0_143_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23813__396 clknet_1_0__leaf__10207_ VGND VGND VPWR VPWR net522 sky130_fd_sc_hd__inv_2
XFILLER_0_131_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24001_ clknet_1_0__leaf__10224_ VGND VGND VPWR VPWR _10241_ sky130_fd_sc_hd__buf_1
X_21213_ _08487_ _07226_ _08490_ VGND VGND VPWR VPWR _04423_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_131_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22193_ _09256_ net3751 _09362_ VGND VGND VPWR VPWR _09369_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_113_3196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__10239_ clknet_0__10239_ VGND VGND VPWR VPWR clknet_1_0__leaf__10239_
+ sky130_fd_sc_hd__clkbuf_16
X_21144_ datamem.data_ram\[57\]\[23\] _06654_ _08432_ _07874_ _06598_ VGND VGND VPWR
+ VPWR _08433_ sky130_fd_sc_hd__o221a_1
XFILLER_0_228_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23054__754 clknet_1_1__leaf__10090_ VGND VGND VPWR VPWR net880 sky130_fd_sc_hd__inv_2
X_25952_ rvcpu.dp.plfd.PCD\[30\] _11155_ VGND VGND VPWR VPWR _11298_ sky130_fd_sc_hd__or2_1
X_21075_ datamem.data_ram\[45\]\[7\] _07831_ _08363_ _05371_ VGND VGND VPWR VPWR _08364_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28740_ _12737_ net3353 net41 VGND VGND VPWR VPWR _12870_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_126_3513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_3524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_1209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20026_ _06752_ _07314_ _07319_ _06860_ VGND VGND VPWR VPWR _07320_ sky130_fd_sc_hd__a31o_1
X_24903_ _10668_ _10640_ _10611_ VGND VGND VPWR VPWR _10669_ sky130_fd_sc_hd__a21oi_4
X_28671_ _12833_ VGND VGND VPWR VPWR _04127_ sky130_fd_sc_hd__clkbuf_1
X_25883_ _11146_ VGND VGND VPWR VPWR _11258_ sky130_fd_sc_hd__buf_2
XFILLER_0_225_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24834_ _10439_ net3023 _10631_ VGND VGND VPWR VPWR _10632_ sky130_fd_sc_hd__mux2_1
X_27622_ _12087_ net3952 net80 VGND VGND VPWR VPWR _12246_ sky130_fd_sc_hd__mux2_1
X_23169__841 clknet_1_0__leaf__10110_ VGND VGND VPWR VPWR net967 sky130_fd_sc_hd__inv_2
XFILLER_0_197_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_87_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27553_ _12209_ VGND VGND VPWR VPWR _03633_ sky130_fd_sc_hd__clkbuf_1
X_24765_ _10592_ VGND VGND VPWR VPWR _02462_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_201_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21977_ rvcpu.dp.rf.reg_file_arr\[8\]\[31\] rvcpu.dp.rf.reg_file_arr\[10\]\[31\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[31\] rvcpu.dp.rf.reg_file_arr\[11\]\[31\] rvcpu.dp.plfd.InstrD\[16\]
+ _08524_ VGND VGND VPWR VPWR _09208_ sky130_fd_sc_hd__mux4_1
XFILLER_0_150_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20928_ datamem.data_ram\[38\]\[22\] datamem.data_ram\[39\]\[22\] _07827_ VGND VGND
+ VPWR VPWR _08218_ sky130_fd_sc_hd__mux2_1
X_27484_ _12172_ VGND VGND VPWR VPWR _03601_ sky130_fd_sc_hd__clkbuf_1
X_24696_ _10555_ VGND VGND VPWR VPWR _02430_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0__10104_ _10104_ VGND VGND VPWR VPWR clknet_0__10104_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_16_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26435_ net1869 _11542_ _11567_ _11534_ VGND VGND VPWR VPWR _03157_ sky130_fd_sc_hd__o211a_1
XFILLER_0_194_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29223_ _10075_ _13123_ VGND VGND VPWR VPWR _13131_ sky130_fd_sc_hd__and2_1
XFILLER_0_127_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23647_ _09291_ net2376 _10182_ VGND VGND VPWR VPWR _10190_ sky130_fd_sc_hd__mux2_1
X_20859_ _07635_ datamem.data_ram\[13\]\[14\] _07833_ datamem.data_ram\[12\]\[14\]
+ _07863_ VGND VGND VPWR VPWR _08149_ sky130_fd_sc_hd__a221o_1
XFILLER_0_154_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_840 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29154_ _13093_ VGND VGND VPWR VPWR _04350_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_46_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26366_ _11104_ VGND VGND VPWR VPWR _11517_ sky130_fd_sc_hd__buf_2
XFILLER_0_119_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28105_ _12517_ VGND VGND VPWR VPWR _03877_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25317_ _10903_ VGND VGND VPWR VPWR _02703_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29085_ _12766_ net2032 _13049_ VGND VGND VPWR VPWR _13057_ sky130_fd_sc_hd__mux2_1
X_22529_ rvcpu.dp.rf.reg_file_arr\[12\]\[11\] rvcpu.dp.rf.reg_file_arr\[13\]\[11\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[11\] rvcpu.dp.rf.reg_file_arr\[15\]\[11\] _09478_
+ _09479_ VGND VGND VPWR VPWR _09684_ sky130_fd_sc_hd__mux4_2
X_26297_ _11481_ VGND VGND VPWR VPWR _03105_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_161_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28036_ _12480_ VGND VGND VPWR VPWR _03845_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16050_ _14365_ VGND VGND VPWR VPWR _01997_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_59_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25248_ _10737_ net2763 _10857_ VGND VGND VPWR VPWR _10864_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15001_ _13545_ _13547_ _13548_ VGND VGND VPWR VPWR _13549_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_55_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25179_ _09329_ VGND VGND VPWR VPWR _10826_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_55_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24007__540 clknet_1_1__leaf__10241_ VGND VGND VPWR VPWR net666 sky130_fd_sc_hd__inv_2
XFILLER_0_209_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29987_ net357 _01722_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[14\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23487__134 clknet_1_0__leaf__10159_ VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__inv_2
X_19740_ _07018_ _07022_ _07027_ _07034_ VGND VGND VPWR VPWR _07035_ sky130_fd_sc_hd__a31o_1
X_28938_ _12764_ net2276 _12968_ VGND VGND VPWR VPWR _12975_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16952_ _04727_ VGND VGND VPWR VPWR _01565_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15903_ net1982 _13213_ _14286_ VGND VGND VPWR VPWR _14287_ sky130_fd_sc_hd__mux2_1
X_19671_ _06810_ VGND VGND VPWR VPWR _06967_ sky130_fd_sc_hd__buf_6
X_16883_ net2514 _14434_ _04684_ VGND VGND VPWR VPWR _04691_ sky130_fd_sc_hd__mux2_1
X_28869_ _12938_ VGND VGND VPWR VPWR _04220_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_218_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18622_ _05346_ _05405_ _05886_ VGND VGND VPWR VPWR _05979_ sky130_fd_sc_hd__a21oi_1
X_30900_ clknet_leaf_150_clk _02635_ VGND VGND VPWR VPWR datamem.data_ram\[41\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15834_ net2055 _13217_ _14247_ VGND VGND VPWR VPWR _14249_ sky130_fd_sc_hd__mux2_1
X_31880_ clknet_leaf_111_clk _03334_ VGND VGND VPWR VPWR datamem.data_ram\[57\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_204_Left_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18553_ _05368_ _05401_ _05886_ VGND VGND VPWR VPWR _05913_ sky130_fd_sc_hd__a21o_1
X_30831_ clknet_leaf_151_clk _02566_ VGND VGND VPWR VPWR datamem.data_ram\[44\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_194_5160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15765_ _14154_ net4009 _14210_ VGND VGND VPWR VPWR _14212_ sky130_fd_sc_hd__mux2_1
X_17504_ _05020_ VGND VGND VPWR VPWR _01290_ sky130_fd_sc_hd__clkbuf_1
X_14716_ _13271_ VGND VGND VPWR VPWR _13272_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_190_5046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30762_ clknet_leaf_136_clk _02497_ VGND VGND VPWR VPWR datamem.data_ram\[47\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_18484_ _05841_ _05845_ _05692_ VGND VGND VPWR VPWR _05846_ sky130_fd_sc_hd__mux2_1
X_15696_ _13237_ VGND VGND VPWR VPWR _14168_ sky130_fd_sc_hd__buf_4
XFILLER_0_59_369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_460 _08634_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_190_5057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_471 _08971_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32501_ clknet_leaf_249_clk _03923_ VGND VGND VPWR VPWR datamem.data_ram\[25\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14647_ _13219_ VGND VGND VPWR VPWR _13220_ sky130_fd_sc_hd__clkbuf_8
XANTENNA_482 _09317_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17435_ _14149_ net4283 _04974_ VGND VGND VPWR VPWR _04984_ sky130_fd_sc_hd__mux2_1
X_30693_ clknet_leaf_156_clk _02428_ VGND VGND VPWR VPWR datamem.data_ram\[4\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_493 _09750_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_18 _06612_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32432_ clknet_leaf_274_clk _03854_ VGND VGND VPWR VPWR datamem.data_ram\[28\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17366_ _04947_ VGND VGND VPWR VPWR _01355_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_29 _06634_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19105_ _06426_ VGND VGND VPWR VPWR rvcpu.dp.lAuiPCE\[11\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16317_ _14521_ VGND VGND VPWR VPWR _01878_ sky130_fd_sc_hd__clkbuf_1
X_32363_ clknet_leaf_93_clk _03785_ VGND VGND VPWR VPWR datamem.data_ram\[2\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17297_ net4430 _13206_ _04902_ VGND VGND VPWR VPWR _04911_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_213_Left_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19036_ _06366_ VGND VGND VPWR VPWR rvcpu.dp.lAuiPCE\[2\] sky130_fd_sc_hd__clkbuf_1
X_31314_ clknet_leaf_44_clk _03017_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCPlus4E\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_16248_ _13274_ VGND VGND VPWR VPWR _14484_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_209_5502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23339__977 clknet_1_1__leaf__10136_ VGND VGND VPWR VPWR net1103 sky130_fd_sc_hd__inv_2
X_32294_ clknet_leaf_215_clk _03716_ VGND VGND VPWR VPWR datamem.data_ram\[32\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_209_5513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31245_ clknet_leaf_21_clk _02948_ VGND VGND VPWR VPWR rvcpu.dp.plfd.InstrD\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16179_ _14437_ VGND VGND VPWR VPWR _01940_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31176_ clknet_leaf_238_clk _02879_ VGND VGND VPWR VPWR datamem.data_ram\[5\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30127_ net489 _01862_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[10\]\[18\] sky130_fd_sc_hd__dfxtp_1
Xhold2905 datamem.data_ram\[24\]\[11\] VGND VGND VPWR VPWR net4055 sky130_fd_sc_hd__dlygate4sd3_1
X_19938_ datamem.data_ram\[39\]\[18\] _06760_ _06782_ datamem.data_ram\[33\]\[18\]
+ _06769_ VGND VGND VPWR VPWR _07232_ sky130_fd_sc_hd__o221a_1
Xhold2916 rvcpu.dp.rf.reg_file_arr\[29\]\[17\] VGND VGND VPWR VPWR net4066 sky130_fd_sc_hd__dlygate4sd3_1
X_23118__795 clknet_1_0__leaf__10105_ VGND VGND VPWR VPWR net921 sky130_fd_sc_hd__inv_2
Xhold2927 datamem.data_ram\[57\]\[14\] VGND VGND VPWR VPWR net4077 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2938 rvcpu.dp.rf.reg_file_arr\[23\]\[10\] VGND VGND VPWR VPWR net4088 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2949 datamem.data_ram\[56\]\[28\] VGND VGND VPWR VPWR net4099 sky130_fd_sc_hd__dlygate4sd3_1
X_30058_ net420 _01793_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[12\]\[13\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_222_Left_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19869_ datamem.data_ram\[12\]\[1\] _07123_ _07160_ _07163_ VGND VGND VPWR VPWR _07164_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_223_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21900_ rvcpu.dp.rf.reg_file_arr\[0\]\[27\] rvcpu.dp.rf.reg_file_arr\[1\]\[27\] rvcpu.dp.rf.reg_file_arr\[2\]\[27\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[27\] _08810_ _08811_ VGND VGND VPWR VPWR _09135_
+ sky130_fd_sc_hd__mux4_1
X_22880_ _09433_ _10015_ _09789_ VGND VGND VPWR VPWR _10016_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_121_3410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21831_ rvcpu.dp.rf.reg_file_arr\[4\]\[23\] rvcpu.dp.rf.reg_file_arr\[5\]\[23\] rvcpu.dp.rf.reg_file_arr\[6\]\[23\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[23\] _08839_ _08840_ VGND VGND VPWR VPWR _09070_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_214_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_223_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_156_4229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24550_ _10472_ net3044 net60 VGND VGND VPWR VPWR _10473_ sky130_fd_sc_hd__mux2_1
X_21762_ rvcpu.dp.rf.reg_file_arr\[16\]\[20\] rvcpu.dp.rf.reg_file_arr\[17\]\[20\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[20\] rvcpu.dp.rf.reg_file_arr\[19\]\[20\] _08799_
+ _08800_ VGND VGND VPWR VPWR _09004_ sky130_fd_sc_hd__mux4_1
XFILLER_0_148_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20713_ datamem.data_ram\[16\]\[5\] _06990_ _06976_ datamem.data_ram\[20\]\[5\] VGND
+ VGND VPWR VPWR _08004_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24481_ _09298_ datamem.data_ram\[52\]\[24\] _10430_ VGND VGND VPWR VPWR _10431_
+ sky130_fd_sc_hd__mux2_1
X_21693_ _08515_ _08938_ VGND VGND VPWR VPWR _08939_ sky130_fd_sc_hd__nor2_1
XFILLER_0_188_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26220_ net1176 _11436_ _11444_ VGND VGND VPWR VPWR _11448_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_3350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20644_ datamem.data_ram\[23\]\[29\] _07020_ _07931_ _07934_ VGND VGND VPWR VPWR
+ _07935_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_119_3361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26151_ net1621 _11408_ VGND VGND VPWR VPWR _11412_ sky130_fd_sc_hd__and2_1
X_20575_ _06641_ VGND VGND VPWR VPWR _07866_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_115_3247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25102_ _10070_ _10779_ _10781_ net1341 VGND VGND VPWR VPWR _02609_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_115_3258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22314_ _09383_ VGND VGND VPWR VPWR _09479_ sky130_fd_sc_hd__buf_6
X_26082_ _11373_ VGND VGND VPWR VPWR _02997_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_41_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_186_4948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_225_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25033_ _10465_ net3231 net90 VGND VGND VPWR VPWR _10743_ sky130_fd_sc_hd__mux2_1
X_29910_ net280 _01645_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[16\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_186_4959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22245_ rvcpu.dp.plfd.InstrD\[23\] VGND VGND VPWR VPWR _09411_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29841_ net219 _01576_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[18\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22176_ _09359_ VGND VGND VPWR VPWR _01106_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_218_515 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_195_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21127_ datamem.data_ram\[36\]\[23\] datamem.data_ram\[37\]\[23\] _07826_ VGND VGND
+ VPWR VPWR _08416_ sky130_fd_sc_hd__mux2_1
X_29772_ net1118 _01507_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[20\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_26984_ _11876_ VGND VGND VPWR VPWR _03397_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28723_ _12754_ net3167 _12859_ VGND VGND VPWR VPWR _12861_ sky130_fd_sc_hd__mux2_1
X_25935_ _11157_ VGND VGND VPWR VPWR _11288_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_145_3966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21058_ _07862_ _08346_ VGND VGND VPWR VPWR _08347_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_145_3977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20009_ datamem.data_ram\[62\]\[2\] _06951_ _06769_ _07302_ VGND VGND VPWR VPWR _07303_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_199_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25866_ rvcpu.dp.plfd.PCPlus4D\[29\] _11244_ _08598_ VGND VGND VPWR VPWR _11245_
+ sky130_fd_sc_hd__mux2_1
X_28654_ _12824_ VGND VGND VPWR VPWR _04119_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27605_ _12149_ net2689 net81 VGND VGND VPWR VPWR _12237_ sky130_fd_sc_hd__mux2_1
X_24817_ _10622_ VGND VGND VPWR VPWR _02484_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_214_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25797_ _11188_ _11189_ _11149_ VGND VGND VPWR VPWR _11190_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_201_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28585_ _12787_ VGND VGND VPWR VPWR _04087_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_198_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_198_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15550_ _13823_ _13435_ VGND VGND VPWR VPWR _14074_ sky130_fd_sc_hd__nand2_1
X_27536_ _12200_ VGND VGND VPWR VPWR _03625_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_48_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24037__566 clknet_1_0__leaf__10245_ VGND VGND VPWR VPWR net692 sky130_fd_sc_hd__inv_2
XFILLER_0_96_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24748_ _10583_ VGND VGND VPWR VPWR _02454_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15481_ _13599_ _13391_ _13510_ _14008_ _14009_ VGND VGND VPWR VPWR _14010_ sky130_fd_sc_hd__o311a_1
X_27467_ _12087_ net2986 net83 VGND VGND VPWR VPWR _12163_ sky130_fd_sc_hd__mux2_1
XFILLER_0_194_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_189_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24679_ _10546_ VGND VGND VPWR VPWR _02422_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_13_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29206_ _10042_ _10947_ VGND VGND VPWR VPWR _13121_ sky130_fd_sc_hd__or2_1
X_17220_ _14139_ net4362 _04865_ VGND VGND VPWR VPWR _04870_ sky130_fd_sc_hd__mux2_1
X_22965__674 clknet_1_0__leaf__10081_ VGND VGND VPWR VPWR net800 sky130_fd_sc_hd__inv_2
X_26418_ _11545_ rvcpu.ALUResultE\[12\] VGND VGND VPWR VPWR _11556_ sky130_fd_sc_hd__and2_1
XFILLER_0_181_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27398_ _12085_ net2301 net85 VGND VGND VPWR VPWR _12119_ sky130_fd_sc_hd__mux2_1
XFILLER_0_182_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17151_ _04833_ VGND VGND VPWR VPWR _01464_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26349_ _10782_ _11507_ _11508_ net1345 VGND VGND VPWR VPWR _03130_ sky130_fd_sc_hd__a22o_1
X_29137_ _13084_ VGND VGND VPWR VPWR _04342_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16102_ net4383 _13204_ _14385_ VGND VGND VPWR VPWR _14393_ sky130_fd_sc_hd__mux2_1
X_29068_ _09290_ net2011 _13040_ VGND VGND VPWR VPWR _13048_ sky130_fd_sc_hd__mux2_1
X_17082_ _14137_ net3943 _04793_ VGND VGND VPWR VPWR _04797_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16033_ _14356_ VGND VGND VPWR VPWR _02005_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28019_ _12471_ VGND VGND VPWR VPWR _03837_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_161_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31030_ clknet_leaf_102_clk _02765_ VGND VGND VPWR VPWR datamem.data_ram\[12\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_209_526 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17984_ _05349_ _05353_ VGND VGND VPWR VPWR _05354_ sky130_fd_sc_hd__and2_1
XFILLER_0_100_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_202_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_200_5307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19723_ datamem.data_ram\[9\]\[25\] _06659_ VGND VGND VPWR VPWR _07018_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_196_5200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16935_ net2404 _14486_ _04683_ VGND VGND VPWR VPWR _04718_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_196_5211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32981_ clknet_leaf_268_clk _04403_ VGND VGND VPWR VPWR datamem.data_ram\[63\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_221_5790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31932_ clknet_leaf_123_clk _03354_ VGND VGND VPWR VPWR datamem.data_ram\[60\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_19654_ rvcpu.dp.plem.ALUResultM\[2\] _06922_ VGND VGND VPWR VPWR _06950_ sky130_fd_sc_hd__nor2_8
X_16866_ _04681_ VGND VGND VPWR VPWR _01605_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_192_5108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18605_ _05960_ _05962_ _05696_ VGND VGND VPWR VPWR _05963_ sky130_fd_sc_hd__mux2_1
X_15817_ net2005 _13190_ _14236_ VGND VGND VPWR VPWR _14240_ sky130_fd_sc_hd__mux2_1
X_31863_ clknet_leaf_124_clk _03317_ VGND VGND VPWR VPWR datamem.data_ram\[63\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_19585_ datamem.data_ram\[44\]\[8\] _06618_ _06781_ datamem.data_ram\[41\]\[8\] VGND
+ VGND VPWR VPWR _06881_ sky130_fd_sc_hd__o22a_1
XFILLER_0_177_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16797_ net2111 _14484_ _04611_ VGND VGND VPWR VPWR _04645_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18536_ _05606_ net102 _05604_ _05596_ _05684_ _05689_ VGND VGND VPWR VPWR _05897_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_133_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30814_ clknet_leaf_280_clk _02549_ VGND VGND VPWR VPWR datamem.data_ram\[45\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15748_ _14137_ net4351 _14199_ VGND VGND VPWR VPWR _14203_ sky130_fd_sc_hd__mux2_1
X_31794_ clknet_leaf_236_clk _03248_ VGND VGND VPWR VPWR datamem.data_ram\[2\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_201_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_103 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18467_ _05824_ _05829_ _05370_ VGND VGND VPWR VPWR _05830_ sky130_fd_sc_hd__mux2_1
X_30745_ clknet_leaf_195_clk _02480_ VGND VGND VPWR VPWR datamem.data_ram\[48\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_290 _13322_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15679_ _14156_ net3588 _14152_ VGND VGND VPWR VPWR _14157_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_4115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17418_ _04975_ VGND VGND VPWR VPWR _01331_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_151_4126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18398_ _05760_ _05761_ _05668_ VGND VGND VPWR VPWR _05762_ sky130_fd_sc_hd__mux2_1
X_30676_ clknet_leaf_190_clk _02411_ VGND VGND VPWR VPWR datamem.data_ram\[50\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32415_ clknet_leaf_184_clk _03837_ VGND VGND VPWR VPWR datamem.data_ram\[28\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_17349_ _14127_ net3598 _04938_ VGND VGND VPWR VPWR _04939_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload210 clknet_leaf_204_clk VGND VGND VPWR VPWR clkload210/Y sky130_fd_sc_hd__clkinvlp_4
X_32346_ clknet_leaf_81_clk _03768_ VGND VGND VPWR VPWR datamem.data_ram\[30\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20360_ datamem.data_ram\[6\]\[28\] _06763_ _06766_ datamem.data_ram\[4\]\[28\] VGND
+ VGND VPWR VPWR _07652_ sky130_fd_sc_hd__o22a_1
Xclkload221 clknet_leaf_280_clk VGND VGND VPWR VPWR clkload221/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_0_67_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload232 clknet_leaf_111_clk VGND VGND VPWR VPWR clkload232/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_31_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload243 clknet_leaf_133_clk VGND VGND VPWR VPWR clkload243/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_130_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19019_ rvcpu.dp.plde.ImmExtE\[0\] rvcpu.dp.plde.PCE\[0\] VGND VGND VPWR VPWR _06352_
+ sky130_fd_sc_hd__nand2_1
Xclkload254 clknet_leaf_192_clk VGND VGND VPWR VPWR clkload254/Y sky130_fd_sc_hd__inv_6
XFILLER_0_114_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23272__917 clknet_1_0__leaf__10129_ VGND VGND VPWR VPWR net1043 sky130_fd_sc_hd__inv_2
Xclkload265 clknet_leaf_121_clk VGND VGND VPWR VPWR clkload265/Y sky130_fd_sc_hd__inv_6
X_20291_ datamem.data_ram\[17\]\[19\] _06659_ _07580_ _07583_ VGND VGND VPWR VPWR
+ _07584_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_228_5966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32277_ clknet_leaf_167_clk _03699_ VGND VGND VPWR VPWR datamem.data_ram\[33\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload276 clknet_leaf_138_clk VGND VGND VPWR VPWR clkload276/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_110_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_228_5977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload287 clknet_1_0__leaf__10241_ VGND VGND VPWR VPWR clkload287/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_149_4066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22030_ rvcpu.dp.plem.WriteDataM\[22\] _09220_ VGND VGND VPWR VPWR _09254_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload298 clknet_1_0__leaf__10208_ VGND VGND VPWR VPWR clkload298/Y sky130_fd_sc_hd__clkinvlp_4
X_31228_ clknet_leaf_42_clk _02931_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCD\[17\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_149_4077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_181_4834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_181_4845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31159_ clknet_leaf_68_clk rvcpu.ALUResultE\[18\] VGND VGND VPWR VPWR rvcpu.dp.plem.ALUResultM\[18\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2702 datamem.data_ram\[40\]\[20\] VGND VGND VPWR VPWR net3852 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2713 datamem.data_ram\[39\]\[12\] VGND VGND VPWR VPWR net3863 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2724 datamem.data_ram\[11\]\[18\] VGND VGND VPWR VPWR net3874 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_71_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2735 rvcpu.dp.rf.reg_file_arr\[23\]\[15\] VGND VGND VPWR VPWR net3885 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2746 rvcpu.dp.rf.reg_file_arr\[21\]\[8\] VGND VGND VPWR VPWR net3896 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2757 datamem.data_ram\[61\]\[20\] VGND VGND VPWR VPWR net3907 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2768 rvcpu.dp.rf.reg_file_arr\[21\]\[6\] VGND VGND VPWR VPWR net3918 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2779 datamem.data_ram\[48\]\[21\] VGND VGND VPWR VPWR net3929 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25720_ _10811_ net3711 _11133_ VGND VGND VPWR VPWR _11134_ sky130_fd_sc_hd__mux2_1
X_22932_ rvcpu.dp.plem.WriteDataM\[3\] VGND VGND VPWR VPWR _10063_ sky130_fd_sc_hd__buf_4
XFILLER_0_138_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_108_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_1231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25651_ _10058_ _11094_ _11095_ net1415 VGND VGND VPWR VPWR _02845_ sky130_fd_sc_hd__a22o_1
XFILLER_0_223_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_3852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22863_ rvcpu.dp.rf.reg_file_arr\[8\]\[29\] rvcpu.dp.rf.reg_file_arr\[10\]\[29\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[29\] rvcpu.dp.rf.reg_file_arr\[11\]\[29\] _09483_
+ _09656_ VGND VGND VPWR VPWR _10000_ sky130_fd_sc_hd__mux4_1
XFILLER_0_155_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_3863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_179_4785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_179_4796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_119_Left_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24602_ _10503_ VGND VGND VPWR VPWR _02388_ sky130_fd_sc_hd__clkbuf_1
X_28370_ _12660_ VGND VGND VPWR VPWR _03999_ sky130_fd_sc_hd__clkbuf_1
X_21814_ _08695_ _09053_ VGND VGND VPWR VPWR _09054_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_80_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25582_ _07019_ _10946_ _10044_ VGND VGND VPWR VPWR _11052_ sky130_fd_sc_hd__or3_1
XFILLER_0_151_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire62 _09341_ VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__buf_4
X_22794_ _09461_ _09932_ _09934_ _09474_ VGND VGND VPWR VPWR _09935_ sky130_fd_sc_hd__o211a_1
XFILLER_0_38_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27321_ _12075_ VGND VGND VPWR VPWR _12076_ sky130_fd_sc_hd__clkbuf_2
X_24533_ _10396_ net4396 _10456_ VGND VGND VPWR VPWR _10462_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21745_ rvcpu.dp.rf.reg_file_arr\[20\]\[19\] rvcpu.dp.rf.reg_file_arr\[21\]\[19\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[19\] rvcpu.dp.rf.reg_file_arr\[23\]\[19\] _08799_
+ _08518_ VGND VGND VPWR VPWR _08988_ sky130_fd_sc_hd__mux4_2
XFILLER_0_136_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27252_ _11980_ _12031_ VGND VGND VPWR VPWR _12040_ sky130_fd_sc_hd__and2_1
XFILLER_0_171_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24464_ _09298_ net3157 _10421_ VGND VGND VPWR VPWR _10422_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21676_ _08742_ _08922_ VGND VGND VPWR VPWR _08923_ sky130_fd_sc_hd__or2_1
X_26203_ _02995_ _02996_ _11439_ VGND VGND VPWR VPWR _11440_ sky130_fd_sc_hd__or3_1
XFILLER_0_164_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27183_ _11991_ net1431 _11995_ _11999_ VGND VGND VPWR VPWR _03473_ sky130_fd_sc_hd__a31o_1
XFILLER_0_190_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20627_ _07177_ _07909_ _07917_ _07154_ _06602_ VGND VGND VPWR VPWR _07918_ sky130_fd_sc_hd__o221a_1
XFILLER_0_184_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24395_ _09267_ net3738 _10376_ VGND VGND VPWR VPWR _10377_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_129_Right_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26134_ net1653 _11397_ VGND VGND VPWR VPWR _11403_ sky130_fd_sc_hd__and2_1
XFILLER_0_117_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20558_ _07835_ VGND VGND VPWR VPWR _07849_ sky130_fd_sc_hd__clkbuf_8
X_23670__267 clknet_1_0__leaf__10193_ VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__inv_2
XFILLER_0_34_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23438__89 clknet_1_1__leaf__10155_ VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_128_Left_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_225_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26065_ _08622_ VGND VGND VPWR VPWR _11362_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_131_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_225_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20489_ _06596_ _07747_ _07758_ _07780_ VGND VGND VPWR VPWR _07781_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_14_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25016_ _09278_ VGND VGND VPWR VPWR _10731_ sky130_fd_sc_hd__clkbuf_2
X_22228_ _08595_ VGND VGND VPWR VPWR _09394_ sky130_fd_sc_hd__buf_4
XFILLER_0_219_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29824_ net202 _01559_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[1\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_22159_ _09349_ VGND VGND VPWR VPWR _01099_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_219_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29755_ net1101 _01490_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[21\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14981_ _13528_ _13473_ _13463_ VGND VGND VPWR VPWR _13529_ sky130_fd_sc_hd__o21ai_1
X_26967_ _11863_ net1555 _11865_ _11867_ VGND VGND VPWR VPWR _03389_ sky130_fd_sc_hd__a31o_1
XFILLER_0_156_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_1115 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16720_ _04604_ VGND VGND VPWR VPWR _01682_ sky130_fd_sc_hd__clkbuf_1
X_28706_ _12690_ net3206 _12850_ VGND VGND VPWR VPWR _12852_ sky130_fd_sc_hd__mux2_1
X_25918_ net1904 _11275_ _11273_ _11278_ VGND VGND VPWR VPWR _02929_ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29686_ net1032 _01421_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[23\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_26898_ _10297_ _10921_ _10922_ VGND VGND VPWR VPWR _11823_ sky130_fd_sc_hd__and3_2
XFILLER_0_89_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_137_Left_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_198_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28637_ _12815_ VGND VGND VPWR VPWR _04111_ sky130_fd_sc_hd__clkbuf_1
X_16651_ _14183_ net3180 _04562_ VGND VGND VPWR VPWR _04568_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25849_ rvcpu.dp.pcreg.q\[26\] _11226_ VGND VGND VPWR VPWR _11231_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_18_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_639 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15602_ net2989 _13229_ _14103_ VGND VGND VPWR VPWR _14109_ sky130_fd_sc_hd__mux2_1
X_19370_ rvcpu.dp.plem.ALUResultM\[2\] VGND VGND VPWR VPWR _06666_ sky130_fd_sc_hd__clkbuf_16
X_28568_ _12778_ VGND VGND VPWR VPWR _04079_ sky130_fd_sc_hd__clkbuf_1
X_16582_ _14183_ net3243 _04525_ VGND VGND VPWR VPWR _04531_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18321_ _05382_ _05662_ VGND VGND VPWR VPWR _05686_ sky130_fd_sc_hd__nand2_1
X_15533_ _13682_ _13665_ _13348_ _13597_ VGND VGND VPWR VPWR _14059_ sky130_fd_sc_hd__a31o_1
Xclkbuf_5_21__f_clk clknet_2_2_0_clk VGND VGND VPWR VPWR clknet_5_21__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_27519_ _12191_ VGND VGND VPWR VPWR _03617_ sky130_fd_sc_hd__clkbuf_1
X_28499_ _09266_ VGND VGND VPWR VPWR _12734_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_56_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15464_ _13528_ _13435_ VGND VGND VPWR VPWR _13994_ sky130_fd_sc_hd__nor2_1
X_18252_ _05488_ _05497_ _05504_ _05512_ VGND VGND VPWR VPWR _05617_ sky130_fd_sc_hd__or4_1
X_30530_ clknet_leaf_268_clk _02265_ VGND VGND VPWR VPWR datamem.data_ram\[56\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17203_ _04860_ VGND VGND VPWR VPWR _01439_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30461_ net139 _02196_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[19\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_15395_ _13327_ _13926_ _13927_ _13504_ _13521_ VGND VGND VPWR VPWR _13928_ sky130_fd_sc_hd__a221o_1
X_18183_ _05545_ _05546_ VGND VGND VPWR VPWR _05548_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_146_Left_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32200_ clknet_leaf_199_clk _03622_ VGND VGND VPWR VPWR datamem.data_ram\[36\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17134_ _14189_ net3518 _04815_ VGND VGND VPWR VPWR _04824_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30392_ net730 _02127_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[31\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold608 datamem.data_ram\[54\]\[7\] VGND VGND VPWR VPWR net1758 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17065_ _04787_ VGND VGND VPWR VPWR _01504_ sky130_fd_sc_hd__clkbuf_1
X_32131_ clknet_leaf_213_clk _03553_ VGND VGND VPWR VPWR datamem.data_ram\[10\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold619 datamem.data_ram\[7\]\[4\] VGND VGND VPWR VPWR net1769 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16016_ rvcpu.dp.plmw.RdW\[0\] VGND VGND VPWR VPWR _14346_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_228_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32062_ clknet_leaf_119_clk _03484_ VGND VGND VPWR VPWR datamem.data_ram\[48\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31013_ clknet_leaf_154_clk _02748_ VGND VGND VPWR VPWR datamem.data_ram\[42\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_223_5841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_223_5852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2009 rvcpu.dp.rf.reg_file_arr\[25\]\[10\] VGND VGND VPWR VPWR net3159 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17967_ _05337_ VGND VGND VPWR VPWR _05338_ sky130_fd_sc_hd__inv_2
Xhold1308 rvcpu.dp.rf.reg_file_arr\[21\]\[26\] VGND VGND VPWR VPWR net2458 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1319 rvcpu.dp.rf.reg_file_arr\[15\]\[4\] VGND VGND VPWR VPWR net2469 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19706_ datamem.data_ram\[2\]\[0\] _07000_ _06966_ datamem.data_ram\[3\]\[0\] _07001_
+ VGND VGND VPWR VPWR _07002_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_155_Left_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16918_ _04709_ VGND VGND VPWR VPWR _01581_ sky130_fd_sc_hd__clkbuf_1
X_32964_ clknet_leaf_204_clk _04386_ VGND VGND VPWR VPWR datamem.data_ram\[63\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_17898_ _05270_ VGND VGND VPWR VPWR _05271_ sky130_fd_sc_hd__buf_4
X_31915_ _04427_ net120 VGND VGND VPWR VPWR datamem.rd_data_mem\[20\] sky130_fd_sc_hd__dlxtn_1
X_19637_ _06651_ VGND VGND VPWR VPWR _06933_ sky130_fd_sc_hd__buf_6
XFILLER_0_215_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_205_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16849_ net2603 _14468_ _04670_ VGND VGND VPWR VPWR _04673_ sky130_fd_sc_hd__mux2_1
X_32895_ clknet_leaf_157_clk _04317_ VGND VGND VPWR VPWR datamem.data_ram\[10\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31846_ clknet_leaf_152_clk _03300_ VGND VGND VPWR VPWR datamem.data_ram\[8\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_19568_ datamem.data_ram\[3\]\[8\] _06863_ VGND VGND VPWR VPWR _06864_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24133__638 clknet_1_1__leaf__10261_ VGND VGND VPWR VPWR net764 sky130_fd_sc_hd__inv_2
XFILLER_0_215_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18519_ _05378_ _05726_ _05729_ _05377_ VGND VGND VPWR VPWR _05880_ sky130_fd_sc_hd__a22o_1
XFILLER_0_220_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_4660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19499_ _06774_ _06775_ _06787_ _06794_ VGND VGND VPWR VPWR _06795_ sky130_fd_sc_hd__a31o_1
XFILLER_0_8_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31777_ clknet_leaf_255_clk _03231_ VGND VGND VPWR VPWR datamem.data_ram\[6\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_174_4671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_174_4682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21530_ _08686_ _08783_ _08748_ VGND VGND VPWR VPWR _08784_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_168_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30728_ clknet_leaf_219_clk _02463_ VGND VGND VPWR VPWR datamem.data_ram\[48\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_170_4568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_164_Left_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21461_ _08572_ _08718_ VGND VGND VPWR VPWR _08719_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_170_4579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30659_ clknet_leaf_194_clk _02394_ VGND VGND VPWR VPWR datamem.data_ram\[50\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23200_ _09252_ datamem.data_ram\[5\]\[21\] _10115_ VGND VGND VPWR VPWR _10121_ sky130_fd_sc_hd__mux2_1
X_20412_ datamem.data_ram\[61\]\[12\] _06661_ _06820_ datamem.data_ram\[56\]\[12\]
+ VGND VGND VPWR VPWR _07704_ sky130_fd_sc_hd__o22a_1
X_21392_ _08565_ _08648_ _08651_ _08652_ VGND VGND VPWR VPWR _08653_ sky130_fd_sc_hd__o211a_1
XFILLER_0_226_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20343_ _06666_ VGND VGND VPWR VPWR _07635_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_4_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32329_ clknet_leaf_248_clk _03751_ VGND VGND VPWR VPWR datamem.data_ram\[31\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_222_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23062_ _10042_ _09268_ VGND VGND VPWR VPWR _10092_ sky130_fd_sc_hd__nor2_8
XTAP_TAPCELL_ROW_73_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20274_ datamem.data_ram\[32\]\[19\] _06698_ _07563_ _07566_ VGND VGND VPWR VPWR
+ _07567_ sky130_fd_sc_hd__o211a_1
XFILLER_0_80_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold3200 datamem.data_ram\[58\]\[21\] VGND VGND VPWR VPWR net4350 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22013_ _09240_ net4355 _09232_ VGND VGND VPWR VPWR _09241_ sky130_fd_sc_hd__mux2_1
Xhold3211 datamem.data_ram\[55\]\[20\] VGND VGND VPWR VPWR net4361 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_179_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold3222 datamem.data_ram\[55\]\[16\] VGND VGND VPWR VPWR net4372 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3233 rvcpu.dp.rf.reg_file_arr\[7\]\[24\] VGND VGND VPWR VPWR net4383 sky130_fd_sc_hd__dlygate4sd3_1
X_27870_ _12145_ net3299 net77 VGND VGND VPWR VPWR _12384_ sky130_fd_sc_hd__mux2_1
Xhold3244 rvcpu.dp.rf.reg_file_arr\[29\]\[16\] VGND VGND VPWR VPWR net4394 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3255 datamem.data_ram\[62\]\[16\] VGND VGND VPWR VPWR net4405 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2510 datamem.data_ram\[32\]\[27\] VGND VGND VPWR VPWR net3660 sky130_fd_sc_hd__dlygate4sd3_1
X_26821_ _11767_ net1624 _11773_ _11776_ VGND VGND VPWR VPWR _03334_ sky130_fd_sc_hd__a31o_1
Xhold3266 rvcpu.dp.rf.reg_file_arr\[7\]\[27\] VGND VGND VPWR VPWR net4416 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2521 datamem.data_ram\[8\]\[24\] VGND VGND VPWR VPWR net3671 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2532 datamem.data_ram\[11\]\[22\] VGND VGND VPWR VPWR net3682 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3277 datamem.data_ram\[52\]\[16\] VGND VGND VPWR VPWR net4427 sky130_fd_sc_hd__dlygate4sd3_1
X_23706__300 clknet_1_0__leaf__10196_ VGND VGND VPWR VPWR net426 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_142_3903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3288 datamem.data_ram\[53\]\[15\] VGND VGND VPWR VPWR net4438 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2543 datamem.data_ram\[47\]\[8\] VGND VGND VPWR VPWR net3693 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold3299 rvcpu.dp.plfd.InstrD\[11\] VGND VGND VPWR VPWR net4449 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2554 datamem.data_ram\[43\]\[17\] VGND VGND VPWR VPWR net3704 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1820 rvcpu.dp.rf.reg_file_arr\[13\]\[1\] VGND VGND VPWR VPWR net2970 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2565 datamem.data_ram\[8\]\[26\] VGND VGND VPWR VPWR net3715 sky130_fd_sc_hd__dlygate4sd3_1
X_29540_ net894 _01275_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[27\]\[7\] sky130_fd_sc_hd__dfxtp_1
Xhold1831 datamem.data_ram\[59\]\[31\] VGND VGND VPWR VPWR net2981 sky130_fd_sc_hd__dlygate4sd3_1
X_26752_ _10783_ _08356_ _11724_ VGND VGND VPWR VPWR _11734_ sky130_fd_sc_hd__mux2_1
X_23964_ _09256_ net3504 _10229_ VGND VGND VPWR VPWR _10236_ sky130_fd_sc_hd__mux2_1
Xhold2576 datamem.data_ram\[40\]\[17\] VGND VGND VPWR VPWR net3726 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1842 datamem.data_ram\[45\]\[9\] VGND VGND VPWR VPWR net2992 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2587 datamem.data_ram\[53\]\[31\] VGND VGND VPWR VPWR net3737 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2598 datamem.data_ram\[18\]\[27\] VGND VGND VPWR VPWR net3748 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1853 datamem.data_ram\[27\]\[9\] VGND VGND VPWR VPWR net3003 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1864 datamem.data_ram\[39\]\[9\] VGND VGND VPWR VPWR net3014 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22915_ _06604_ _07154_ VGND VGND VPWR VPWR _10049_ sky130_fd_sc_hd__nor2_1
X_25703_ _10811_ net3797 _11124_ VGND VGND VPWR VPWR _11125_ sky130_fd_sc_hd__mux2_1
Xhold1875 datamem.data_ram\[6\]\[28\] VGND VGND VPWR VPWR net3025 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26683_ _11683_ net1782 _11693_ _11695_ VGND VGND VPWR VPWR _03277_ sky130_fd_sc_hd__a31o_1
Xhold1886 datamem.data_ram\[26\]\[26\] VGND VGND VPWR VPWR net3036 sky130_fd_sc_hd__dlygate4sd3_1
X_29471_ net833 _01206_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[2\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_196_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23895_ clknet_1_1__leaf__10203_ VGND VGND VPWR VPWR _10223_ sky130_fd_sc_hd__buf_1
Xhold1897 rvcpu.dp.rf.reg_file_arr\[30\]\[9\] VGND VGND VPWR VPWR net3047 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28422_ _12687_ net3745 _12688_ VGND VGND VPWR VPWR _12689_ sky130_fd_sc_hd__mux2_1
X_25634_ _10055_ VGND VGND VPWR VPWR _11085_ sky130_fd_sc_hd__buf_2
XFILLER_0_116_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22846_ rvcpu.dp.rf.reg_file_arr\[8\]\[28\] rvcpu.dp.rf.reg_file_arr\[10\]\[28\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[28\] rvcpu.dp.rf.reg_file_arr\[11\]\[28\] _09424_
+ _09485_ VGND VGND VPWR VPWR _09984_ sky130_fd_sc_hd__mux4_1
XFILLER_0_211_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_935 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25565_ _10405_ _11042_ VGND VGND VPWR VPWR _11043_ sky130_fd_sc_hd__and2_1
X_28353_ _12651_ VGND VGND VPWR VPWR _03991_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22777_ _09918_ VGND VGND VPWR VPWR _01148_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27304_ _11965_ _12066_ VGND VGND VPWR VPWR _12067_ sky130_fd_sc_hd__and2_1
X_24516_ _09255_ VGND VGND VPWR VPWR _10452_ sky130_fd_sc_hd__clkbuf_2
X_21728_ rvcpu.dp.rf.reg_file_arr\[28\]\[18\] rvcpu.dp.rf.reg_file_arr\[30\]\[18\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[18\] rvcpu.dp.rf.reg_file_arr\[31\]\[18\] _08629_
+ _08683_ VGND VGND VPWR VPWR _08972_ sky130_fd_sc_hd__mux4_1
XFILLER_0_94_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28284_ _12614_ VGND VGND VPWR VPWR _03959_ sky130_fd_sc_hd__clkbuf_1
X_25496_ _10818_ net3960 _10999_ VGND VGND VPWR VPWR _11003_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27235_ _12029_ VGND VGND VPWR VPWR _12030_ sky130_fd_sc_hd__clkbuf_2
X_24447_ _10410_ _10406_ VGND VGND VPWR VPWR _10411_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_62_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23752__342 clknet_1_0__leaf__10200_ VGND VGND VPWR VPWR net468 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_62_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21659_ _08901_ _08903_ _08906_ _08626_ _08808_ VGND VGND VPWR VPWR _08907_ sky130_fd_sc_hd__a221o_1
XFILLER_0_136_388 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15180_ _13513_ _13722_ VGND VGND VPWR VPWR _13723_ sky130_fd_sc_hd__or2_1
X_27166_ _11946_ _11984_ VGND VGND VPWR VPWR _11989_ sky130_fd_sc_hd__and2_1
X_24378_ _09224_ net4354 _10367_ VGND VGND VPWR VPWR _10368_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26117_ net1728 _11386_ VGND VGND VPWR VPWR _11394_ sky130_fd_sc_hd__and2_1
XFILLER_0_201_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27097_ _11829_ _11941_ VGND VGND VPWR VPWR _11945_ sky130_fd_sc_hd__and2_1
XFILLER_0_127_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26048_ _11121_ net1810 _11350_ _11352_ VGND VGND VPWR VPWR _02985_ sky130_fd_sc_hd__a31o_1
XFILLER_0_132_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18870_ _05622_ _05478_ _05473_ VGND VGND VPWR VPWR _06213_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_219_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17821_ _05208_ VGND VGND VPWR VPWR rvcpu.dp.SrcBFW_Mux.y\[26\] sky130_fd_sc_hd__buf_1
X_29807_ net1145 _01542_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[1\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27999_ _09287_ VGND VGND VPWR VPWR _12460_ sky130_fd_sc_hd__clkbuf_2
Xhold5 rvcpu.dp.plem.lAuiPCM\[28\] VGND VGND VPWR VPWR net1155 sky130_fd_sc_hd__dlygate4sd3_1
X_29738_ net1084 _01473_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[21\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_17752_ _05151_ VGND VGND VPWR VPWR _01165_ sky130_fd_sc_hd__clkbuf_1
X_14964_ rvcpu.dp.pcreg.q\[7\] rvcpu.dp.pcreg.q\[6\] VGND VGND VPWR VPWR _13513_ sky130_fd_sc_hd__nand2_4
X_16703_ _04595_ VGND VGND VPWR VPWR _01690_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_169_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29669_ net1015 _01404_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[23\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_17683_ net2168 _13274_ _05081_ VGND VGND VPWR VPWR _05115_ sky130_fd_sc_hd__mux2_1
X_14895_ _13287_ _13288_ VGND VGND VPWR VPWR _13446_ sky130_fd_sc_hd__and2b_1
XFILLER_0_159_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31700_ clknet_leaf_43_clk _03158_ VGND VGND VPWR VPWR rvcpu.dp.pcreg.q\[18\] sky130_fd_sc_hd__dfxtp_1
X_19422_ _06717_ VGND VGND VPWR VPWR _06718_ sky130_fd_sc_hd__buf_4
XFILLER_0_199_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16634_ _14166_ net4042 _04551_ VGND VGND VPWR VPWR _04559_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32680_ clknet_leaf_181_clk _04102_ VGND VGND VPWR VPWR datamem.data_ram\[18\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31631_ clknet_leaf_48_clk net1235 VGND VGND VPWR VPWR rvcpu.dp.plmw.lAuiPCW\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19353_ _06648_ VGND VGND VPWR VPWR _06649_ sky130_fd_sc_hd__buf_6
XFILLER_0_168_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16565_ _14166_ net4301 _04514_ VGND VGND VPWR VPWR _04522_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18304_ _05668_ VGND VGND VPWR VPWR _05669_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_139_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15516_ _13767_ _13389_ _13780_ _13430_ VGND VGND VPWR VPWR _14043_ sky130_fd_sc_hd__o22a_1
XFILLER_0_167_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31562_ clknet_leaf_71_clk datamem.rd_data_mem\[12\] VGND VGND VPWR VPWR rvcpu.dp.plmw.ReadDataW\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_19284_ rvcpu.dp.plem.funct3M\[1\] rvcpu.dp.plem.funct3M\[0\] VGND VGND VPWR VPWR
+ _06580_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_139_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16496_ _04485_ VGND VGND VPWR VPWR _01795_ sky130_fd_sc_hd__clkbuf_1
X_23080__761 clknet_1_1__leaf__10091_ VGND VGND VPWR VPWR net887 sky130_fd_sc_hd__inv_2
XFILLER_0_84_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18235_ _05311_ _05318_ _05436_ _05438_ VGND VGND VPWR VPWR _05600_ sky130_fd_sc_hd__or4_1
X_30513_ clknet_leaf_219_clk _02248_ VGND VGND VPWR VPWR datamem.data_ram\[56\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_15447_ _13573_ _13973_ _13976_ _13977_ VGND VGND VPWR VPWR _13978_ sky130_fd_sc_hd__o211a_1
XFILLER_0_170_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_212_5575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31493_ clknet_leaf_45_clk rvcpu.dp.lAuiPCE\[19\] VGND VGND VPWR VPWR rvcpu.dp.plem.lAuiPCM\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_212_5586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23002__707 clknet_1_1__leaf__10085_ VGND VGND VPWR VPWR net833 sky130_fd_sc_hd__inv_2
XFILLER_0_111_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18166_ _05529_ _05530_ VGND VGND VPWR VPWR _05531_ sky130_fd_sc_hd__nor2_2
X_30444_ net782 _02179_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[29\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_15378_ _13419_ _13370_ _13416_ VGND VGND VPWR VPWR _13912_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_52_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap102 _05429_ VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_2
X_17117_ _04792_ VGND VGND VPWR VPWR _04815_ sky130_fd_sc_hd__clkbuf_4
Xhold405 datamem.data_ram\[54\]\[0\] VGND VGND VPWR VPWR net1555 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_208_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold416 datamem.data_ram\[6\]\[0\] VGND VGND VPWR VPWR net1566 sky130_fd_sc_hd__dlygate4sd3_1
X_18097_ _05463_ _05464_ VGND VGND VPWR VPWR _05465_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30375_ net721 _02110_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[3\]\[26\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_225_5903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold427 datamem.data_ram\[56\]\[2\] VGND VGND VPWR VPWR net1577 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32114_ clknet_leaf_97_clk _03536_ VGND VGND VPWR VPWR datamem.data_ram\[0\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold438 rvcpu.dp.plfd.PCD\[28\] VGND VGND VPWR VPWR net1588 sky130_fd_sc_hd__dlygate4sd3_1
Xhold449 datamem.data_ram\[47\]\[1\] VGND VGND VPWR VPWR net1599 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_4003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17048_ _04778_ VGND VGND VPWR VPWR _01512_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32045_ clknet_leaf_132_clk _03467_ VGND VGND VPWR VPWR datamem.data_ram\[49\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1105 datamem.data_ram\[13\]\[16\] VGND VGND VPWR VPWR net2255 sky130_fd_sc_hd__dlygate4sd3_1
X_18999_ _05645_ _06324_ _06325_ _06333_ VGND VGND VPWR VPWR _06334_ sky130_fd_sc_hd__a31o_1
XFILLER_0_104_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1116 datamem.data_ram\[28\]\[14\] VGND VGND VPWR VPWR net2266 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1127 rvcpu.dp.rf.reg_file_arr\[1\]\[26\] VGND VGND VPWR VPWR net2277 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1138 rvcpu.dp.rf.reg_file_arr\[20\]\[2\] VGND VGND VPWR VPWR net2288 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_105_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1149 rvcpu.dp.rf.reg_file_arr\[9\]\[21\] VGND VGND VPWR VPWR net2299 sky130_fd_sc_hd__dlygate4sd3_1
X_23922__478 clknet_1_1__leaf__10226_ VGND VGND VPWR VPWR net604 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_105_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20961_ datamem.data_ram\[62\]\[15\] datamem.data_ram\[63\]\[15\] _06651_ VGND VGND
+ VPWR VPWR _08250_ sky130_fd_sc_hd__mux2_1
X_32947_ clknet_leaf_211_clk _04369_ VGND VGND VPWR VPWR datamem.data_ram\[6\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_176_4711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_176_4722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22700_ rvcpu.dp.rf.reg_file_arr\[12\]\[20\] rvcpu.dp.rf.reg_file_arr\[13\]\[20\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[20\] rvcpu.dp.rf.reg_file_arr\[15\]\[20\] _09462_
+ _09721_ VGND VGND VPWR VPWR _09846_ sky130_fd_sc_hd__mux4_1
XFILLER_0_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23621__239 clknet_1_1__leaf__10180_ VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__inv_2
XFILLER_0_152_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32878_ clknet_leaf_54_clk _04300_ VGND VGND VPWR VPWR datamem.data_ram\[10\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20892_ _08125_ _08131_ _08153_ _08181_ VGND VGND VPWR VPWR _08182_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_49_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_778 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22631_ rvcpu.dp.rf.reg_file_arr\[20\]\[17\] rvcpu.dp.rf.reg_file_arr\[21\]\[17\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[17\] rvcpu.dp.rf.reg_file_arr\[23\]\[17\] _09517_
+ _09577_ VGND VGND VPWR VPWR _09780_ sky130_fd_sc_hd__mux4_2
X_31829_ clknet_leaf_106_clk _03283_ VGND VGND VPWR VPWR datamem.data_ram\[16\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_172_4619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_172_Left_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25350_ _10405_ _10923_ VGND VGND VPWR VPWR _10924_ sky130_fd_sc_hd__and2_1
XFILLER_0_193_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22562_ rvcpu.dp.rf.reg_file_arr\[0\]\[13\] rvcpu.dp.rf.reg_file_arr\[1\]\[13\] rvcpu.dp.rf.reg_file_arr\[2\]\[13\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[13\] _09714_ _09585_ VGND VGND VPWR VPWR _09715_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_91_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24301_ _09291_ net3821 _10316_ VGND VGND VPWR VPWR _10324_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21513_ _08511_ _08767_ VGND VGND VPWR VPWR _08768_ sky130_fd_sc_hd__nor2_1
X_23278__923 clknet_1_1__leaf__10129_ VGND VGND VPWR VPWR net1049 sky130_fd_sc_hd__inv_2
X_25281_ _10733_ net3216 _10878_ VGND VGND VPWR VPWR _10883_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_135_3740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22493_ _09482_ _09649_ VGND VGND VPWR VPWR _09650_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27020_ _11896_ VGND VGND VPWR VPWR _11897_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_17_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24232_ _09260_ net4006 _10279_ VGND VGND VPWR VPWR _10287_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_25_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21444_ _08702_ VGND VGND VPWR VPWR _01031_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_3637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23368__1004 clknet_1_0__leaf__10138_ VGND VGND VPWR VPWR net1130 sky130_fd_sc_hd__inv_2
XFILLER_0_47_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_131_3648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_550 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21375_ _08535_ VGND VGND VPWR VPWR _08636_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_96_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_1160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20326_ datamem.data_ram\[19\]\[4\] _06943_ _06993_ datamem.data_ram\[23\]\[4\] VGND
+ VGND VPWR VPWR _07618_ sky130_fd_sc_hd__a22o_1
X_28971_ _10066_ _12989_ VGND VGND VPWR VPWR _12994_ sky130_fd_sc_hd__and2_1
Xhold950 datamem.data_ram\[49\]\[22\] VGND VGND VPWR VPWR net2100 sky130_fd_sc_hd__dlygate4sd3_1
Xhold961 rvcpu.dp.rf.reg_file_arr\[16\]\[1\] VGND VGND VPWR VPWR net2111 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_181_Left_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold972 rvcpu.dp.rf.reg_file_arr\[1\]\[27\] VGND VGND VPWR VPWR net2122 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27922_ _12125_ net4435 _12412_ VGND VGND VPWR VPWR _12413_ sky130_fd_sc_hd__mux2_1
X_20257_ _06753_ _07544_ _07549_ _06985_ VGND VGND VPWR VPWR _07550_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_34_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold983 rvcpu.dp.rf.reg_file_arr\[10\]\[24\] VGND VGND VPWR VPWR net2133 sky130_fd_sc_hd__dlygate4sd3_1
Xhold994 datamem.data_ram\[0\]\[15\] VGND VGND VPWR VPWR net2144 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3030 datamem.data_ram\[53\]\[30\] VGND VGND VPWR VPWR net4180 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_34_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3041 datamem.data_ram\[18\]\[11\] VGND VGND VPWR VPWR net4191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3052 datamem.data_ram\[56\]\[9\] VGND VGND VPWR VPWR net4202 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27853_ _12128_ net2490 _12373_ VGND VGND VPWR VPWR _12375_ sky130_fd_sc_hd__mux2_1
Xhold3063 rvcpu.dp.rf.reg_file_arr\[24\]\[8\] VGND VGND VPWR VPWR net4213 sky130_fd_sc_hd__dlygate4sd3_1
X_23782__368 clknet_1_1__leaf__10204_ VGND VGND VPWR VPWR net494 sky130_fd_sc_hd__inv_2
Xhold3074 datamem.data_ram\[28\]\[12\] VGND VGND VPWR VPWR net4224 sky130_fd_sc_hd__dlygate4sd3_1
X_20188_ datamem.data_ram\[3\]\[11\] _06739_ _07477_ _07480_ VGND VGND VPWR VPWR _07481_
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_129_3588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2340 datamem.data_ram\[59\]\[11\] VGND VGND VPWR VPWR net3490 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3085 rvcpu.dp.rf.reg_file_arr\[0\]\[14\] VGND VGND VPWR VPWR net4235 sky130_fd_sc_hd__dlygate4sd3_1
X_26804_ _11684_ _11762_ VGND VGND VPWR VPWR _11766_ sky130_fd_sc_hd__and2_1
XFILLER_0_216_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2351 datamem.data_ram\[11\]\[20\] VGND VGND VPWR VPWR net3501 sky130_fd_sc_hd__dlygate4sd3_1
X_23250__897 clknet_1_1__leaf__10127_ VGND VGND VPWR VPWR net1023 sky130_fd_sc_hd__inv_2
Xhold3096 rvcpu.dp.rf.reg_file_arr\[13\]\[8\] VGND VGND VPWR VPWR net4246 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2362 rvcpu.dp.rf.reg_file_arr\[24\]\[12\] VGND VGND VPWR VPWR net3512 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2373 datamem.data_ram\[21\]\[20\] VGND VGND VPWR VPWR net3523 sky130_fd_sc_hd__dlygate4sd3_1
X_27784_ _12093_ net2792 _12326_ VGND VGND VPWR VPWR _12333_ sky130_fd_sc_hd__mux2_1
X_24996_ _10446_ net3024 _10715_ VGND VGND VPWR VPWR _10719_ sky130_fd_sc_hd__mux2_1
Xhold2384 datamem.data_ram\[16\]\[20\] VGND VGND VPWR VPWR net3534 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1650 datamem.data_ram\[47\]\[9\] VGND VGND VPWR VPWR net2800 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29523_ net885 _01258_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[28\]\[30\] sky130_fd_sc_hd__dfxtp_1
Xhold2395 datamem.data_ram\[2\]\[24\] VGND VGND VPWR VPWR net3545 sky130_fd_sc_hd__dlygate4sd3_1
X_26735_ _11723_ VGND VGND VPWR VPWR _11724_ sky130_fd_sc_hd__clkbuf_4
Xhold1661 datamem.data_ram\[10\]\[31\] VGND VGND VPWR VPWR net2811 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1672 datamem.data_ram\[48\]\[11\] VGND VGND VPWR VPWR net2822 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1683 rvcpu.dp.rf.reg_file_arr\[29\]\[15\] VGND VGND VPWR VPWR net2833 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1694 datamem.data_ram\[24\]\[9\] VGND VGND VPWR VPWR net2844 sky130_fd_sc_hd__dlygate4sd3_1
X_14680_ _13180_ VGND VGND VPWR VPWR _13245_ sky130_fd_sc_hd__buf_4
X_29454_ net816 _01189_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[30\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_26666_ _10063_ VGND VGND VPWR VPWR _11684_ sky130_fd_sc_hd__buf_2
XFILLER_0_19_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_190_Left_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28405_ _12679_ VGND VGND VPWR VPWR _04015_ sky130_fd_sc_hd__clkbuf_1
X_23596__216 clknet_1_0__leaf__10178_ VGND VGND VPWR VPWR net342 sky130_fd_sc_hd__inv_2
XFILLER_0_211_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__10266_ _10266_ VGND VGND VPWR VPWR clknet_0__10266_ sky130_fd_sc_hd__clkbuf_16
X_22829_ _09452_ _09965_ _09967_ _09795_ VGND VGND VPWR VPWR _09968_ sky130_fd_sc_hd__a211o_1
X_25617_ _10737_ net2720 net53 VGND VGND VPWR VPWR _11073_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29385_ clknet_leaf_269_clk _01120_ VGND VGND VPWR VPWR datamem.data_ram\[60\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_26597_ _11645_ _11640_ VGND VGND VPWR VPWR _11646_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_183_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28336_ _12642_ VGND VGND VPWR VPWR _03983_ sky130_fd_sc_hd__clkbuf_1
X_16350_ _14539_ VGND VGND VPWR VPWR _01863_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25548_ _11032_ VGND VGND VPWR VPWR _02805_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__10197_ _10197_ VGND VGND VPWR VPWR clknet_0__10197_ sky130_fd_sc_hd__clkbuf_16
X_23676__273 clknet_1_1__leaf__10193_ VGND VGND VPWR VPWR net399 sky130_fd_sc_hd__inv_2
XFILLER_0_54_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15301_ _13463_ _13838_ VGND VGND VPWR VPWR _13839_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_181_Right_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16281_ net2508 _14447_ _14500_ VGND VGND VPWR VPWR _14503_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_229_6003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25479_ _10048_ net35 _10996_ net1328 VGND VGND VPWR VPWR _02772_ sky130_fd_sc_hd__a22o_1
X_28267_ _12359_ net3435 _12603_ VGND VGND VPWR VPWR _12605_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_229_6014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_160_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_160_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_129_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_229_6025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18020_ rvcpu.dp.plde.ImmExtE\[0\] _05321_ VGND VGND VPWR VPWR _05390_ sky130_fd_sc_hd__nand2_1
X_27218_ _12005_ net1612 _12018_ _12020_ VGND VGND VPWR VPWR _03487_ sky130_fd_sc_hd__a31o_1
X_15232_ _13331_ _13284_ VGND VGND VPWR VPWR _13773_ sky130_fd_sc_hd__or2_1
XFILLER_0_151_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28198_ _12452_ net3477 net46 VGND VGND VPWR VPWR _12567_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15163_ _13419_ _13603_ _13673_ VGND VGND VPWR VPWR _13707_ sky130_fd_sc_hd__o21ai_1
X_27149_ _10072_ VGND VGND VPWR VPWR _11978_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30160_ net522 _01895_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[0\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_15094_ _13401_ _13484_ VGND VGND VPWR VPWR _13639_ sky130_fd_sc_hd__nor2_2
X_19971_ datamem.data_ram\[29\]\[18\] _06662_ _06646_ datamem.data_ram\[24\]\[18\]
+ VGND VGND VPWR VPWR _07265_ sky130_fd_sc_hd__o22a_1
XFILLER_0_120_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18922_ _06258_ _06259_ _06260_ _06261_ VGND VGND VPWR VPWR _06262_ sky130_fd_sc_hd__or4b_1
X_30091_ net453 _01826_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[11\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_219_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18853_ _06137_ _06196_ VGND VGND VPWR VPWR _06197_ sky130_fd_sc_hd__and2_1
X_17804_ _13172_ rvcpu.dp.plde.RD2E\[31\] _05196_ VGND VGND VPWR VPWR _05197_ sky130_fd_sc_hd__mux2_1
X_18784_ _05454_ _05513_ VGND VGND VPWR VPWR _06132_ sky130_fd_sc_hd__nor2_1
XFILLER_0_175_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15996_ net2090 _13251_ _14333_ VGND VGND VPWR VPWR _14336_ sky130_fd_sc_hd__mux2_1
X_32801_ clknet_leaf_159_clk _04223_ VGND VGND VPWR VPWR datamem.data_ram\[13\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17735_ _13251_ net3047 _05140_ VGND VGND VPWR VPWR _05143_ sky130_fd_sc_hd__mux2_1
X_14947_ _13353_ VGND VGND VPWR VPWR _13496_ sky130_fd_sc_hd__clkbuf_4
X_30993_ clknet_leaf_55_clk _02728_ VGND VGND VPWR VPWR datamem.data_ram\[13\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32732_ clknet_leaf_80_clk _04154_ VGND VGND VPWR VPWR datamem.data_ram\[16\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17666_ _05106_ VGND VGND VPWR VPWR _01206_ sky130_fd_sc_hd__clkbuf_1
X_14878_ _13303_ VGND VGND VPWR VPWR _13430_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23759__348 clknet_1_0__leaf__10201_ VGND VGND VPWR VPWR net474 sky130_fd_sc_hd__inv_2
X_19405_ _06700_ VGND VGND VPWR VPWR _06701_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_134_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16617_ _14149_ net3125 _04540_ VGND VGND VPWR VPWR _04550_ sky130_fd_sc_hd__mux2_1
X_32663_ clknet_leaf_86_clk _04085_ VGND VGND VPWR VPWR datamem.data_ram\[19\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_17597_ _13248_ net3515 _05068_ VGND VGND VPWR VPWR _05070_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_214_5626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_214_5637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31614_ clknet_leaf_13_clk net1251 VGND VGND VPWR VPWR rvcpu.dp.plmw.RdW\[0\] sky130_fd_sc_hd__dfxtp_2
X_19336_ _06631_ VGND VGND VPWR VPWR _06632_ sky130_fd_sc_hd__buf_8
XFILLER_0_169_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16548_ _14149_ net2328 _04503_ VGND VGND VPWR VPWR _04513_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32594_ clknet_leaf_285_clk _04016_ VGND VGND VPWR VPWR datamem.data_ram\[21\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19267_ _06566_ rvcpu.dp.plfd.InstrD\[6\] rvcpu.dp.plfd.InstrD\[4\] VGND VGND VPWR
+ VPWR _06567_ sky130_fd_sc_hd__nor3b_2
X_31545_ clknet_leaf_15_clk net1252 VGND VGND VPWR VPWR rvcpu.dp.plem.RdM\[3\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_151_clk clknet_5_28__leaf_clk VGND VGND VPWR VPWR clknet_leaf_151_clk
+ sky130_fd_sc_hd__clkbuf_8
X_16479_ _04476_ VGND VGND VPWR VPWR _01803_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18218_ _05380_ _05382_ VGND VGND VPWR VPWR _05583_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31476_ clknet_leaf_65_clk rvcpu.dp.lAuiPCE\[2\] VGND VGND VPWR VPWR rvcpu.dp.plem.lAuiPCM\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_19198_ rvcpu.dp.plde.ImmExtE\[23\] rvcpu.dp.plde.PCE\[23\] VGND VGND VPWR VPWR _06508_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_578 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18149_ _05498_ _05504_ _05513_ VGND VGND VPWR VPWR _05514_ sky130_fd_sc_hd__and3_1
X_30427_ net765 _02162_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[29\]\[6\] sky130_fd_sc_hd__dfxtp_1
Xhold202 datamem.data_ram\[18\]\[7\] VGND VGND VPWR VPWR net1352 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold213 _02930_ VGND VGND VPWR VPWR net1363 sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 datamem.data_ram\[3\]\[7\] VGND VGND VPWR VPWR net1374 sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 datamem.data_ram\[32\]\[6\] VGND VGND VPWR VPWR net1385 sky130_fd_sc_hd__dlygate4sd3_1
X_21160_ datamem.data_ram\[0\]\[23\] _06645_ _08448_ _06940_ _06676_ VGND VGND VPWR
+ VPWR _08449_ sky130_fd_sc_hd__o221a_1
Xhold246 datamem.data_ram\[32\]\[1\] VGND VGND VPWR VPWR net1396 sky130_fd_sc_hd__dlygate4sd3_1
X_30358_ net704 _02093_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[3\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold257 datamem.data_ram\[19\]\[3\] VGND VGND VPWR VPWR net1407 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_229_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold268 datamem.data_ram\[48\]\[0\] VGND VGND VPWR VPWR net1418 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_165_4445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20111_ datamem.data_ram\[18\]\[10\] _06804_ _07401_ _07404_ VGND VGND VPWR VPWR
+ _07405_ sky130_fd_sc_hd__o211a_1
Xhold279 datamem.data_ram\[5\]\[4\] VGND VGND VPWR VPWR net1429 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_165_4456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21091_ _07858_ _08375_ _08379_ _08355_ _06741_ VGND VGND VPWR VPWR _08380_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_165_4467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30289_ net635 _02024_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[5\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32028_ clknet_leaf_128_clk _03450_ VGND VGND VPWR VPWR datamem.data_ram\[26\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_20042_ datamem.data_ram\[3\]\[26\] _06729_ _06668_ datamem.data_ram\[7\]\[26\] _06677_
+ VGND VGND VPWR VPWR _07336_ sky130_fd_sc_hd__o221a_1
X_24850_ net112 _10599_ VGND VGND VPWR VPWR _10640_ sky130_fd_sc_hd__nor2_8
XFILLER_0_77_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24139__644 clknet_1_0__leaf__10261_ VGND VGND VPWR VPWR net770 sky130_fd_sc_hd__inv_2
X_24781_ _10465_ net2955 net94 VGND VGND VPWR VPWR _10603_ sky130_fd_sc_hd__mux2_1
X_21993_ rvcpu.dp.plem.WriteDataM\[0\] _09215_ _09219_ _09222_ VGND VGND VPWR VPWR
+ _09223_ sky130_fd_sc_hd__a31o_4
XTAP_TAPCELL_ROW_124_3463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_3474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_108 _07028_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26520_ _10048_ _11604_ _11605_ net1333 VGND VGND VPWR VPWR _03204_ sky130_fd_sc_hd__a22o_1
XANTENNA_119 _07203_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20944_ datamem.data_ram\[58\]\[22\] _06940_ _06934_ datamem.data_ram\[56\]\[22\]
+ VGND VGND VPWR VPWR _08234_ sky130_fd_sc_hd__o22a_1
X_23087__767 clknet_1_1__leaf__10102_ VGND VGND VPWR VPWR net893 sky130_fd_sc_hd__inv_2
XFILLER_0_221_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26451_ _11524_ rvcpu.ALUResultE\[22\] _11288_ VGND VGND VPWR VPWR _11579_ sky130_fd_sc_hd__a21o_1
XFILLER_0_138_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23818__401 clknet_1_0__leaf__10207_ VGND VGND VPWR VPWR net527 sky130_fd_sc_hd__inv_2
XFILLER_0_163_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20875_ datamem.data_ram\[55\]\[14\] _07020_ _08164_ rvcpu.dp.plem.ALUResultM\[6\]
+ VGND VGND VPWR VPWR _08165_ sky130_fd_sc_hd__o211a_1
XFILLER_0_178_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25402_ _10067_ _10950_ VGND VGND VPWR VPWR _10956_ sky130_fd_sc_hd__and2_1
XFILLER_0_113_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22614_ rvcpu.dp.rf.reg_file_arr\[28\]\[16\] rvcpu.dp.rf.reg_file_arr\[30\]\[16\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[16\] rvcpu.dp.rf.reg_file_arr\[31\]\[16\] _09446_
+ _09402_ VGND VGND VPWR VPWR _09764_ sky130_fd_sc_hd__mux4_1
X_26382_ _11525_ VGND VGND VPWR VPWR _11529_ sky130_fd_sc_hd__clkbuf_4
X_29170_ _09259_ net3713 net64 VGND VGND VPWR VPWR _13102_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23594_ clknet_1_1__leaf__10172_ VGND VGND VPWR VPWR _10178_ sky130_fd_sc_hd__buf_1
XFILLER_0_64_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25333_ _10912_ VGND VGND VPWR VPWR _02710_ sky130_fd_sc_hd__clkbuf_1
X_28121_ _12369_ net3464 _12519_ VGND VGND VPWR VPWR _12526_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22545_ _09622_ _09696_ _09698_ VGND VGND VPWR VPWR _09699_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_142_clk clknet_5_29__leaf_clk VGND VGND VPWR VPWR clknet_leaf_142_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_63_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_174_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_908 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25264_ _10538_ net1390 _10867_ _10873_ VGND VGND VPWR VPWR _02680_ sky130_fd_sc_hd__a31o_1
XFILLER_0_133_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28052_ _12489_ VGND VGND VPWR VPWR _03852_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_336 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22476_ rvcpu.dp.rf.reg_file_arr\[16\]\[9\] rvcpu.dp.rf.reg_file_arr\[17\]\[9\] rvcpu.dp.rf.reg_file_arr\[18\]\[9\]
+ rvcpu.dp.rf.reg_file_arr\[19\]\[9\] _09445_ _09447_ VGND VGND VPWR VPWR _09633_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_17_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27003_ _11863_ net1546 _11885_ _11887_ VGND VGND VPWR VPWR _03405_ sky130_fd_sc_hd__a31o_1
X_24215_ _09330_ net3279 _10270_ VGND VGND VPWR VPWR _10278_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21427_ _08540_ VGND VGND VPWR VPWR _08686_ sky130_fd_sc_hd__buf_4
X_25195_ _10835_ VGND VGND VPWR VPWR _02649_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21358_ _08612_ _08619_ rvcpu.dp.plde.BranchE VGND VGND VPWR VPWR _08620_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_60_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20309_ datamem.data_ram\[2\]\[4\] _06932_ _06976_ datamem.data_ram\[4\]\[4\] VGND
+ VGND VPWR VPWR _07601_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_57_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24077_ _10250_ VGND VGND VPWR VPWR _02116_ sky130_fd_sc_hd__clkbuf_1
X_28954_ _12745_ net3308 net67 VGND VGND VPWR VPWR _12984_ sky130_fd_sc_hd__mux2_1
Xhold780 rvcpu.dp.rf.reg_file_arr\[3\]\[31\] VGND VGND VPWR VPWR net1930 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21289_ _08550_ VGND VGND VPWR VPWR _08551_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold791 rvcpu.dp.rf.reg_file_arr\[5\]\[14\] VGND VGND VPWR VPWR net1941 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27905_ _12142_ net2962 net47 VGND VGND VPWR VPWR _12404_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28885_ _12762_ net3290 _12941_ VGND VGND VPWR VPWR _12947_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_216_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_53_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27836_ _12363_ net4216 _12357_ VGND VGND VPWR VPWR _12364_ sky130_fd_sc_hd__mux2_1
X_15850_ net2137 _13241_ _14247_ VGND VGND VPWR VPWR _14257_ sky130_fd_sc_hd__mux2_1
XFILLER_0_216_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23031__733 clknet_1_1__leaf__10088_ VGND VGND VPWR VPWR net859 sky130_fd_sc_hd__inv_2
Xhold2170 rvcpu.dp.rf.reg_file_arr\[8\]\[12\] VGND VGND VPWR VPWR net3320 sky130_fd_sc_hd__dlygate4sd3_1
X_14801_ _13312_ _13353_ VGND VGND VPWR VPWR _13354_ sky130_fd_sc_hd__nand2_1
Xhold2181 rvcpu.dp.rf.reg_file_arr\[8\]\[31\] VGND VGND VPWR VPWR net3331 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2192 datamem.data_ram\[57\]\[9\] VGND VGND VPWR VPWR net3342 sky130_fd_sc_hd__dlygate4sd3_1
X_15781_ _14170_ net2580 _14210_ VGND VGND VPWR VPWR _14220_ sky130_fd_sc_hd__mux2_1
X_27767_ _12323_ VGND VGND VPWR VPWR _03733_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_207_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24979_ _10472_ net4084 net101 VGND VGND VPWR VPWR _10710_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1480 datamem.data_ram\[2\]\[29\] VGND VGND VPWR VPWR net2630 sky130_fd_sc_hd__dlygate4sd3_1
X_29506_ net868 _01241_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[28\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_17520_ _13235_ net2798 _05021_ VGND VGND VPWR VPWR _05029_ sky130_fd_sc_hd__mux2_1
X_14732_ _13283_ _13284_ VGND VGND VPWR VPWR _13285_ sky130_fd_sc_hd__nand2_1
XFILLER_0_207_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26718_ _10751_ net3597 _11714_ VGND VGND VPWR VPWR _11715_ sky130_fd_sc_hd__mux2_1
Xhold1491 rvcpu.dp.rf.reg_file_arr\[16\]\[30\] VGND VGND VPWR VPWR net2641 sky130_fd_sc_hd__dlygate4sd3_1
X_27698_ _12138_ net2637 _12280_ VGND VGND VPWR VPWR _12287_ sky130_fd_sc_hd__mux2_1
XFILLER_0_200_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17451_ _04992_ VGND VGND VPWR VPWR _01315_ sky130_fd_sc_hd__clkbuf_1
X_29437_ net799 _01172_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[30\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_26649_ _11665_ net1372 _11662_ _11671_ VGND VGND VPWR VPWR _03267_ sky130_fd_sc_hd__a31o_1
X_14663_ _13231_ VGND VGND VPWR VPWR _13232_ sky130_fd_sc_hd__buf_4
XFILLER_0_131_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_211_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16402_ net3395 _14432_ _14561_ VGND VGND VPWR VPWR _14567_ sky130_fd_sc_hd__mux2_1
XFILLER_0_200_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17382_ _14164_ net2348 _04949_ VGND VGND VPWR VPWR _04956_ sky130_fd_sc_hd__mux2_1
X_29368_ clknet_leaf_202_clk _01103_ VGND VGND VPWR VPWR datamem.data_ram\[60\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_14594_ rvcpu.dp.plmw.RdW\[1\] _13178_ VGND VGND VPWR VPWR _13179_ sky130_fd_sc_hd__or2_4
XFILLER_0_82_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19121_ _06434_ VGND VGND VPWR VPWR _06440_ sky130_fd_sc_hd__inv_2
XFILLER_0_184_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28319_ _12633_ VGND VGND VPWR VPWR _03975_ sky130_fd_sc_hd__clkbuf_1
X_16333_ _14530_ VGND VGND VPWR VPWR _01871_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_211_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_133_clk clknet_5_27__leaf_clk VGND VGND VPWR VPWR clknet_leaf_133_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_171_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29299_ clknet_leaf_1_clk _01034_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD1E\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19052_ _06374_ _06376_ _06379_ VGND VGND VPWR VPWR _06380_ sky130_fd_sc_hd__o21a_1
X_31330_ clknet_leaf_16_clk _03033_ VGND VGND VPWR VPWR rvcpu.dp.plde.RdE\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16264_ net2455 _14430_ _14489_ VGND VGND VPWR VPWR _14494_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_656 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_201_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18003_ rvcpu.dp.plde.RD1E\[3\] _05265_ _05269_ _13268_ _05372_ VGND VGND VPWR VPWR
+ _05373_ sky130_fd_sc_hd__a221o_2
XTAP_TAPCELL_ROW_11_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15215_ _13361_ _13456_ _13555_ _13756_ VGND VGND VPWR VPWR _13757_ sky130_fd_sc_hd__or4_1
XFILLER_0_180_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31261_ clknet_leaf_20_clk _02964_ VGND VGND VPWR VPWR rvcpu.dp.plfd.InstrD\[19\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_152_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16195_ _14448_ VGND VGND VPWR VPWR _01935_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30212_ net566 _01947_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[8\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_15146_ _13403_ _13507_ VGND VGND VPWR VPWR _13690_ sky130_fd_sc_hd__and2_1
XFILLER_0_168_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31192_ clknet_leaf_49_clk _02895_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCPlus4D\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15077_ _13496_ _13621_ _13622_ _13429_ VGND VGND VPWR VPWR _13623_ sky130_fd_sc_hd__a22o_1
X_19954_ datamem.data_ram\[59\]\[18\] _06632_ _06704_ datamem.data_ram\[63\]\[18\]
+ VGND VGND VPWR VPWR _07248_ sky130_fd_sc_hd__o22a_1
X_30143_ net505 _01878_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[0\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_207_5452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_207_5463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_207_5474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18905_ _05698_ _05661_ _05691_ _06245_ VGND VGND VPWR VPWR _06246_ sky130_fd_sc_hd__a31o_1
X_19885_ datamem.data_ram\[24\]\[17\] _06698_ _07021_ datamem.data_ram\[31\]\[17\]
+ VGND VGND VPWR VPWR _07180_ sky130_fd_sc_hd__o22a_1
X_30074_ net436 _01809_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[12\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_4331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18836_ _06169_ _06170_ _06176_ _06181_ VGND VGND VPWR VPWR _06182_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_160_4342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_5264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_5275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23464__113 clknet_1_1__leaf__10157_ VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__inv_2
XFILLER_0_117_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_223_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18767_ _05311_ _05727_ _05730_ _06116_ _05820_ VGND VGND VPWR VPWR _06117_ sky130_fd_sc_hd__a221o_1
XFILLER_0_223_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15979_ net2106 _13226_ _14322_ VGND VGND VPWR VPWR _14327_ sky130_fd_sc_hd__mux2_1
XFILLER_0_175_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23993__527 clknet_1_0__leaf__10240_ VGND VGND VPWR VPWR net653 sky130_fd_sc_hd__inv_2
XFILLER_0_222_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23367__1003 clknet_1_0__leaf__10138_ VGND VGND VPWR VPWR net1129 sky130_fd_sc_hd__inv_2
X_17718_ _13226_ net2051 _05129_ VGND VGND VPWR VPWR _05134_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18698_ _06032_ _06051_ VGND VGND VPWR VPWR _06052_ sky130_fd_sc_hd__or2_1
X_30976_ clknet_leaf_161_clk _02711_ VGND VGND VPWR VPWR datamem.data_ram\[39\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32715_ clknet_leaf_252_clk _04137_ VGND VGND VPWR VPWR datamem.data_ram\[17\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17649_ _05097_ VGND VGND VPWR VPWR _01214_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_4282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_158_4293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23008__713 clknet_1_0__leaf__10085_ VGND VGND VPWR VPWR net839 sky130_fd_sc_hd__inv_2
X_32646_ clknet_leaf_157_clk _04068_ VGND VGND VPWR VPWR datamem.data_ram\[1\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_20660_ datamem.data_ram\[47\]\[29\] _07020_ _07947_ _07950_ VGND VGND VPWR VPWR
+ _07951_ sky130_fd_sc_hd__o211a_1
XFILLER_0_212_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19319_ rvcpu.dp.plem.ALUResultM\[3\] _06614_ VGND VGND VPWR VPWR _06615_ sky130_fd_sc_hd__nor2_8
XFILLER_0_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_124_clk clknet_5_27__leaf_clk VGND VGND VPWR VPWR clknet_leaf_124_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_129_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32577_ clknet_leaf_245_clk _03999_ VGND VGND VPWR VPWR datamem.data_ram\[21\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_20591_ datamem.data_ram\[19\]\[13\] _07831_ _07881_ _07820_ VGND VGND VPWR VPWR
+ _07882_ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22330_ _09492_ _09493_ _09449_ VGND VGND VPWR VPWR _09494_ sky130_fd_sc_hd__mux2_1
XFILLER_0_190_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31528_ clknet_leaf_28_clk net1201 VGND VGND VPWR VPWR rvcpu.dp.plem.PCPlus4M\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24030__561 clknet_1_0__leaf__10243_ VGND VGND VPWR VPWR net687 sky130_fd_sc_hd__inv_2
XFILLER_0_2_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22261_ _09422_ _09425_ _09426_ VGND VGND VPWR VPWR _09427_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_167_4507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31459_ clknet_leaf_75_clk rvcpu.dp.SrcBFW_Mux.y\[17\] VGND VGND VPWR VPWR rvcpu.dp.plem.WriteDataM\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21212_ _08487_ _06799_ _08490_ VGND VGND VPWR VPWR _04422_ sky130_fd_sc_hd__o21ai_1
X_22192_ _09368_ VGND VGND VPWR VPWR _01113_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_113_3197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__10238_ clknet_0__10238_ VGND VGND VPWR VPWR clknet_1_0__leaf__10238_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_130_158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23316__956 clknet_1_1__leaf__10134_ VGND VGND VPWR VPWR net1082 sky130_fd_sc_hd__inv_2
X_21143_ datamem.data_ram\[62\]\[23\] _06922_ _06917_ datamem.data_ram\[60\]\[23\]
+ VGND VGND VPWR VPWR _08432_ sky130_fd_sc_hd__o22a_1
X_23928__484 clknet_1_0__leaf__10226_ VGND VGND VPWR VPWR net610 sky130_fd_sc_hd__inv_2
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25951_ net2321 _11290_ _11286_ _11297_ VGND VGND VPWR VPWR _02943_ sky130_fd_sc_hd__o211a_1
X_21074_ datamem.data_ram\[44\]\[7\] _07825_ VGND VGND VPWR VPWR _08363_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_126_3514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_3525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20025_ _06769_ _07316_ _07318_ VGND VGND VPWR VPWR _07319_ sky130_fd_sc_hd__or3_1
X_24902_ _09225_ VGND VGND VPWR VPWR _10668_ sky130_fd_sc_hd__buf_8
X_28670_ _12751_ net4074 _12832_ VGND VGND VPWR VPWR _12833_ sky130_fd_sc_hd__mux2_1
X_25882_ net1679 _11256_ _11177_ _11257_ VGND VGND VPWR VPWR _02914_ sky130_fd_sc_hd__o211a_1
X_27621_ _12245_ VGND VGND VPWR VPWR _03665_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_225_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24833_ _10598_ _10630_ _10611_ VGND VGND VPWR VPWR _10631_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_87_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27552_ _12147_ net3087 net98 VGND VGND VPWR VPWR _12209_ sky130_fd_sc_hd__mux2_1
X_24764_ _10470_ net3434 _10589_ VGND VGND VPWR VPWR _10592_ sky130_fd_sc_hd__mux2_1
X_21976_ rvcpu.dp.rf.reg_file_arr\[12\]\[31\] rvcpu.dp.rf.reg_file_arr\[13\]\[31\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[31\] rvcpu.dp.rf.reg_file_arr\[15\]\[31\] _08628_
+ _08629_ VGND VGND VPWR VPWR _09207_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_29_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_5_2__f_clk clknet_2_0_0_clk VGND VGND VPWR VPWR clknet_5_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_55_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_179_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20927_ _07860_ _08211_ _08216_ VGND VGND VPWR VPWR _08217_ sky130_fd_sc_hd__o21a_1
X_27483_ _12130_ net3008 _12169_ VGND VGND VPWR VPWR _12172_ sky130_fd_sc_hd__mux2_1
X_24695_ _10444_ net4134 _10552_ VGND VGND VPWR VPWR _10555_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0__10103_ _10103_ VGND VGND VPWR VPWR clknet_0__10103_ sky130_fd_sc_hd__clkbuf_16
X_29222_ _11533_ net1383 _13122_ _13130_ VGND VGND VPWR VPWR _04381_ sky130_fd_sc_hd__a31o_1
X_23362__998 clknet_1_1__leaf__10138_ VGND VGND VPWR VPWR net1124 sky130_fd_sc_hd__inv_2
X_26434_ _06468_ _11539_ _11529_ _11196_ _11566_ VGND VGND VPWR VPWR _11567_ sky130_fd_sc_hd__a221o_1
XFILLER_0_166_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23646_ _10189_ VGND VGND VPWR VPWR _01746_ sky130_fd_sc_hd__clkbuf_1
X_20858_ _08146_ _08147_ _07840_ VGND VGND VPWR VPWR _08148_ sky130_fd_sc_hd__a21o_1
XFILLER_0_49_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29153_ _09290_ net2144 _13085_ VGND VGND VPWR VPWR _13093_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26365_ _11501_ net1524 _11510_ _11516_ VGND VGND VPWR VPWR _03138_ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_115_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_115_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_14_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_852 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20789_ datamem.data_ram\[23\]\[30\] _06761_ _07024_ datamem.data_ram\[20\]\[30\]
+ _06714_ VGND VGND VPWR VPWR _08079_ sky130_fd_sc_hd__o221a_1
XFILLER_0_148_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28104_ _12460_ net4412 net75 VGND VGND VPWR VPWR _12517_ sky130_fd_sc_hd__mux2_1
X_25316_ _10818_ net4038 _10899_ VGND VGND VPWR VPWR _10903_ sky130_fd_sc_hd__mux2_1
X_22528_ _09461_ _09680_ _09682_ _09474_ VGND VGND VPWR VPWR _09683_ sky130_fd_sc_hd__o211a_1
XFILLER_0_107_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26296_ net1720 _11478_ VGND VGND VPWR VPWR _11481_ sky130_fd_sc_hd__and2_1
X_29084_ _13056_ VGND VGND VPWR VPWR _04317_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28035_ _12443_ net2416 _12473_ VGND VGND VPWR VPWR _12480_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22459_ _09451_ _09616_ _09404_ VGND VGND VPWR VPWR _09617_ sky130_fd_sc_hd__o21a_1
X_25247_ _10863_ VGND VGND VPWR VPWR _02673_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15000_ _13391_ _13484_ VGND VGND VPWR VPWR _13548_ sky130_fd_sc_hd__or2_1
XFILLER_0_150_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25178_ _10825_ VGND VGND VPWR VPWR _02642_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23788__374 clknet_1_0__leaf__10204_ VGND VGND VPWR VPWR net500 sky130_fd_sc_hd__inv_2
XFILLER_0_32_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24129_ clknet_1_0__leaf__10244_ VGND VGND VPWR VPWR _10261_ sky130_fd_sc_hd__buf_1
XFILLER_0_20_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29986_ net356 _01721_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[14\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_28937_ _12974_ VGND VGND VPWR VPWR _04252_ sky130_fd_sc_hd__clkbuf_1
X_16951_ net3368 _14434_ _04720_ VGND VGND VPWR VPWR _04727_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15902_ _14274_ VGND VGND VPWR VPWR _14286_ sky130_fd_sc_hd__buf_4
XFILLER_0_218_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19670_ _06943_ VGND VGND VPWR VPWR _06966_ sky130_fd_sc_hd__buf_4
XFILLER_0_99_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_194_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16882_ _04690_ VGND VGND VPWR VPWR _01598_ sky130_fd_sc_hd__clkbuf_1
X_28868_ _12698_ net2796 _12932_ VGND VGND VPWR VPWR _12938_ sky130_fd_sc_hd__mux2_1
XFILLER_0_218_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_205_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18621_ _05978_ VGND VGND VPWR VPWR rvcpu.ALUResultE\[6\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_189_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27819_ _12352_ VGND VGND VPWR VPWR _03756_ sky130_fd_sc_hd__clkbuf_1
X_15833_ _14248_ VGND VGND VPWR VPWR _02105_ sky130_fd_sc_hd__clkbuf_1
X_28799_ _12901_ VGND VGND VPWR VPWR _04187_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_205_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30830_ clknet_leaf_155_clk _02565_ VGND VGND VPWR VPWR datamem.data_ram\[44\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_18552_ _05368_ _05401_ VGND VGND VPWR VPWR _05912_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_194_5150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15764_ _14211_ VGND VGND VPWR VPWR _02145_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_194_5161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17503_ _13210_ net2316 _05010_ VGND VGND VPWR VPWR _05020_ sky130_fd_sc_hd__mux2_1
X_14715_ rvcpu.dp.plmw.ALUResultW\[2\] rvcpu.dp.plmw.ReadDataW\[2\] rvcpu.dp.plmw.PCPlus4W\[2\]
+ rvcpu.dp.plmw.lAuiPCW\[2\] rvcpu.dp.plmw.ResultSrcW\[0\] rvcpu.dp.plmw.ResultSrcW\[1\]
+ VGND VGND VPWR VPWR _13271_ sky130_fd_sc_hd__mux4_2
XFILLER_0_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18483_ _05676_ _05843_ _05844_ VGND VGND VPWR VPWR _05845_ sky130_fd_sc_hd__o21ai_2
X_30761_ clknet_leaf_152_clk _02496_ VGND VGND VPWR VPWR datamem.data_ram\[47\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15695_ _14167_ VGND VGND VPWR VPWR _02170_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_213_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_190_5047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_450 _07860_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_190_5058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32500_ clknet_leaf_253_clk _03922_ VGND VGND VPWR VPWR datamem.data_ram\[25\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_461 _08735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17434_ _04983_ VGND VGND VPWR VPWR _01323_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_472 _09059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14646_ rvcpu.dp.plmw.ALUResultW\[19\] rvcpu.dp.plmw.ReadDataW\[19\] rvcpu.dp.plmw.PCPlus4W\[19\]
+ rvcpu.dp.plmw.lAuiPCW\[19\] _13169_ _13171_ VGND VGND VPWR VPWR _13219_ sky130_fd_sc_hd__mux4_2
XFILLER_0_28_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_483 _09317_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_30692_ clknet_leaf_280_clk _02427_ VGND VGND VPWR VPWR datamem.data_ram\[4\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_494 _09892_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32431_ clknet_leaf_274_clk _03853_ VGND VGND VPWR VPWR datamem.data_ram\[28\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_106_clk clknet_5_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_106_clk
+ sky130_fd_sc_hd__clkbuf_8
X_17365_ _14147_ net2930 _04938_ VGND VGND VPWR VPWR _04947_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_19 _06613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19104_ _06425_ rvcpu.dp.plde.ImmExtE\[11\] _06419_ VGND VGND VPWR VPWR _06426_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16316_ net2608 _14482_ _14511_ VGND VGND VPWR VPWR _14521_ sky130_fd_sc_hd__mux2_1
X_32362_ clknet_leaf_93_clk _03784_ VGND VGND VPWR VPWR datamem.data_ram\[2\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_17296_ _04910_ VGND VGND VPWR VPWR _01396_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19035_ _06365_ rvcpu.dp.plde.ImmExtE\[2\] _06355_ VGND VGND VPWR VPWR _06366_ sky130_fd_sc_hd__mux2_1
X_31313_ clknet_leaf_45_clk _03016_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCPlus4E\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23574__196 clknet_1_1__leaf__10176_ VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__inv_2
XFILLER_0_141_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16247_ _14483_ VGND VGND VPWR VPWR _01918_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_209_5503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32293_ clknet_leaf_226_clk _03715_ VGND VGND VPWR VPWR datamem.data_ram\[32\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_209_5514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31244_ clknet_leaf_21_clk _02947_ VGND VGND VPWR VPWR rvcpu.dp.plfd.InstrD\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_16178_ net3134 _14436_ _14422_ VGND VGND VPWR VPWR _14437_ sky130_fd_sc_hd__mux2_1
X_15129_ _13346_ _13389_ _13317_ VGND VGND VPWR VPWR _13674_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23038__739 clknet_1_1__leaf__10089_ VGND VGND VPWR VPWR net865 sky130_fd_sc_hd__inv_2
X_31175_ clknet_leaf_210_clk _02878_ VGND VGND VPWR VPWR datamem.data_ram\[5\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30126_ net488 _01861_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[10\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_19937_ datamem.data_ram\[35\]\[18\] _06634_ _07230_ datamem.data_ram\[36\]\[18\]
+ VGND VGND VPWR VPWR _07231_ sky130_fd_sc_hd__o22a_1
Xhold2906 datamem.data_ram\[19\]\[24\] VGND VGND VPWR VPWR net4056 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2917 rvcpu.dp.rf.reg_file_arr\[10\]\[12\] VGND VGND VPWR VPWR net4067 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2928 datamem.data_ram\[23\]\[13\] VGND VGND VPWR VPWR net4078 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2939 rvcpu.dp.rf.reg_file_arr\[27\]\[30\] VGND VGND VPWR VPWR net4089 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24060__587 clknet_1_1__leaf__10247_ VGND VGND VPWR VPWR net713 sky130_fd_sc_hd__inv_2
X_19868_ datamem.data_ram\[11\]\[1\] _06966_ _07161_ _07162_ VGND VGND VPWR VPWR _07163_
+ sky130_fd_sc_hd__a211o_1
X_30057_ net419 _01792_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[12\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_218_1221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18819_ _05338_ _05453_ _05504_ _05513_ VGND VGND VPWR VPWR _06165_ sky130_fd_sc_hd__o211a_1
X_19799_ datamem.data_ram\[59\]\[9\] _06636_ _07090_ _07093_ VGND VGND VPWR VPWR _07094_
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_121_3400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_3411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21830_ _08682_ _09066_ _09068_ _08558_ VGND VGND VPWR VPWR _09069_ sky130_fd_sc_hd__o211a_1
XFILLER_0_211_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21761_ _09003_ VGND VGND VPWR VPWR _01047_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30959_ clknet_leaf_163_clk _02694_ VGND VGND VPWR VPWR datamem.data_ram\[3\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20712_ datamem.data_ram\[28\]\[5\] _07123_ _07999_ _08002_ VGND VGND VPWR VPWR _08003_
+ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_82_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_854 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24480_ _09351_ _10327_ _10366_ VGND VGND VPWR VPWR _10430_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_148_556 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21692_ rvcpu.dp.rf.reg_file_arr\[24\]\[16\] rvcpu.dp.rf.reg_file_arr\[25\]\[16\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[16\] rvcpu.dp.rf.reg_file_arr\[27\]\[16\] _08525_
+ _08528_ VGND VGND VPWR VPWR _08938_ sky130_fd_sc_hd__mux4_1
XFILLER_0_77_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32629_ clknet_leaf_95_clk _04051_ VGND VGND VPWR VPWR datamem.data_ram\[1\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20643_ datamem.data_ram\[19\]\[29\] _06829_ _07932_ _07933_ VGND VGND VPWR VPWR
+ _07934_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_119_3351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26150_ _11411_ VGND VGND VPWR VPWR _03027_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20574_ datamem.data_ram\[32\]\[13\] datamem.data_ram\[33\]\[13\] datamem.data_ram\[34\]\[13\]
+ datamem.data_ram\[35\]\[13\] _07835_ _07821_ VGND VGND VPWR VPWR _07865_ sky130_fd_sc_hd__mux4_1
XFILLER_0_33_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_115_3248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25101_ _10782_ _10779_ _10781_ net1466 VGND VGND VPWR VPWR _02608_ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22313_ _09477_ VGND VGND VPWR VPWR _09478_ sky130_fd_sc_hd__buf_6
X_26081_ _06573_ _11372_ VGND VGND VPWR VPWR _11373_ sky130_fd_sc_hd__and2_1
XFILLER_0_144_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_115_3259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25032_ _10741_ _10601_ _10705_ VGND VGND VPWR VPWR _10742_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_186_4949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22244_ _09407_ _09409_ _09380_ VGND VGND VPWR VPWR _09410_ sky130_fd_sc_hd__mux2_1
XFILLER_0_225_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29840_ net218 _01575_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[18\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22175_ _09326_ net3909 _09352_ VGND VGND VPWR VPWR _09359_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_218_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21126_ _07820_ _08413_ _08414_ _07844_ VGND VGND VPWR VPWR _08415_ sky130_fd_sc_hd__o211a_1
X_29771_ net1117 _01506_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[20\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_26983_ _10751_ net3670 _11875_ VGND VGND VPWR VPWR _11876_ sky130_fd_sc_hd__mux2_1
X_23861__424 clknet_1_0__leaf__10219_ VGND VGND VPWR VPWR net550 sky130_fd_sc_hd__inv_2
XFILLER_0_195_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_50_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28722_ _12860_ VGND VGND VPWR VPWR _04151_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_89_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25934_ net1668 _11275_ _11286_ _11287_ VGND VGND VPWR VPWR _02936_ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_89_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21057_ datamem.data_ram\[44\]\[31\] datamem.data_ram\[45\]\[31\] _07825_ VGND VGND
+ VPWR VPWR _08346_ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_145_3967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20008_ datamem.data_ram\[56\]\[2\] _06936_ _06953_ datamem.data_ram\[60\]\[2\] VGND
+ VGND VPWR VPWR _07302_ sky130_fd_sc_hd__a22o_1
X_28653_ _12687_ net4117 _12823_ VGND VGND VPWR VPWR _12824_ sky130_fd_sc_hd__mux2_1
XFILLER_0_213_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25865_ rvcpu.dp.pcreg.q\[29\] _11239_ VGND VGND VPWR VPWR _11244_ sky130_fd_sc_hd__xor2_1
XFILLER_0_92_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_213_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_202_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_198_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27604_ _12236_ VGND VGND VPWR VPWR _03657_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24816_ _10385_ net2849 _10621_ VGND VGND VPWR VPWR _10622_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28584_ _12734_ net2928 _12786_ VGND VGND VPWR VPWR _12787_ sky130_fd_sc_hd__mux2_1
XFILLER_0_213_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25796_ rvcpu.dp.pcreg.q\[14\] _11182_ rvcpu.dp.pcreg.q\[15\] VGND VGND VPWR VPWR
+ _11189_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_96_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27535_ _12130_ net2679 _12197_ VGND VGND VPWR VPWR _12200_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24747_ _10390_ net3841 _10580_ VGND VGND VPWR VPWR _10583_ sky130_fd_sc_hd__mux2_1
X_21959_ rvcpu.dp.rf.reg_file_arr\[12\]\[30\] rvcpu.dp.rf.reg_file_arr\[13\]\[30\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[30\] rvcpu.dp.rf.reg_file_arr\[15\]\[30\] _08549_
+ _08553_ VGND VGND VPWR VPWR _09191_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_48_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15480_ _13320_ _13285_ _13349_ VGND VGND VPWR VPWR _14009_ sky130_fd_sc_hd__or3_2
X_27466_ _12162_ VGND VGND VPWR VPWR _03593_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_104_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24678_ _10390_ net3823 _10543_ VGND VGND VPWR VPWR _10546_ sky130_fd_sc_hd__mux2_1
XFILLER_0_204_54 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29205_ _13120_ VGND VGND VPWR VPWR _04374_ sky130_fd_sc_hd__clkbuf_1
X_26417_ net4450 _11542_ _11555_ _11534_ VGND VGND VPWR VPWR _03151_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_13_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27397_ _12118_ VGND VGND VPWR VPWR _03568_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_193_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29136_ _09259_ net4164 _13076_ VGND VGND VPWR VPWR _13084_ sky130_fd_sc_hd__mux2_1
X_17150_ _14137_ net3935 _04829_ VGND VGND VPWR VPWR _04833_ sky130_fd_sc_hd__mux2_1
X_26348_ _10064_ _11507_ _11508_ net1329 VGND VGND VPWR VPWR _03129_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16101_ _14392_ VGND VGND VPWR VPWR _01973_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17081_ _04796_ VGND VGND VPWR VPWR _01497_ sky130_fd_sc_hd__clkbuf_1
X_29067_ _13047_ VGND VGND VPWR VPWR _04309_ sky130_fd_sc_hd__clkbuf_1
X_26279_ net1840 _11467_ VGND VGND VPWR VPWR _11472_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_220_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28018_ _12369_ net4138 net97 VGND VGND VPWR VPWR _12471_ sky130_fd_sc_hd__mux2_1
X_16032_ net2119 _13201_ _14349_ VGND VGND VPWR VPWR _14356_ sky130_fd_sc_hd__mux2_1
XFILLER_0_204_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23366__1002 clknet_1_0__leaf__10138_ VGND VGND VPWR VPWR net1128 sky130_fd_sc_hd__inv_2
XFILLER_0_21_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_204_5400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_199_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17983_ rvcpu.dp.plde.ImmExtE\[6\] rvcpu.dp.SrcBFW_Mux.y\[6\] _05277_ VGND VGND VPWR
+ VPWR _05353_ sky130_fd_sc_hd__mux2_1
X_29969_ net339 _01704_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[15\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_24169__11 clknet_1_0__leaf__10264_ VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__inv_2
X_19722_ _06590_ _06913_ _07017_ VGND VGND VPWR VPWR _04415_ sky130_fd_sc_hd__o21ai_1
X_16934_ _04717_ VGND VGND VPWR VPWR _01573_ sky130_fd_sc_hd__clkbuf_1
X_32980_ clknet_leaf_272_clk _04402_ VGND VGND VPWR VPWR datamem.data_ram\[63\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_196_5201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19653_ _06948_ VGND VGND VPWR VPWR _06949_ sky130_fd_sc_hd__clkbuf_8
X_31931_ clknet_leaf_122_clk _03353_ VGND VGND VPWR VPWR datamem.data_ram\[60\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_221_5791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16865_ net2480 _14484_ _04647_ VGND VGND VPWR VPWR _04681_ sky130_fd_sc_hd__mux2_1
XFILLER_0_189_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18604_ _05799_ _05843_ _05961_ VGND VGND VPWR VPWR _05962_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_192_5109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15816_ _14239_ VGND VGND VPWR VPWR _02113_ sky130_fd_sc_hd__clkbuf_1
X_31862_ clknet_leaf_110_clk _03316_ VGND VGND VPWR VPWR datamem.data_ram\[62\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_19584_ datamem.data_ram\[38\]\[8\] _06628_ _06876_ _06879_ VGND VGND VPWR VPWR _06880_
+ sky130_fd_sc_hd__o211a_1
X_16796_ _04644_ VGND VGND VPWR VPWR _01646_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18535_ _05803_ _05895_ _05668_ VGND VGND VPWR VPWR _05896_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30813_ clknet_leaf_264_clk _02548_ VGND VGND VPWR VPWR datamem.data_ram\[45\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15747_ _14202_ VGND VGND VPWR VPWR _02153_ sky130_fd_sc_hd__clkbuf_1
X_31793_ clknet_leaf_210_clk _03247_ VGND VGND VPWR VPWR datamem.data_ram\[2\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30744_ clknet_leaf_142_clk _02479_ VGND VGND VPWR VPWR datamem.data_ram\[48\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_18466_ _05825_ _05828_ _05380_ VGND VGND VPWR VPWR _05829_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15678_ _13219_ VGND VGND VPWR VPWR _14156_ sky130_fd_sc_hd__buf_4
XFILLER_0_74_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_280 _13257_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_291 _13348_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_185_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17417_ _14127_ net3236 _04974_ VGND VGND VPWR VPWR _04975_ sky130_fd_sc_hd__mux2_1
X_14629_ rvcpu.dp.plmw.ALUResultW\[23\] rvcpu.dp.plmw.ReadDataW\[23\] rvcpu.dp.plmw.PCPlus4W\[23\]
+ rvcpu.dp.plmw.lAuiPCW\[23\] _13169_ _13171_ VGND VGND VPWR VPWR _13206_ sky130_fd_sc_hd__mux4_2
XFILLER_0_157_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_695 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_4116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18397_ _05539_ _05545_ _05682_ VGND VGND VPWR VPWR _05761_ sky130_fd_sc_hd__mux2_1
X_30675_ clknet_leaf_178_clk _02410_ VGND VGND VPWR VPWR datamem.data_ram\[50\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_151_4127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32414_ clknet_leaf_245_clk _03836_ VGND VGND VPWR VPWR datamem.data_ram\[28\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17348_ _04937_ VGND VGND VPWR VPWR _04938_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_16_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32345_ clknet_leaf_77_clk _03767_ VGND VGND VPWR VPWR datamem.data_ram\[30\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload200 clknet_leaf_193_clk VGND VGND VPWR VPWR clkload200/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_130_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload211 clknet_leaf_205_clk VGND VGND VPWR VPWR clkload211/X sky130_fd_sc_hd__clkbuf_4
X_17279_ _04464_ _04900_ VGND VGND VPWR VPWR _04901_ sky130_fd_sc_hd__and2_2
Xclkload222 clknet_leaf_159_clk VGND VGND VPWR VPWR clkload222/Y sky130_fd_sc_hd__bufinv_16
Xclkload233 clknet_leaf_112_clk VGND VGND VPWR VPWR clkload233/Y sky130_fd_sc_hd__inv_6
X_19018_ _06337_ _06338_ _06351_ VGND VGND VPWR VPWR rvcpu.ALUResultE\[30\] sky130_fd_sc_hd__o21bai_2
XFILLER_0_70_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload244 clknet_leaf_134_clk VGND VGND VPWR VPWR clkload244/Y sky130_fd_sc_hd__clkinv_4
Xclkload255 clknet_leaf_141_clk VGND VGND VPWR VPWR clkload255/Y sky130_fd_sc_hd__inv_6
X_20290_ datamem.data_ram\[20\]\[19\] _06688_ _07581_ _07582_ VGND VGND VPWR VPWR
+ _07583_ sky130_fd_sc_hd__o211a_1
X_32276_ clknet_leaf_161_clk _03698_ VGND VGND VPWR VPWR datamem.data_ram\[33\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_228_5956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload266 clknet_leaf_125_clk VGND VGND VPWR VPWR clkload266/Y sky130_fd_sc_hd__clkinv_1
XFILLER_0_24_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_228_5967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload277 clknet_leaf_140_clk VGND VGND VPWR VPWR clkload277/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_228_5978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload288 clknet_1_1__leaf__10240_ VGND VGND VPWR VPWR clkload288/Y sky130_fd_sc_hd__clkinvlp_4
X_31227_ clknet_leaf_43_clk net1363 VGND VGND VPWR VPWR rvcpu.dp.plfd.PCD\[16\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_149_4067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload299 clknet_1_0__leaf__10206_ VGND VGND VPWR VPWR clkload299/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_149_4078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_181_4835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_181_4846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31158_ clknet_leaf_69_clk rvcpu.ALUResultE\[17\] VGND VGND VPWR VPWR rvcpu.dp.plem.ALUResultM\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2703 datamem.data_ram\[50\]\[16\] VGND VGND VPWR VPWR net3853 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2714 rvcpu.dp.rf.reg_file_arr\[16\]\[11\] VGND VGND VPWR VPWR net3864 sky130_fd_sc_hd__dlygate4sd3_1
X_23999__533 clknet_1_0__leaf__10240_ VGND VGND VPWR VPWR net659 sky130_fd_sc_hd__inv_2
Xhold2725 datamem.data_ram\[23\]\[8\] VGND VGND VPWR VPWR net3875 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30109_ net471 _01844_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[10\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_71_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2736 datamem.data_ram\[47\]\[29\] VGND VGND VPWR VPWR net3886 sky130_fd_sc_hd__dlygate4sd3_1
X_31089_ clknet_leaf_107_clk _02824_ VGND VGND VPWR VPWR datamem.data_ram\[21\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2747 datamem.data_ram\[1\]\[10\] VGND VGND VPWR VPWR net3897 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2758 datamem.data_ram\[41\]\[16\] VGND VGND VPWR VPWR net3908 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2769 datamem.data_ram\[41\]\[29\] VGND VGND VPWR VPWR net3919 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22931_ _10056_ net1569 _10046_ _10062_ VGND VGND VPWR VPWR _01158_ sky130_fd_sc_hd__a31o_1
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_84_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25650_ _10048_ _11094_ _11095_ net1318 VGND VGND VPWR VPWR _02844_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22862_ _09429_ _09996_ _09998_ VGND VGND VPWR VPWR _09999_ sky130_fd_sc_hd__a21o_1
XFILLER_0_74_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_140_3853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_3864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_179_4786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24601_ _10465_ net2572 _10502_ VGND VGND VPWR VPWR _10503_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_179_4797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21813_ rvcpu.dp.rf.reg_file_arr\[12\]\[22\] rvcpu.dp.rf.reg_file_arr\[13\]\[22\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[22\] rvcpu.dp.rf.reg_file_arr\[15\]\[22\] _08696_
+ _08553_ VGND VGND VPWR VPWR _09053_ sky130_fd_sc_hd__mux4_1
Xwire41 _12868_ VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__buf_4
X_25581_ _11018_ net1444 _11041_ _11051_ VGND VGND VPWR VPWR _02819_ sky130_fd_sc_hd__a31o_1
XFILLER_0_195_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_1276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22793_ _09469_ _09933_ VGND VGND VPWR VPWR _09934_ sky130_fd_sc_hd__or2_1
X_27320_ _10979_ _10049_ _10051_ VGND VGND VPWR VPWR _12075_ sky130_fd_sc_hd__and3_1
XFILLER_0_148_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21744_ _08514_ _08986_ VGND VGND VPWR VPWR _08987_ sky130_fd_sc_hd__or2_1
X_24532_ _10461_ VGND VGND VPWR VPWR _02360_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_176_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27251_ _12036_ net1459 _12030_ _12039_ VGND VGND VPWR VPWR _03501_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_43_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24463_ _10113_ _10327_ _10366_ VGND VGND VPWR VPWR _10421_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_43_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21675_ rvcpu.dp.rf.reg_file_arr\[24\]\[15\] rvcpu.dp.rf.reg_file_arr\[25\]\[15\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[15\] rvcpu.dp.rf.reg_file_arr\[27\]\[15\] _08548_
+ _08526_ VGND VGND VPWR VPWR _08922_ sky130_fd_sc_hd__mux4_1
X_24110__617 clknet_1_0__leaf__10259_ VGND VGND VPWR VPWR net743 sky130_fd_sc_hd__inv_2
XFILLER_0_108_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26202_ _11362_ net116 VGND VGND VPWR VPWR _11439_ sky130_fd_sc_hd__and2_1
XFILLER_0_136_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20626_ datamem.data_ram\[8\]\[13\] _06647_ _06634_ datamem.data_ram\[11\]\[13\]
+ _07916_ VGND VGND VPWR VPWR _07917_ sky130_fd_sc_hd__o221a_1
X_27182_ _11970_ _11996_ VGND VGND VPWR VPWR _11999_ sky130_fd_sc_hd__and2_1
X_24394_ _09226_ _10347_ _10366_ VGND VGND VPWR VPWR _10376_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_46_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26133_ _11402_ VGND VGND VPWR VPWR _03019_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20557_ datamem.data_ram\[15\]\[21\] _07020_ _06688_ datamem.data_ram\[12\]\[21\]
+ VGND VGND VPWR VPWR _07848_ sky130_fd_sc_hd__o22a_1
XFILLER_0_61_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26064_ rvcpu.c.ad.opb5 _06572_ VGND VGND VPWR VPWR _11361_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20488_ _06715_ _07763_ _07768_ _07779_ VGND VGND VPWR VPWR _07780_ sky130_fd_sc_hd__o31a_1
XFILLER_0_85_1199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_225_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22227_ _09392_ VGND VGND VPWR VPWR _09393_ sky130_fd_sc_hd__buf_4
X_25015_ _10730_ VGND VGND VPWR VPWR _02574_ sky130_fd_sc_hd__clkbuf_1
X_29823_ net201 _01558_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[1\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_22158_ _09291_ net2759 net62 VGND VGND VPWR VPWR _09349_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21109_ _07838_ _08395_ _08397_ _07844_ VGND VGND VPWR VPWR _08398_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_7_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29754_ net1100 _01489_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[21\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_14980_ _13335_ _13369_ VGND VGND VPWR VPWR _13528_ sky130_fd_sc_hd__nor2_4
X_26966_ _11822_ _11866_ VGND VGND VPWR VPWR _11867_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_7_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22089_ _09298_ net2946 _09302_ VGND VGND VPWR VPWR _09303_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28705_ _12851_ VGND VGND VPWR VPWR _04143_ sky130_fd_sc_hd__clkbuf_1
X_25917_ net1803 _11263_ VGND VGND VPWR VPWR _11278_ sky130_fd_sc_hd__or2_1
XFILLER_0_156_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29685_ net1031 _01420_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[23\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26897_ _10047_ VGND VGND VPWR VPWR _11822_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_191_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28636_ _12734_ net3088 net71 VGND VGND VPWR VPWR _12815_ sky130_fd_sc_hd__mux2_1
X_16650_ _04567_ VGND VGND VPWR VPWR _01715_ sky130_fd_sc_hd__clkbuf_1
X_25848_ _11230_ VGND VGND VPWR VPWR _02907_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_198_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15601_ _14108_ VGND VGND VPWR VPWR _02205_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_18_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28567_ _12751_ net2060 _12777_ VGND VGND VPWR VPWR _12778_ sky130_fd_sc_hd__mux2_1
X_16581_ _04530_ VGND VGND VPWR VPWR _01755_ sky130_fd_sc_hd__clkbuf_1
X_25779_ _11174_ _11175_ _11157_ VGND VGND VPWR VPWR _11176_ sky130_fd_sc_hd__a21o_1
XFILLER_0_85_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18320_ _05580_ _05684_ _05395_ VGND VGND VPWR VPWR _05685_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15532_ _13319_ _14057_ _13572_ VGND VGND VPWR VPWR _14058_ sky130_fd_sc_hd__a21oi_1
X_27518_ _12085_ net3788 net99 VGND VGND VPWR VPWR _12191_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_201_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28498_ _12727_ net1640 _12723_ _12733_ VGND VGND VPWR VPWR _04054_ sky130_fd_sc_hd__a31o_1
XFILLER_0_167_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18251_ _05599_ _05602_ _05615_ VGND VGND VPWR VPWR _05616_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_127_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15463_ _13988_ _13989_ _13992_ _13499_ VGND VGND VPWR VPWR _13993_ sky130_fd_sc_hd__a31o_1
X_27449_ _12151_ net3843 net84 VGND VGND VPWR VPWR _12152_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_182_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17202_ _14189_ net2546 _04851_ VGND VGND VPWR VPWR _04860_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_131 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18182_ _05545_ _05546_ VGND VGND VPWR VPWR _05547_ sky130_fd_sc_hd__and2_1
X_30460_ net138 _02195_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[19\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15394_ _13665_ _13323_ _13666_ VGND VGND VPWR VPWR _13927_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_64_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17133_ _04823_ VGND VGND VPWR VPWR _01472_ sky130_fd_sc_hd__clkbuf_1
X_29119_ _09290_ net2448 _13067_ VGND VGND VPWR VPWR _13075_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30391_ net729 _02126_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[31\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32130_ clknet_leaf_212_clk _03552_ VGND VGND VPWR VPWR datamem.data_ram\[10\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold609 datamem.data_ram\[58\]\[1\] VGND VGND VPWR VPWR net1759 sky130_fd_sc_hd__dlygate4sd3_1
X_17064_ net3904 _14478_ _04779_ VGND VGND VPWR VPWR _04787_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16015_ _14345_ VGND VGND VPWR VPWR _02020_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32061_ clknet_leaf_118_clk _03483_ VGND VGND VPWR VPWR datamem.data_ram\[48\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31012_ clknet_leaf_165_clk _02747_ VGND VGND VPWR VPWR datamem.data_ram\[11\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_223_5842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_223_5853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17966_ _05311_ _05318_ _05333_ _05336_ VGND VGND VPWR VPWR _05337_ sky130_fd_sc_hd__a31oi_1
Xhold1309 datamem.data_ram\[3\]\[14\] VGND VGND VPWR VPWR net2459 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19705_ datamem.data_ram\[6\]\[0\] _06952_ _06973_ datamem.data_ram\[0\]\[0\] VGND
+ VGND VPWR VPWR _07001_ sky130_fd_sc_hd__a22o_1
X_16917_ net2161 _14468_ _04706_ VGND VGND VPWR VPWR _04709_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32963_ clknet_leaf_199_clk _04385_ VGND VGND VPWR VPWR datamem.data_ram\[63\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_17897_ _05269_ VGND VGND VPWR VPWR _05270_ sky130_fd_sc_hd__clkbuf_4
X_19636_ _06931_ VGND VGND VPWR VPWR _06932_ sky130_fd_sc_hd__buf_4
XFILLER_0_189_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31914_ _04425_ net120 VGND VGND VPWR VPWR datamem.rd_data_mem\[19\] sky130_fd_sc_hd__dlxtn_1
X_16848_ _04672_ VGND VGND VPWR VPWR _01614_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_192_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32894_ clknet_leaf_158_clk _04316_ VGND VGND VPWR VPWR datamem.data_ram\[10\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_195_Right_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_205_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_220_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31845_ clknet_leaf_157_clk _03299_ VGND VGND VPWR VPWR datamem.data_ram\[8\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_19567_ _06829_ VGND VGND VPWR VPWR _06863_ sky130_fd_sc_hd__buf_8
XFILLER_0_215_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16779_ net3455 _14466_ _04634_ VGND VGND VPWR VPWR _04636_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18518_ _05370_ _05719_ _05820_ VGND VGND VPWR VPWR _05879_ sky130_fd_sc_hd__and3_1
X_19498_ datamem.data_ram\[27\]\[16\] _06636_ _06788_ _06793_ VGND VGND VPWR VPWR
+ _06794_ sky130_fd_sc_hd__o211a_1
XFILLER_0_73_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31776_ clknet_leaf_272_clk _03230_ VGND VGND VPWR VPWR datamem.data_ram\[6\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_174_4661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_4672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_4683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18449_ rvcpu.dp.plde.ALUControlE\[0\] _00003_ VGND VGND VPWR VPWR _05812_ sky130_fd_sc_hd__or2_1
X_30727_ clknet_leaf_196_clk _02462_ VGND VGND VPWR VPWR datamem.data_ram\[48\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23890__450 clknet_1_0__leaf__10222_ VGND VGND VPWR VPWR net576 sky130_fd_sc_hd__inv_2
XFILLER_0_200_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21460_ rvcpu.dp.rf.reg_file_arr\[8\]\[4\] rvcpu.dp.rf.reg_file_arr\[10\]\[4\] rvcpu.dp.rf.reg_file_arr\[9\]\[4\]
+ rvcpu.dp.rf.reg_file_arr\[11\]\[4\] _08649_ _08537_ VGND VGND VPWR VPWR _08718_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_170_4569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30658_ clknet_leaf_216_clk _02393_ VGND VGND VPWR VPWR datamem.data_ram\[50\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20411_ datamem.data_ram\[62\]\[12\] _06744_ _07243_ datamem.data_ram\[57\]\[12\]
+ VGND VGND VPWR VPWR _07703_ sky130_fd_sc_hd__o22a_1
XFILLER_0_114_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21391_ _08558_ VGND VGND VPWR VPWR _08652_ sky130_fd_sc_hd__buf_2
X_30589_ clknet_leaf_117_clk _02324_ VGND VGND VPWR VPWR datamem.data_ram\[53\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_226_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20342_ datamem.data_ram\[62\]\[4\] _06978_ _06948_ datamem.data_ram\[57\]\[4\] VGND
+ VGND VPWR VPWR _07634_ sky130_fd_sc_hd__a22o_1
XFILLER_0_160_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32328_ clknet_leaf_170_clk _03750_ VGND VGND VPWR VPWR datamem.data_ram\[31\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_133_3690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20273_ datamem.data_ram\[37\]\[19\] _06724_ _07564_ _07565_ VGND VGND VPWR VPWR
+ _07566_ sky130_fd_sc_hd__o211a_1
X_32259_ clknet_leaf_243_clk _03681_ VGND VGND VPWR VPWR datamem.data_ram\[34\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_73_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24066__593 clknet_1_0__leaf__10247_ VGND VGND VPWR VPWR net719 sky130_fd_sc_hd__inv_2
XFILLER_0_102_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_73_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22012_ _09239_ VGND VGND VPWR VPWR _09240_ sky130_fd_sc_hd__clkbuf_2
Xhold3201 rvcpu.dp.rf.reg_file_arr\[31\]\[28\] VGND VGND VPWR VPWR net4351 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3212 rvcpu.dp.rf.reg_file_arr\[23\]\[27\] VGND VGND VPWR VPWR net4362 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3223 datamem.data_ram\[59\]\[16\] VGND VGND VPWR VPWR net4373 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3234 rvcpu.dp.rf.reg_file_arr\[24\]\[18\] VGND VGND VPWR VPWR net4384 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2500 datamem.data_ram\[42\]\[12\] VGND VGND VPWR VPWR net3650 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3245 rvcpu.dp.rf.reg_file_arr\[29\]\[28\] VGND VGND VPWR VPWR net4395 sky130_fd_sc_hd__dlygate4sd3_1
X_26820_ _11679_ _11774_ VGND VGND VPWR VPWR _11776_ sky130_fd_sc_hd__and2_1
Xhold3256 datamem.data_ram\[55\]\[19\] VGND VGND VPWR VPWR net4406 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2511 datamem.data_ram\[27\]\[24\] VGND VGND VPWR VPWR net3661 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2522 datamem.data_ram\[51\]\[28\] VGND VGND VPWR VPWR net3672 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3267 datamem.data_ram\[1\]\[14\] VGND VGND VPWR VPWR net4417 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2533 datamem.data_ram\[50\]\[19\] VGND VGND VPWR VPWR net3683 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3278 rvcpu.dp.rf.reg_file_arr\[21\]\[22\] VGND VGND VPWR VPWR net4428 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_880 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_3904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3289 rvcpu.dp.rf.reg_file_arr\[24\]\[26\] VGND VGND VPWR VPWR net4439 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2544 rvcpu.dp.rf.reg_file_arr\[28\]\[14\] VGND VGND VPWR VPWR net3694 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2555 datamem.data_ram\[26\]\[18\] VGND VGND VPWR VPWR net3705 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1810 datamem.data_ram\[49\]\[8\] VGND VGND VPWR VPWR net2960 sky130_fd_sc_hd__dlygate4sd3_1
X_26751_ _11700_ net1818 _11724_ _11733_ VGND VGND VPWR VPWR _03307_ sky130_fd_sc_hd__a31o_1
Xhold2566 datamem.data_ram\[13\]\[27\] VGND VGND VPWR VPWR net3716 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1821 datamem.data_ram\[55\]\[27\] VGND VGND VPWR VPWR net2971 sky130_fd_sc_hd__dlygate4sd3_1
X_23963_ _10235_ VGND VGND VPWR VPWR _02017_ sky130_fd_sc_hd__clkbuf_1
Xhold2577 datamem.data_ram\[3\]\[17\] VGND VGND VPWR VPWR net3727 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1832 datamem.data_ram\[14\]\[13\] VGND VGND VPWR VPWR net2982 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1843 datamem.data_ram\[50\]\[18\] VGND VGND VPWR VPWR net2993 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2588 datamem.data_ram\[54\]\[8\] VGND VGND VPWR VPWR net3738 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_95_clk clknet_5_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_95_clk sky130_fd_sc_hd__clkbuf_8
Xhold1854 datamem.data_ram\[37\]\[26\] VGND VGND VPWR VPWR net3004 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2599 datamem.data_ram\[46\]\[20\] VGND VGND VPWR VPWR net3749 sky130_fd_sc_hd__dlygate4sd3_1
X_25702_ _10542_ _11123_ _10998_ VGND VGND VPWR VPWR _11124_ sky130_fd_sc_hd__a21oi_4
X_22914_ _10047_ VGND VGND VPWR VPWR _10048_ sky130_fd_sc_hd__buf_2
Xhold1865 datamem.data_ram\[29\]\[24\] VGND VGND VPWR VPWR net3015 sky130_fd_sc_hd__dlygate4sd3_1
X_29470_ net832 _01205_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[2\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_26682_ _11676_ _11694_ VGND VGND VPWR VPWR _11695_ sky130_fd_sc_hd__and2_1
Xhold1876 rvcpu.dp.rf.reg_file_arr\[24\]\[13\] VGND VGND VPWR VPWR net3026 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1887 rvcpu.dp.rf.reg_file_arr\[18\]\[31\] VGND VGND VPWR VPWR net3037 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_162_Right_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1898 datamem.data_ram\[9\]\[11\] VGND VGND VPWR VPWR net3048 sky130_fd_sc_hd__dlygate4sd3_1
X_28421_ _09350_ _12602_ _12668_ VGND VGND VPWR VPWR _12688_ sky130_fd_sc_hd__a21oi_4
X_25633_ _11057_ net1488 _11077_ _11084_ VGND VGND VPWR VPWR _02838_ sky130_fd_sc_hd__a31o_1
XFILLER_0_116_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22845_ rvcpu.dp.rf.reg_file_arr\[12\]\[28\] rvcpu.dp.rf.reg_file_arr\[13\]\[28\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[28\] rvcpu.dp.rf.reg_file_arr\[15\]\[28\] _09464_
+ _09467_ VGND VGND VPWR VPWR _09983_ sky130_fd_sc_hd__mux4_1
X_23365__1001 clknet_1_0__leaf__10138_ VGND VGND VPWR VPWR net1127 sky130_fd_sc_hd__inv_2
XFILLER_0_196_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28352_ _12447_ net4140 net95 VGND VGND VPWR VPWR _12651_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25564_ _10946_ _11039_ VGND VGND VPWR VPWR _11042_ sky130_fd_sc_hd__nor2_2
XFILLER_0_112_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_588 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22776_ _09705_ _09909_ _09913_ _09917_ VGND VGND VPWR VPWR _09918_ sky130_fd_sc_hd__and4_1
XFILLER_0_195_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27303_ _10209_ _08066_ _11898_ VGND VGND VPWR VPWR _12066_ sky130_fd_sc_hd__and3_1
XFILLER_0_149_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24515_ _10451_ VGND VGND VPWR VPWR _02353_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28283_ _12430_ net3081 _12613_ VGND VGND VPWR VPWR _12614_ sky130_fd_sc_hd__mux2_1
X_21727_ _08969_ _08970_ _08743_ VGND VGND VPWR VPWR _08971_ sky130_fd_sc_hd__mux2_2
XFILLER_0_137_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25495_ _11002_ VGND VGND VPWR VPWR _02782_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23140__815 clknet_1_0__leaf__10107_ VGND VGND VPWR VPWR net941 sky130_fd_sc_hd__inv_2
XFILLER_0_191_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27234_ _07808_ _10043_ _10897_ VGND VGND VPWR VPWR _12029_ sky130_fd_sc_hd__or3_1
XFILLER_0_192_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24446_ _10060_ VGND VGND VPWR VPWR _10410_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_164_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21658_ _08904_ _08905_ _08540_ VGND VGND VPWR VPWR _08906_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27165_ _11974_ net1674 _11983_ _11988_ VGND VGND VPWR VPWR _03466_ sky130_fd_sc_hd__a31o_1
X_20609_ datamem.data_ram\[47\]\[13\] _06784_ _06790_ datamem.data_ram\[41\]\[13\]
+ _07899_ VGND VGND VPWR VPWR _07900_ sky130_fd_sc_hd__o221a_1
XFILLER_0_151_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24377_ _09226_ _10337_ _10366_ VGND VGND VPWR VPWR _10367_ sky130_fd_sc_hd__a21oi_4
X_21589_ rvcpu.dp.rf.reg_file_arr\[12\]\[10\] rvcpu.dp.rf.reg_file_arr\[13\]\[10\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[10\] rvcpu.dp.rf.reg_file_arr\[15\]\[10\] _08839_
+ _08840_ VGND VGND VPWR VPWR _08841_ sky130_fd_sc_hd__mux4_1
XFILLER_0_201_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23255__902 clknet_1_0__leaf__10127_ VGND VGND VPWR VPWR net1028 sky130_fd_sc_hd__inv_2
X_26116_ _11393_ VGND VGND VPWR VPWR _03011_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27096_ _11938_ net1664 _11940_ _11944_ VGND VGND VPWR VPWR _03441_ sky130_fd_sc_hd__a31o_1
XFILLER_0_22_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26047_ _11078_ _11351_ VGND VGND VPWR VPWR _11352_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17820_ rvcpu.dp.plem.ALUResultM\[26\] _05207_ _05178_ VGND VGND VPWR VPWR _05208_
+ sky130_fd_sc_hd__mux2_1
X_29806_ net1144 _01541_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[1\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27998_ _12459_ VGND VGND VPWR VPWR _03828_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_17 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17751_ _13275_ net2743 _05117_ VGND VGND VPWR VPWR _05151_ sky130_fd_sc_hd__mux2_1
X_26949_ _11849_ net1497 _11853_ _11856_ VGND VGND VPWR VPWR _03382_ sky130_fd_sc_hd__a31o_1
X_14963_ _13304_ _13335_ _13348_ VGND VGND VPWR VPWR _13512_ sky130_fd_sc_hd__and3_1
Xhold6 rvcpu.dp.plem.lAuiPCM\[24\] VGND VGND VPWR VPWR net1156 sky130_fd_sc_hd__dlygate4sd3_1
X_29737_ net1083 _01472_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[21\]\[4\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_86_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_86_clk sky130_fd_sc_hd__clkbuf_8
X_16702_ _14166_ net4305 _04587_ VGND VGND VPWR VPWR _04595_ sky130_fd_sc_hd__mux2_1
XFILLER_0_226_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29668_ net1014 _01403_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[24\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_17682_ _05114_ VGND VGND VPWR VPWR _01198_ sky130_fd_sc_hd__clkbuf_1
X_14894_ _13442_ _13444_ VGND VGND VPWR VPWR _13445_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19421_ _06625_ VGND VGND VPWR VPWR _06717_ sky130_fd_sc_hd__buf_6
XFILLER_0_226_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28619_ _12751_ net3914 _12805_ VGND VGND VPWR VPWR _12806_ sky130_fd_sc_hd__mux2_1
X_16633_ _04558_ VGND VGND VPWR VPWR _01723_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29599_ net953 _01334_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[25\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31630_ clknet_leaf_48_clk net1242 VGND VGND VPWR VPWR rvcpu.dp.plmw.lAuiPCW\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_19352_ _06647_ VGND VGND VPWR VPWR _06648_ sky130_fd_sc_hd__clkbuf_8
X_16564_ _04521_ VGND VGND VPWR VPWR _01763_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18303_ _05667_ VGND VGND VPWR VPWR _05668_ sky130_fd_sc_hd__clkbuf_4
X_15515_ _13542_ _13531_ _13698_ _13648_ _14021_ VGND VGND VPWR VPWR _14042_ sky130_fd_sc_hd__o32a_1
XFILLER_0_155_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31561_ clknet_leaf_62_clk datamem.rd_data_mem\[11\] VGND VGND VPWR VPWR rvcpu.dp.plmw.ReadDataW\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_19283_ _06570_ _06575_ _06574_ _06567_ VGND VGND VPWR VPWR _04450_ sky130_fd_sc_hd__o211a_1
X_16495_ net2250 _14455_ _04478_ VGND VGND VPWR VPWR _04485_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_216_5690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18234_ _05346_ _05356_ _05589_ _05598_ VGND VGND VPWR VPWR _05599_ sky130_fd_sc_hd__o31ai_4
X_30512_ clknet_leaf_203_clk _02247_ VGND VGND VPWR VPWR datamem.data_ram\[56\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_15446_ _13561_ _13656_ _13353_ VGND VGND VPWR VPWR _13977_ sky130_fd_sc_hd__o21ai_1
X_31492_ clknet_leaf_46_clk rvcpu.dp.lAuiPCE\[18\] VGND VGND VPWR VPWR rvcpu.dp.plem.lAuiPCM\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_212_5576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_212_5587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18165_ _05527_ _05528_ VGND VGND VPWR VPWR _05530_ sky130_fd_sc_hd__nor2_1
X_30443_ net781 _02178_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[29\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_15377_ _13359_ _13474_ _13634_ _13910_ _13409_ VGND VGND VPWR VPWR _13911_ sky130_fd_sc_hd__o311a_1
XFILLER_0_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17116_ _04814_ VGND VGND VPWR VPWR _01480_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap103 _05408_ VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_64_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18096_ rvcpu.dp.plde.ImmExtE\[22\] rvcpu.dp.SrcBFW_Mux.y\[22\] _05279_ VGND VGND
+ VPWR VPWR _05464_ sky130_fd_sc_hd__mux2_1
Xmax_cap114 net115 VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_68_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30374_ net720 _02109_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[3\]\[25\] sky130_fd_sc_hd__dfxtp_1
Xhold406 datamem.data_ram\[23\]\[1\] VGND VGND VPWR VPWR net1556 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold417 datamem.data_ram\[4\]\[5\] VGND VGND VPWR VPWR net1567 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_225_5904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold428 datamem.data_ram\[29\]\[1\] VGND VGND VPWR VPWR net1578 sky130_fd_sc_hd__dlygate4sd3_1
X_32113_ clknet_leaf_98_clk _03535_ VGND VGND VPWR VPWR datamem.data_ram\[0\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold439 datamem.data_ram\[22\]\[3\] VGND VGND VPWR VPWR net1589 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17047_ net2196 _14461_ _04768_ VGND VGND VPWR VPWR _04778_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_4004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22978__685 clknet_1_0__leaf__10083_ VGND VGND VPWR VPWR net811 sky130_fd_sc_hd__inv_2
X_32044_ clknet_leaf_132_clk _03466_ VGND VGND VPWR VPWR datamem.data_ram\[49\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18998_ _06315_ _06327_ _06332_ VGND VGND VPWR VPWR _06333_ sky130_fd_sc_hd__or3_1
Xhold1106 datamem.data_ram\[35\]\[23\] VGND VGND VPWR VPWR net2256 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1117 datamem.data_ram\[14\]\[15\] VGND VGND VPWR VPWR net2267 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1128 datamem.data_ram\[32\]\[13\] VGND VGND VPWR VPWR net2278 sky130_fd_sc_hd__dlygate4sd3_1
X_17949_ rvcpu.dp.plde.ALUSrcE VGND VGND VPWR VPWR _05321_ sky130_fd_sc_hd__buf_4
XFILLER_0_139_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_77_clk clknet_5_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_77_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_105_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1139 rvcpu.dp.rf.reg_file_arr\[7\]\[5\] VGND VGND VPWR VPWR net2289 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20960_ datamem.data_ram\[58\]\[15\] _06608_ _06917_ _08248_ VGND VGND VPWR VPWR
+ _08249_ sky130_fd_sc_hd__o22a_1
X_32946_ clknet_leaf_211_clk _04368_ VGND VGND VPWR VPWR datamem.data_ram\[6\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_176_4712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_177_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_176_4723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19619_ _06914_ VGND VGND VPWR VPWR _06915_ sky130_fd_sc_hd__buf_2
XFILLER_0_71_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20891_ _08166_ _08180_ _06985_ VGND VGND VPWR VPWR _08181_ sky130_fd_sc_hd__a21o_1
XFILLER_0_45_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32877_ clknet_leaf_54_clk _04299_ VGND VGND VPWR VPWR datamem.data_ram\[10\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22630_ _09511_ _09778_ VGND VGND VPWR VPWR _09779_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31828_ clknet_leaf_105_clk _03282_ VGND VGND VPWR VPWR datamem.data_ram\[16\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22561_ _09416_ VGND VGND VPWR VPWR _09714_ sky130_fd_sc_hd__buf_4
X_31759_ clknet_leaf_105_clk _03213_ VGND VGND VPWR VPWR datamem.data_ram\[18\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_23736__327 clknet_1_1__leaf__10199_ VGND VGND VPWR VPWR net453 sky130_fd_sc_hd__inv_2
XFILLER_0_174_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21512_ _08627_ _08762_ _08764_ _08766_ VGND VGND VPWR VPWR _08767_ sky130_fd_sc_hd__o2bb2a_1
X_24300_ _10323_ VGND VGND VPWR VPWR _02266_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_3730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25280_ _10882_ VGND VGND VPWR VPWR _02687_ sky130_fd_sc_hd__clkbuf_1
X_22492_ rvcpu.dp.rf.reg_file_arr\[0\]\[9\] rvcpu.dp.rf.reg_file_arr\[1\]\[9\] rvcpu.dp.rf.reg_file_arr\[2\]\[9\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[9\] _09477_ _09383_ VGND VGND VPWR VPWR _09649_ sky130_fd_sc_hd__mux4_1
XFILLER_0_111_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_3741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24231_ _10286_ VGND VGND VPWR VPWR _02234_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_161_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21443_ _08672_ _08681_ _08691_ _08701_ VGND VGND VPWR VPWR _08702_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_25_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_3638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24162_ clknet_1_1__leaf__10079_ VGND VGND VPWR VPWR _10264_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_131_3649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21374_ _08559_ VGND VGND VPWR VPWR _08635_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_96_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_1172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20325_ datamem.data_ram\[22\]\[4\] _07159_ _07081_ _07616_ VGND VGND VPWR VPWR _07617_
+ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_9_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28970_ _12727_ net1750 _12988_ _12993_ VGND VGND VPWR VPWR _04266_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_9_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold940 rvcpu.dp.rf.reg_file_arr\[5\]\[9\] VGND VGND VPWR VPWR net2090 sky130_fd_sc_hd__dlygate4sd3_1
Xhold951 datamem.data_ram\[9\]\[25\] VGND VGND VPWR VPWR net2101 sky130_fd_sc_hd__dlygate4sd3_1
X_27921_ _10777_ _10114_ _12356_ VGND VGND VPWR VPWR _12412_ sky130_fd_sc_hd__a21oi_4
Xhold962 rvcpu.dp.rf.reg_file_arr\[25\]\[19\] VGND VGND VPWR VPWR net2112 sky130_fd_sc_hd__dlygate4sd3_1
X_23044_ clknet_1_1__leaf__10087_ VGND VGND VPWR VPWR _10090_ sky130_fd_sc_hd__buf_1
X_20256_ _06680_ _07546_ _07548_ VGND VGND VPWR VPWR _07549_ sky130_fd_sc_hd__or3_2
Xhold973 rvcpu.dp.rf.reg_file_arr\[5\]\[18\] VGND VGND VPWR VPWR net2123 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold984 rvcpu.dp.rf.reg_file_arr\[30\]\[22\] VGND VGND VPWR VPWR net2134 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3020 rvcpu.dp.rf.reg_file_arr\[22\]\[17\] VGND VGND VPWR VPWR net4170 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_34_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold995 rvcpu.dp.rf.reg_file_arr\[4\]\[18\] VGND VGND VPWR VPWR net2145 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_34_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3031 datamem.data_ram\[47\]\[12\] VGND VGND VPWR VPWR net4181 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold3042 rvcpu.dp.rf.reg_file_arr\[16\]\[26\] VGND VGND VPWR VPWR net4192 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27852_ _12374_ VGND VGND VPWR VPWR _03767_ sky130_fd_sc_hd__clkbuf_1
Xhold3053 datamem.data_ram\[31\]\[21\] VGND VGND VPWR VPWR net4203 sky130_fd_sc_hd__dlygate4sd3_1
X_20187_ datamem.data_ram\[2\]\[11\] _06692_ _07031_ _07479_ VGND VGND VPWR VPWR _07480_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_216_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3064 datamem.data_ram\[53\]\[20\] VGND VGND VPWR VPWR net4214 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2330 datamem.data_ram\[63\]\[9\] VGND VGND VPWR VPWR net3480 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3075 datamem.data_ram\[8\]\[31\] VGND VGND VPWR VPWR net4225 sky130_fd_sc_hd__dlygate4sd3_1
X_26803_ _11753_ net1577 _11761_ _11765_ VGND VGND VPWR VPWR _03327_ sky130_fd_sc_hd__a31o_1
Xhold3086 datamem.data_ram\[55\]\[17\] VGND VGND VPWR VPWR net4236 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2341 datamem.data_ram\[13\]\[24\] VGND VGND VPWR VPWR net3491 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2352 datamem.data_ram\[23\]\[19\] VGND VGND VPWR VPWR net3502 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3097 datamem.data_ram\[25\]\[14\] VGND VGND VPWR VPWR net4247 sky130_fd_sc_hd__dlygate4sd3_1
X_27783_ _12332_ VGND VGND VPWR VPWR _03740_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24995_ _10718_ VGND VGND VPWR VPWR _02566_ sky130_fd_sc_hd__clkbuf_1
Xhold2363 datamem.data_ram\[50\]\[26\] VGND VGND VPWR VPWR net3513 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_68_clk clknet_5_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_68_clk sky130_fd_sc_hd__clkbuf_8
X_23285__928 clknet_1_1__leaf__10131_ VGND VGND VPWR VPWR net1054 sky130_fd_sc_hd__inv_2
Xhold2374 rvcpu.dp.rf.reg_file_arr\[22\]\[31\] VGND VGND VPWR VPWR net3524 sky130_fd_sc_hd__dlygate4sd3_1
X_29522_ net884 _01257_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[28\]\[29\] sky130_fd_sc_hd__dfxtp_1
Xhold2385 datamem.data_ram\[17\]\[29\] VGND VGND VPWR VPWR net3535 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1640 datamem.data_ram\[28\]\[9\] VGND VGND VPWR VPWR net2790 sky130_fd_sc_hd__dlygate4sd3_1
X_26734_ _09227_ _11603_ VGND VGND VPWR VPWR _11723_ sky130_fd_sc_hd__or2_1
Xhold2396 datamem.data_ram\[45\]\[19\] VGND VGND VPWR VPWR net3546 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1651 datamem.data_ram\[31\]\[13\] VGND VGND VPWR VPWR net2801 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1662 datamem.data_ram\[59\]\[29\] VGND VGND VPWR VPWR net2812 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1673 rvcpu.dp.rf.reg_file_arr\[17\]\[10\] VGND VGND VPWR VPWR net2823 sky130_fd_sc_hd__dlygate4sd3_1
X_23897__456 clknet_1_0__leaf__10223_ VGND VGND VPWR VPWR net582 sky130_fd_sc_hd__inv_2
XFILLER_0_193_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1684 rvcpu.dp.rf.reg_file_arr\[25\]\[7\] VGND VGND VPWR VPWR net2834 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1695 rvcpu.dp.rf.reg_file_arr\[30\]\[13\] VGND VGND VPWR VPWR net2845 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29453_ net815 _01188_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[30\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_26665_ _11104_ VGND VGND VPWR VPWR _11683_ sky130_fd_sc_hd__buf_2
XFILLER_0_98_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24116__623 clknet_1_1__leaf__10259_ VGND VGND VPWR VPWR net749 sky130_fd_sc_hd__inv_2
X_28404_ _12447_ net2774 _12678_ VGND VGND VPWR VPWR _12679_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0__10265_ _10265_ VGND VGND VPWR VPWR clknet_0__10265_ sky130_fd_sc_hd__clkbuf_16
X_25616_ _11072_ VGND VGND VPWR VPWR _02833_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_169_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22828_ _09481_ _09966_ VGND VGND VPWR VPWR _09967_ sky130_fd_sc_hd__and2_1
X_29384_ clknet_leaf_266_clk _01119_ VGND VGND VPWR VPWR datamem.data_ram\[60\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_26596_ _10066_ VGND VGND VPWR VPWR _11645_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_39_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_183_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28335_ _12430_ net2623 _12641_ VGND VGND VPWR VPWR _12642_ sky130_fd_sc_hd__mux2_1
X_25547_ _10754_ net3811 _11030_ VGND VGND VPWR VPWR _11032_ sky130_fd_sc_hd__mux2_1
Xclkbuf_0__10196_ _10196_ VGND VGND VPWR VPWR clknet_0__10196_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_94_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22759_ _09901_ VGND VGND VPWR VPWR _01147_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15300_ _13449_ _13389_ _13509_ _13763_ VGND VGND VPWR VPWR _13838_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28266_ _12604_ VGND VGND VPWR VPWR _03951_ sky130_fd_sc_hd__clkbuf_1
X_16280_ _14502_ VGND VGND VPWR VPWR _01896_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25478_ _10780_ net35 VGND VGND VPWR VPWR _10996_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_229_6004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_229_6015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_229_6026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27217_ _11965_ _12019_ VGND VGND VPWR VPWR _12020_ sky130_fd_sc_hd__and2_1
X_15231_ _13360_ _13771_ _13315_ VGND VGND VPWR VPWR _13772_ sky130_fd_sc_hd__a21o_1
XFILLER_0_129_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24429_ _10397_ VGND VGND VPWR VPWR _02321_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28197_ _12566_ VGND VGND VPWR VPWR _03920_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27148_ _11974_ net1643 _11964_ _11977_ VGND VGND VPWR VPWR _03460_ sky130_fd_sc_hd__a31o_1
X_15162_ _13475_ VGND VGND VPWR VPWR _13706_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_151_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27079_ _11919_ net1735 _11923_ _11932_ VGND VGND VPWR VPWR _03436_ sky130_fd_sc_hd__a31o_1
X_15093_ _13521_ VGND VGND VPWR VPWR _13638_ sky130_fd_sc_hd__clkbuf_4
X_19970_ datamem.data_ram\[30\]\[18\] _06763_ _06782_ datamem.data_ram\[25\]\[18\]
+ VGND VGND VPWR VPWR _07264_ sky130_fd_sc_hd__o22a_1
XFILLER_0_26_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18921_ _05535_ _06108_ _06136_ _06001_ VGND VGND VPWR VPWR _06261_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_31_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30090_ net452 _01825_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[11\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18852_ _05275_ _06031_ _05944_ _05819_ VGND VGND VPWR VPWR _06196_ sky130_fd_sc_hd__a31o_1
XFILLER_0_219_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17803_ _05195_ VGND VGND VPWR VPWR _05196_ sky130_fd_sc_hd__clkbuf_4
X_18783_ _06131_ VGND VGND VPWR VPWR rvcpu.ALUResultE\[15\] sky130_fd_sc_hd__clkbuf_1
X_15995_ _14335_ VGND VGND VPWR VPWR _02030_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_59_clk clknet_5_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_59_clk sky130_fd_sc_hd__clkbuf_8
X_17734_ _05142_ VGND VGND VPWR VPWR _01174_ sky130_fd_sc_hd__clkbuf_1
X_32800_ clknet_leaf_186_clk _04222_ VGND VGND VPWR VPWR datamem.data_ram\[13\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_14946_ _13401_ _13494_ VGND VGND VPWR VPWR _13495_ sky130_fd_sc_hd__nor2_1
X_30992_ clknet_leaf_102_clk _02727_ VGND VGND VPWR VPWR datamem.data_ram\[13\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_216_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32731_ clknet_leaf_171_clk _04153_ VGND VGND VPWR VPWR datamem.data_ram\[16\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_17665_ net1972 _13247_ _05104_ VGND VGND VPWR VPWR _05106_ sky130_fd_sc_hd__mux2_1
X_14877_ _13428_ VGND VGND VPWR VPWR _13429_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_106_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_218_5730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16616_ _04549_ VGND VGND VPWR VPWR _01731_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19404_ _06699_ VGND VGND VPWR VPWR _06700_ sky130_fd_sc_hd__buf_6
XFILLER_0_203_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_202_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32662_ clknet_leaf_83_clk _04084_ VGND VGND VPWR VPWR datamem.data_ram\[19\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_212_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_203_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17596_ _05069_ VGND VGND VPWR VPWR _01239_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_214_5627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31613_ clknet_leaf_26_clk net1212 VGND VGND VPWR VPWR rvcpu.dp.plmw.PCPlus4W\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_214_5638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16547_ _04512_ VGND VGND VPWR VPWR _01771_ sky130_fd_sc_hd__clkbuf_1
X_19335_ net122 _06607_ VGND VGND VPWR VPWR _06631_ sky130_fd_sc_hd__nand2_8
X_32593_ clknet_leaf_252_clk _04015_ VGND VGND VPWR VPWR datamem.data_ram\[21\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_222_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19266_ rvcpu.dp.plfd.InstrD\[3\] rvcpu.dp.plfd.InstrD\[2\] rvcpu.dp.plfd.InstrD\[0\]
+ VGND VGND VPWR VPWR _06566_ sky130_fd_sc_hd__or3b_1
X_31544_ clknet_leaf_15_clk net1278 VGND VGND VPWR VPWR rvcpu.dp.plem.RdM\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16478_ net3234 _14438_ _04467_ VGND VGND VPWR VPWR _04476_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18217_ _05577_ _05581_ _05383_ VGND VGND VPWR VPWR _05582_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15429_ _13858_ _13959_ _13423_ VGND VGND VPWR VPWR _13960_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31475_ clknet_leaf_66_clk rvcpu.dp.lAuiPCE\[1\] VGND VGND VPWR VPWR rvcpu.dp.plem.lAuiPCM\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_19197_ rvcpu.dp.plde.ImmExtE\[23\] rvcpu.dp.plde.PCE\[23\] VGND VGND VPWR VPWR _06507_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_182_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18148_ _05512_ VGND VGND VPWR VPWR _05513_ sky130_fd_sc_hd__buf_2
X_30426_ net764 _02161_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[29\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_47 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold203 datamem.data_ram\[30\]\[6\] VGND VGND VPWR VPWR net1353 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold214 rvcpu.dp.pcreg.q\[1\] VGND VGND VPWR VPWR net1364 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_169_4560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold225 datamem.data_ram\[40\]\[6\] VGND VGND VPWR VPWR net1375 sky130_fd_sc_hd__dlygate4sd3_1
X_18079_ _05446_ _05409_ VGND VGND VPWR VPWR _05447_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30357_ net703 _02092_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[3\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_223_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold236 datamem.data_ram\[29\]\[6\] VGND VGND VPWR VPWR net1386 sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 datamem.data_ram\[27\]\[6\] VGND VGND VPWR VPWR net1397 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold258 datamem.data_ram\[14\]\[1\] VGND VGND VPWR VPWR net1408 sky130_fd_sc_hd__dlygate4sd3_1
X_20110_ datamem.data_ram\[21\]\[10\] _06723_ _07402_ _07403_ VGND VGND VPWR VPWR
+ _07404_ sky130_fd_sc_hd__o211a_1
X_23364__1000 clknet_1_0__leaf__10138_ VGND VGND VPWR VPWR net1126 sky130_fd_sc_hd__inv_2
Xhold269 datamem.data_ram\[38\]\[0\] VGND VGND VPWR VPWR net1419 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_165_4446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21090_ datamem.data_ram\[54\]\[7\] _06950_ _06946_ datamem.data_ram\[49\]\[7\] _08378_
+ VGND VGND VPWR VPWR _08379_ sky130_fd_sc_hd__a221o_1
XFILLER_0_229_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_165_4457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30288_ net634 _02023_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[5\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32027_ clknet_leaf_127_clk _03449_ VGND VGND VPWR VPWR datamem.data_ram\[26\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_20041_ datamem.data_ram\[0\]\[26\] _06645_ _07242_ datamem.data_ram\[1\]\[26\] VGND
+ VGND VPWR VPWR _07335_ sky130_fd_sc_hd__o22a_1
XFILLER_0_42_1164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_13_Left_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23800_ clknet_1_0__leaf__10203_ VGND VGND VPWR VPWR _10206_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_68_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_68_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_307 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24780_ _10598_ _10601_ _10501_ VGND VGND VPWR VPWR _10602_ sky130_fd_sc_hd__a21oi_1
X_21992_ rvcpu.dp.plem.WriteDataM\[16\] _09221_ VGND VGND VPWR VPWR _09222_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_124_3464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_3475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20943_ datamem.data_ram\[63\]\[22\] _07860_ _07863_ datamem.data_ram\[61\]\[22\]
+ _08232_ VGND VGND VPWR VPWR _08233_ sky130_fd_sc_hd__o221a_1
X_32929_ clknet_leaf_142_clk _04351_ VGND VGND VPWR VPWR datamem.data_ram\[7\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_109 _07031_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26450_ net1867 _11573_ _11578_ _11570_ VGND VGND VPWR VPWR _03161_ sky130_fd_sc_hd__o211a_1
X_20874_ datamem.data_ram\[48\]\[14\] _06647_ _06790_ datamem.data_ram\[49\]\[14\]
+ VGND VGND VPWR VPWR _08164_ sky130_fd_sc_hd__o22a_1
X_23970__506 clknet_1_0__leaf__10238_ VGND VGND VPWR VPWR net632 sky130_fd_sc_hd__inv_2
XFILLER_0_7_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_178_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25401_ _10954_ net1589 _10949_ _10955_ VGND VGND VPWR VPWR _02735_ sky130_fd_sc_hd__a31o_1
XFILLER_0_138_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22613_ _09516_ _09762_ VGND VGND VPWR VPWR _09763_ sky130_fd_sc_hd__or2_1
X_26381_ _11524_ rvcpu.ALUResultE\[3\] _06371_ _11522_ VGND VGND VPWR VPWR _11528_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_27_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28120_ _12525_ VGND VGND VPWR VPWR _03884_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_22_Left_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_187_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25332_ _10756_ net3405 _10909_ VGND VGND VPWR VPWR _10912_ sky130_fd_sc_hd__mux2_1
X_22544_ _09528_ _09697_ _09426_ VGND VGND VPWR VPWR _09698_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28051_ _12458_ net3619 net96 VGND VGND VPWR VPWR _12489_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_98_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25263_ _10067_ _10868_ VGND VGND VPWR VPWR _10873_ sky130_fd_sc_hd__and2_1
XFILLER_0_173_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22475_ _09632_ VGND VGND VPWR VPWR _01132_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27002_ _11822_ _11886_ VGND VGND VPWR VPWR _11887_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24214_ _10277_ VGND VGND VPWR VPWR _02226_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21426_ rvcpu.dp.rf.reg_file_arr\[0\]\[3\] rvcpu.dp.rf.reg_file_arr\[1\]\[3\] rvcpu.dp.rf.reg_file_arr\[2\]\[3\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[3\] _08683_ _08684_ VGND VGND VPWR VPWR _08685_ sky130_fd_sc_hd__mux4_1
XFILLER_0_133_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25194_ _10735_ net3901 net57 VGND VGND VPWR VPWR _10835_ sky130_fd_sc_hd__mux2_1
X_21357_ _08611_ _08613_ _08614_ _08618_ VGND VGND VPWR VPWR _08619_ sky130_fd_sc_hd__o211a_1
X_20308_ datamem.data_ram\[7\]\[4\] _06927_ _07133_ datamem.data_ram\[1\]\[4\] VGND
+ VGND VPWR VPWR _07600_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_57_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28953_ _12983_ VGND VGND VPWR VPWR _04259_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_57_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24076_ _09267_ net4027 _10249_ VGND VGND VPWR VPWR _10250_ sky130_fd_sc_hd__mux2_1
X_21288_ _08549_ VGND VGND VPWR VPWR _08550_ sky130_fd_sc_hd__buf_4
Xhold770 datamem.data_ram\[50\]\[14\] VGND VGND VPWR VPWR net1920 sky130_fd_sc_hd__dlygate4sd3_1
Xhold781 rvcpu.dp.rf.reg_file_arr\[10\]\[9\] VGND VGND VPWR VPWR net1931 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_31_Left_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold792 rvcpu.dp.rf.reg_file_arr\[5\]\[5\] VGND VGND VPWR VPWR net1942 sky130_fd_sc_hd__dlygate4sd3_1
X_20239_ datamem.data_ram\[53\]\[3\] _06920_ _06937_ datamem.data_ram\[48\]\[3\] _07531_
+ VGND VGND VPWR VPWR _07532_ sky130_fd_sc_hd__a221o_1
X_27904_ _10520_ _10092_ _12356_ VGND VGND VPWR VPWR _12403_ sky130_fd_sc_hd__a21oi_1
X_28884_ _12946_ VGND VGND VPWR VPWR _04227_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_53_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27835_ _09313_ VGND VGND VPWR VPWR _12363_ sky130_fd_sc_hd__clkbuf_2
Xhold2160 rvcpu.dp.rf.reg_file_arr\[4\]\[28\] VGND VGND VPWR VPWR net3310 sky130_fd_sc_hd__dlygate4sd3_1
X_14800_ _13352_ VGND VGND VPWR VPWR _13353_ sky130_fd_sc_hd__buf_2
Xhold2171 datamem.data_ram\[41\]\[24\] VGND VGND VPWR VPWR net3321 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2182 rvcpu.dp.rf.reg_file_arr\[26\]\[12\] VGND VGND VPWR VPWR net3332 sky130_fd_sc_hd__dlygate4sd3_1
X_15780_ _14219_ VGND VGND VPWR VPWR _02137_ sky130_fd_sc_hd__clkbuf_1
X_27766_ _12155_ net3622 _12316_ VGND VGND VPWR VPWR _12323_ sky130_fd_sc_hd__mux2_1
XFILLER_0_188_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2193 datamem.data_ram\[22\]\[31\] VGND VGND VPWR VPWR net3343 sky130_fd_sc_hd__dlygate4sd3_1
X_24978_ _10709_ VGND VGND VPWR VPWR _02558_ sky130_fd_sc_hd__clkbuf_1
Xhold1470 datamem.data_ram\[31\]\[18\] VGND VGND VPWR VPWR net2620 sky130_fd_sc_hd__dlygate4sd3_1
X_23604__224 clknet_1_1__leaf__10178_ VGND VGND VPWR VPWR net350 sky130_fd_sc_hd__inv_2
X_14731_ rvcpu.dp.pcreg.q\[5\] VGND VGND VPWR VPWR _13284_ sky130_fd_sc_hd__buf_4
X_26717_ _10838_ _10960_ _11713_ VGND VGND VPWR VPWR _11714_ sky130_fd_sc_hd__a21oi_4
X_29505_ net867 _01240_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[28\]\[12\] sky130_fd_sc_hd__dfxtp_1
Xhold1481 datamem.data_ram\[39\]\[13\] VGND VGND VPWR VPWR net2631 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1492 rvcpu.dp.rf.reg_file_arr\[22\]\[25\] VGND VGND VPWR VPWR net2642 sky130_fd_sc_hd__dlygate4sd3_1
X_23929_ clknet_1_1__leaf__10224_ VGND VGND VPWR VPWR _10227_ sky130_fd_sc_hd__buf_1
X_27697_ _12286_ VGND VGND VPWR VPWR _03700_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17450_ _14164_ net3250 _04985_ VGND VGND VPWR VPWR _04992_ sky130_fd_sc_hd__mux2_1
X_29436_ net798 _01171_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[30\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_23146__821 clknet_1_0__leaf__10107_ VGND VGND VPWR VPWR net947 sky130_fd_sc_hd__inv_2
X_26648_ _11091_ _11663_ VGND VGND VPWR VPWR _11671_ sky130_fd_sc_hd__and2_1
X_14662_ rvcpu.dp.plmw.ALUResultW\[15\] rvcpu.dp.plmw.ReadDataW\[15\] rvcpu.dp.plmw.PCPlus4W\[15\]
+ rvcpu.dp.plmw.lAuiPCW\[15\] _13168_ _13170_ VGND VGND VPWR VPWR _13231_ sky130_fd_sc_hd__mux4_2
XFILLER_0_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1300 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_40_Left_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16401_ _14566_ VGND VGND VPWR VPWR _01839_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_200_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__10248_ _10248_ VGND VGND VPWR VPWR clknet_0__10248_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_95_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17381_ _04955_ VGND VGND VPWR VPWR _01348_ sky130_fd_sc_hd__clkbuf_1
X_29367_ clknet_leaf_198_clk _01102_ VGND VGND VPWR VPWR datamem.data_ram\[60\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_14593_ rvcpu.dp.plmw.RegWriteW rvcpu.dp.plmw.RdW\[0\] VGND VGND VPWR VPWR _13178_
+ sky130_fd_sc_hd__nand2_2
X_26579_ _10735_ net2463 _11629_ VGND VGND VPWR VPWR _11635_ sky130_fd_sc_hd__mux2_1
X_19120_ _06439_ VGND VGND VPWR VPWR rvcpu.dp.lAuiPCE\[13\] sky130_fd_sc_hd__clkbuf_1
X_28318_ _12355_ net3376 _12632_ VGND VGND VPWR VPWR _12633_ sky130_fd_sc_hd__mux2_1
X_16332_ net2450 _14430_ _14525_ VGND VGND VPWR VPWR _14530_ sky130_fd_sc_hd__mux2_1
XFILLER_0_229_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0__10179_ _10179_ VGND VGND VPWR VPWR clknet_0__10179_ sky130_fd_sc_hd__clkbuf_16
X_29298_ clknet_leaf_1_clk _01033_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD1E\[5\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__10079_ clknet_0__10079_ VGND VGND VPWR VPWR clknet_1_1__leaf__10079_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_82_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19051_ rvcpu.dp.plde.ImmExtE\[4\] rvcpu.dp.plde.PCE\[4\] VGND VGND VPWR VPWR _06379_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_164_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28249_ _12594_ VGND VGND VPWR VPWR _03944_ sky130_fd_sc_hd__clkbuf_1
X_16263_ _14493_ VGND VGND VPWR VPWR _01904_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18002_ _05371_ _05293_ VGND VGND VPWR VPWR _05372_ sky130_fd_sc_hd__nor2_1
X_15214_ _13504_ _13754_ _13755_ _13409_ VGND VGND VPWR VPWR _13756_ sky130_fd_sc_hd__a22o_1
XFILLER_0_180_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31260_ clknet_leaf_15_clk _02963_ VGND VGND VPWR VPWR rvcpu.dp.plfd.InstrD\[18\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_125_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16194_ net2127 _14447_ _14443_ VGND VGND VPWR VPWR _14448_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_498 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30211_ net565 _01946_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[8\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_15145_ _13430_ _13447_ VGND VGND VPWR VPWR _13689_ sky130_fd_sc_hd__nor2_2
X_31191_ clknet_leaf_50_clk _02894_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCPlus4D\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30142_ net504 _01877_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[0\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_15076_ _13509_ _13489_ VGND VGND VPWR VPWR _13622_ sky130_fd_sc_hd__nor2_1
X_19953_ datamem.data_ram\[61\]\[18\] _06663_ _06782_ datamem.data_ram\[57\]\[18\]
+ VGND VGND VPWR VPWR _07247_ sky130_fd_sc_hd__o22a_1
XFILLER_0_227_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_207_5453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_207_5464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_207_5475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18904_ _05461_ _05728_ _06179_ _06244_ VGND VGND VPWR VPWR _06245_ sky130_fd_sc_hd__a211o_1
X_30073_ net435 _01808_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[12\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_19884_ _07154_ _07165_ _07178_ _06988_ VGND VGND VPWR VPWR _07179_ sky130_fd_sc_hd__o211a_1
X_23233__882 clknet_1_1__leaf__10125_ VGND VGND VPWR VPWR net1008 sky130_fd_sc_hd__inv_2
XFILLER_0_219_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_160_4332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18835_ _05889_ _05846_ _06178_ _06180_ VGND VGND VPWR VPWR _06181_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_199_5265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_4343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_208_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_199_5276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18766_ _05334_ _05310_ VGND VGND VPWR VPWR _06116_ sky130_fd_sc_hd__or2_1
XFILLER_0_136_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15978_ _14326_ VGND VGND VPWR VPWR _02038_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14929_ _13432_ _13422_ _13477_ VGND VGND VPWR VPWR _13478_ sky130_fd_sc_hd__or3_1
X_17717_ _05133_ VGND VGND VPWR VPWR _01182_ sky130_fd_sc_hd__clkbuf_1
X_30975_ clknet_leaf_166_clk _02710_ VGND VGND VPWR VPWR datamem.data_ram\[39\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_222_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18697_ _05749_ _06044_ _06048_ _05702_ _06050_ VGND VGND VPWR VPWR _06051_ sky130_fd_sc_hd__a221o_1
XFILLER_0_89_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_188_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23579__201 clknet_1_1__leaf__10176_ VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_63_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32714_ clknet_leaf_285_clk _04136_ VGND VGND VPWR VPWR datamem.data_ram\[17\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_17648_ net2617 _13222_ _05093_ VGND VGND VPWR VPWR _05097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_4283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_4294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_552 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32645_ clknet_leaf_153_clk _04067_ VGND VGND VPWR VPWR datamem.data_ram\[1\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_17579_ _05060_ VGND VGND VPWR VPWR _01247_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19318_ _06585_ rvcpu.dp.plem.ALUResultM\[4\] VGND VGND VPWR VPWR _06614_ sky130_fd_sc_hd__nand2_4
X_32576_ clknet_leaf_274_clk _03998_ VGND VGND VPWR VPWR datamem.data_ram\[22\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_20590_ _06666_ datamem.data_ram\[18\]\[13\] VGND VGND VPWR VPWR _07881_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31527_ clknet_leaf_29_clk net1193 VGND VGND VPWR VPWR rvcpu.dp.plem.PCPlus4M\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_19249_ _06552_ VGND VGND VPWR VPWR rvcpu.dp.lAuiPCE\[29\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22260_ _09387_ VGND VGND VPWR VPWR _09426_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_170_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31458_ clknet_leaf_75_clk rvcpu.dp.SrcBFW_Mux.y\[16\] VGND VGND VPWR VPWR rvcpu.dp.plem.WriteDataM\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_4508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21211_ _08489_ VGND VGND VPWR VPWR _08490_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_115_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30409_ net747 _02144_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[31\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_22191_ _09252_ net4387 _09362_ VGND VGND VPWR VPWR _09368_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31389_ clknet_leaf_41_clk _03092_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCE\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23551__175 clknet_1_0__leaf__10174_ VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_113_3198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21142_ datamem.data_ram\[63\]\[23\] _07859_ _06917_ datamem.data_ram\[61\]\[23\]
+ VGND VGND VPWR VPWR _08431_ sky130_fd_sc_hd__o22a_1
XFILLER_0_112_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25950_ net1651 _11155_ VGND VGND VPWR VPWR _11297_ sky130_fd_sc_hd__or2_1
X_21073_ _07635_ datamem.data_ram\[46\]\[7\] datamem.data_ram\[47\]\[7\] _07831_ rvcpu.dp.plem.ALUResultM\[3\]
+ VGND VGND VPWR VPWR _08362_ sky130_fd_sc_hd__o221a_1
XFILLER_0_158_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_3515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20024_ datamem.data_ram\[45\]\[2\] _06919_ _06941_ datamem.data_ram\[43\]\[2\] _07317_
+ VGND VGND VPWR VPWR _07318_ sky130_fd_sc_hd__a221o_1
X_24901_ _10667_ VGND VGND VPWR VPWR _02523_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_126_3526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25881_ rvcpu.dp.plfd.PCD\[0\] _11143_ VGND VGND VPWR VPWR _11257_ sky130_fd_sc_hd__or2_1
X_27620_ _12085_ net2653 net80 VGND VGND VPWR VPWR _12245_ sky130_fd_sc_hd__mux2_1
X_24832_ net104 _10600_ VGND VGND VPWR VPWR _10630_ sky130_fd_sc_hd__nor2_8
XFILLER_0_154_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_87_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27551_ _12208_ VGND VGND VPWR VPWR _03632_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_1247 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24763_ _10591_ VGND VGND VPWR VPWR _02461_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_87_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21975_ _08523_ _09203_ _09205_ _08575_ VGND VGND VPWR VPWR _09206_ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26502_ clknet_1_1__leaf__10079_ VGND VGND VPWR VPWR _11602_ sky130_fd_sc_hd__buf_1
XFILLER_0_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20926_ _07868_ _08214_ _08215_ _07863_ VGND VGND VPWR VPWR _08216_ sky130_fd_sc_hd__o22a_1
X_27482_ _12171_ VGND VGND VPWR VPWR _03600_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24694_ _10554_ VGND VGND VPWR VPWR _02429_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_0__10102_ _10102_ VGND VGND VPWR VPWR clknet_0__10102_ sky130_fd_sc_hd__clkbuf_16
X_29221_ _10072_ _13123_ VGND VGND VPWR VPWR _13130_ sky130_fd_sc_hd__and2_1
X_26433_ _11545_ rvcpu.ALUResultE\[17\] VGND VGND VPWR VPWR _11566_ sky130_fd_sc_hd__and2_1
XFILLER_0_95_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23645_ _09288_ net3312 _10182_ VGND VGND VPWR VPWR _10189_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20857_ _07823_ datamem.data_ram\[10\]\[14\] datamem.data_ram\[11\]\[14\] _07849_
+ _07867_ VGND VGND VPWR VPWR _08147_ sky130_fd_sc_hd__a221o_1
XFILLER_0_64_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29152_ _13092_ VGND VGND VPWR VPWR _04349_ sky130_fd_sc_hd__clkbuf_1
X_26364_ _11047_ _11511_ VGND VGND VPWR VPWR _11516_ sky130_fd_sc_hd__and2_1
XFILLER_0_153_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20788_ _08075_ _08076_ _08077_ _07822_ _07868_ VGND VGND VPWR VPWR _08078_ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28103_ _12516_ VGND VGND VPWR VPWR _03876_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25315_ _10902_ VGND VGND VPWR VPWR _02702_ sky130_fd_sc_hd__clkbuf_1
X_29083_ _12764_ net3422 _13049_ VGND VGND VPWR VPWR _13056_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22527_ _09636_ _09681_ VGND VGND VPWR VPWR _09682_ sky130_fd_sc_hd__or2_1
X_26295_ _11480_ VGND VGND VPWR VPWR _03104_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28034_ _12479_ VGND VGND VPWR VPWR _03844_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25246_ _10735_ net3630 net55 VGND VGND VPWR VPWR _10863_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22458_ rvcpu.dp.rf.reg_file_arr\[28\]\[8\] rvcpu.dp.rf.reg_file_arr\[30\]\[8\] rvcpu.dp.rf.reg_file_arr\[29\]\[8\]
+ rvcpu.dp.rf.reg_file_arr\[31\]\[8\] _09446_ _09402_ VGND VGND VPWR VPWR _09616_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_59_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23176__847 clknet_1_0__leaf__10111_ VGND VGND VPWR VPWR net973 sky130_fd_sc_hd__inv_2
X_21409_ rvcpu.dp.rf.reg_file_arr\[0\]\[2\] rvcpu.dp.rf.reg_file_arr\[1\]\[2\] rvcpu.dp.rf.reg_file_arr\[2\]\[2\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[2\] _08566_ _08569_ VGND VGND VPWR VPWR _08669_ sky130_fd_sc_hd__mux4_1
X_25177_ _10824_ net3090 _10812_ VGND VGND VPWR VPWR _10825_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22389_ rvcpu.dp.rf.reg_file_arr\[8\]\[4\] rvcpu.dp.rf.reg_file_arr\[10\]\[4\] rvcpu.dp.rf.reg_file_arr\[9\]\[4\]
+ rvcpu.dp.rf.reg_file_arr\[11\]\[4\] _09431_ _09532_ VGND VGND VPWR VPWR _09551_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_55_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29985_ net355 _01720_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[14\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28936_ _12762_ net2309 _12968_ VGND VGND VPWR VPWR _12974_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16950_ _04726_ VGND VGND VPWR VPWR _01566_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15901_ _14285_ VGND VGND VPWR VPWR _02074_ sky130_fd_sc_hd__clkbuf_1
X_16881_ net2885 _14432_ _04684_ VGND VGND VPWR VPWR _04690_ sky130_fd_sc_hd__mux2_1
XFILLER_0_218_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28867_ _12937_ VGND VGND VPWR VPWR _04219_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_202_5350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18620_ _05955_ _05959_ _05964_ _05977_ VGND VGND VPWR VPWR _05978_ sky130_fd_sc_hd__or4b_1
X_23528__155 clknet_1_1__leaf__10171_ VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__inv_2
X_15832_ net2028 _13213_ _14247_ VGND VGND VPWR VPWR _14248_ sky130_fd_sc_hd__mux2_1
X_27818_ _12153_ net2801 net78 VGND VGND VPWR VPWR _12352_ sky130_fd_sc_hd__mux2_1
X_28798_ _12743_ net3642 net70 VGND VGND VPWR VPWR _12901_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_194_5140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18551_ _05368_ _05585_ _05586_ _05654_ VGND VGND VPWR VPWR _05911_ sky130_fd_sc_hd__a31oi_1
X_15763_ _14151_ net3334 _14210_ VGND VGND VPWR VPWR _14211_ sky130_fd_sc_hd__mux2_1
X_27749_ _12138_ net2178 _12307_ VGND VGND VPWR VPWR _12314_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_194_5151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_194_5162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14714_ _13270_ VGND VGND VPWR VPWR _03175_ sky130_fd_sc_hd__clkbuf_1
X_17502_ _05019_ VGND VGND VPWR VPWR _01291_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_185_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30760_ clknet_leaf_149_clk _02495_ VGND VGND VPWR VPWR datamem.data_ram\[47\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_18482_ _05704_ _05669_ _05758_ VGND VGND VPWR VPWR _05844_ sky130_fd_sc_hd__or3_1
XFILLER_0_87_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15694_ _14166_ net3731 _14152_ VGND VGND VPWR VPWR _14167_ sky130_fd_sc_hd__mux2_1
XANTENNA_440 _07021_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_451 _07860_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_212_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_190_5048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17433_ _14147_ net3902 _04974_ VGND VGND VPWR VPWR _04983_ sky130_fd_sc_hd__mux2_1
XANTENNA_462 _08744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_190_5059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29419_ clknet_leaf_12_clk _01154_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD2E\[30\] sky130_fd_sc_hd__dfxtp_1
X_14645_ _13218_ VGND VGND VPWR VPWR _03192_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_170_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30691_ clknet_leaf_173_clk _02426_ VGND VGND VPWR VPWR datamem.data_ram\[4\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_473 _09281_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_170_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_484 _09386_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_184_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_495 _09892_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32430_ clknet_leaf_249_clk _03852_ VGND VGND VPWR VPWR datamem.data_ram\[28\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17364_ _04946_ VGND VGND VPWR VPWR _01356_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_16_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24014__546 clknet_1_1__leaf__10242_ VGND VGND VPWR VPWR net672 sky130_fd_sc_hd__inv_2
XFILLER_0_200_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19103_ _06423_ _06424_ VGND VGND VPWR VPWR _06425_ sky130_fd_sc_hd__xnor2_1
X_16315_ _14520_ VGND VGND VPWR VPWR _01879_ sky130_fd_sc_hd__clkbuf_1
X_32361_ clknet_leaf_94_clk _03783_ VGND VGND VPWR VPWR datamem.data_ram\[2\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17295_ net4329 _13203_ _04902_ VGND VGND VPWR VPWR _04910_ sky130_fd_sc_hd__mux2_1
X_19034_ _06362_ _06364_ VGND VGND VPWR VPWR _06365_ sky130_fd_sc_hd__xor2_2
X_31312_ clknet_leaf_45_clk _03015_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCPlus4E\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_16246_ net2799 _14482_ _14464_ VGND VGND VPWR VPWR _14483_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32292_ clknet_leaf_225_clk _03714_ VGND VGND VPWR VPWR datamem.data_ram\[32\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_209_5504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_209_5515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31243_ clknet_leaf_21_clk _02946_ VGND VGND VPWR VPWR rvcpu.dp.plfd.InstrD\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_16177_ _13203_ VGND VGND VPWR VPWR _14436_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15128_ _13671_ _13562_ _13672_ VGND VGND VPWR VPWR _13673_ sky130_fd_sc_hd__or3_1
XFILLER_0_23_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31174_ clknet_leaf_214_clk _02877_ VGND VGND VPWR VPWR datamem.data_ram\[5\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_227_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_290_clk clknet_5_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_290_clk
+ sky130_fd_sc_hd__clkbuf_8
X_30125_ net487 _01860_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[10\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_15059_ _13603_ _13605_ _13501_ VGND VGND VPWR VPWR _13606_ sky130_fd_sc_hd__a21oi_1
X_19936_ _06805_ VGND VGND VPWR VPWR _07230_ sky130_fd_sc_hd__buf_6
XFILLER_0_220_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2907 rvcpu.dp.rf.reg_file_arr\[14\]\[10\] VGND VGND VPWR VPWR net4057 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2918 datamem.data_ram\[62\]\[19\] VGND VGND VPWR VPWR net4068 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2929 datamem.data_ram\[61\]\[19\] VGND VGND VPWR VPWR net4079 sky130_fd_sc_hd__dlygate4sd3_1
X_30056_ net418 _01791_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[12\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_19867_ datamem.data_ram\[10\]\[1\] _06932_ _06973_ datamem.data_ram\[8\]\[1\] _07031_
+ VGND VGND VPWR VPWR _07162_ sky130_fd_sc_hd__a221o_1
XFILLER_0_128_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18818_ _05239_ _06152_ _06154_ _06164_ VGND VGND VPWR VPWR rvcpu.ALUResultE\[17\]
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_218_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19798_ datamem.data_ram\[57\]\[9\] _06783_ _07091_ _07092_ VGND VGND VPWR VPWR _07093_
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_121_3401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18749_ _05658_ _06097_ _06099_ _06075_ VGND VGND VPWR VPWR _06100_ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_210_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_222_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1052 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21760_ _08672_ _08994_ _08998_ _09002_ VGND VGND VPWR VPWR _09003_ sky130_fd_sc_hd__and4_1
X_30958_ clknet_leaf_156_clk _02693_ VGND VGND VPWR VPWR datamem.data_ram\[3\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_1074 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20711_ datamem.data_ram\[27\]\[5\] _06966_ _08000_ _08001_ VGND VGND VPWR VPWR _08002_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_4_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21691_ _08935_ _08936_ _08743_ VGND VGND VPWR VPWR _08937_ sky130_fd_sc_hd__mux2_1
XFILLER_0_176_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30889_ clknet_leaf_219_clk _02624_ VGND VGND VPWR VPWR datamem.data_ram\[42\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32628_ clknet_leaf_93_clk _04050_ VGND VGND VPWR VPWR datamem.data_ram\[1\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20642_ datamem.data_ram\[18\]\[29\] _06803_ _06823_ datamem.data_ram\[21\]\[29\]
+ _06733_ VGND VGND VPWR VPWR _07933_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_119_3341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_119_3352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_335 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20573_ datamem.data_ram\[36\]\[13\] datamem.data_ram\[37\]\[13\] _07828_ VGND VGND
+ VPWR VPWR _07864_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32559_ clknet_leaf_184_clk _03981_ VGND VGND VPWR VPWR datamem.data_ram\[22\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25100_ _10067_ VGND VGND VPWR VPWR _10782_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_115_3249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22312_ _09462_ VGND VGND VPWR VPWR _09477_ sky130_fd_sc_hd__buf_4
X_26080_ _11371_ VGND VGND VPWR VPWR _11372_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_41_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23292_ clknet_1_0__leaf__10130_ VGND VGND VPWR VPWR _10132_ sky130_fd_sc_hd__buf_1
XFILLER_0_15_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25031_ _07137_ VGND VGND VPWR VPWR _10741_ sky130_fd_sc_hd__buf_8
X_22243_ rvcpu.dp.rf.reg_file_arr\[20\]\[0\] rvcpu.dp.rf.reg_file_arr\[21\]\[0\] rvcpu.dp.rf.reg_file_arr\[22\]\[0\]
+ rvcpu.dp.rf.reg_file_arr\[23\]\[0\] _09406_ _09408_ VGND VGND VPWR VPWR _09409_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_48_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22174_ _09358_ VGND VGND VPWR VPWR _01105_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_169_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_281_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_281_clk
+ sky130_fd_sc_hd__clkbuf_8
X_21125_ _06666_ datamem.data_ram\[43\]\[23\] _06944_ datamem.data_ram\[42\]\[23\]
+ _07838_ VGND VGND VPWR VPWR _08414_ sky130_fd_sc_hd__a221o_1
X_26982_ _10113_ _10337_ _11713_ VGND VGND VPWR VPWR _11875_ sky130_fd_sc_hd__a21oi_4
X_29770_ net1116 _01505_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[20\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_50_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25933_ rvcpu.dp.plfd.PCD\[22\] _11279_ VGND VGND VPWR VPWR _11287_ sky130_fd_sc_hd__or2_1
X_28721_ _12751_ net2360 _12859_ VGND VGND VPWR VPWR _12860_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_89_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21056_ _07859_ _08339_ _08344_ _06732_ VGND VGND VPWR VPWR _08345_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_89_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20007_ datamem.data_ram\[61\]\[2\] _06920_ _06942_ datamem.data_ram\[59\]\[2\] _07300_
+ VGND VGND VPWR VPWR _07301_ sky130_fd_sc_hd__a221o_1
XFILLER_0_214_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_185_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_145_3979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28652_ _12279_ _12602_ _12795_ VGND VGND VPWR VPWR _12823_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_199_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25864_ _11243_ VGND VGND VPWR VPWR _02910_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_213_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23976__512 clknet_1_1__leaf__10238_ VGND VGND VPWR VPWR net638 sky130_fd_sc_hd__inv_2
X_24815_ _10297_ _10347_ _10611_ VGND VGND VPWR VPWR _10621_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_2_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27603_ _12147_ net3326 net81 VGND VGND VPWR VPWR _12236_ sky130_fd_sc_hd__mux2_1
X_28583_ _10141_ _12622_ _12668_ VGND VGND VPWR VPWR _12786_ sky130_fd_sc_hd__a21oi_4
X_25795_ rvcpu.dp.pcreg.q\[15\] rvcpu.dp.pcreg.q\[14\] _11182_ VGND VGND VPWR VPWR
+ _11188_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_2_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27534_ _12199_ VGND VGND VPWR VPWR _03624_ sky130_fd_sc_hd__clkbuf_1
X_24746_ _10582_ VGND VGND VPWR VPWR _02453_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_179_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21958_ rvcpu.dp.rf.reg_file_arr\[8\]\[30\] rvcpu.dp.rf.reg_file_arr\[10\]\[30\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[30\] rvcpu.dp.rf.reg_file_arr\[11\]\[30\] _08534_
+ _08537_ VGND VGND VPWR VPWR _09190_ sky130_fd_sc_hd__mux4_1
XFILLER_0_69_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20909_ datamem.data_ram\[16\]\[22\] _07829_ VGND VGND VPWR VPWR _08199_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26485__39 clknet_1_1__leaf__10267_ VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__inv_2
X_27465_ _12085_ net3004 net83 VGND VGND VPWR VPWR _12162_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_104_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24677_ _10545_ VGND VGND VPWR VPWR _02421_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21889_ _08547_ _09122_ _09124_ _08575_ VGND VGND VPWR VPWR _09125_ sky130_fd_sc_hd__o211a_1
X_26416_ _06425_ _11539_ _11529_ _11176_ _11554_ VGND VGND VPWR VPWR _11555_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_13_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29204_ _09329_ net2152 _13112_ VGND VGND VPWR VPWR _13120_ sky130_fd_sc_hd__mux2_1
XFILLER_0_204_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27396_ _12083_ net2420 net85 VGND VGND VPWR VPWR _12118_ sky130_fd_sc_hd__mux2_1
X_29135_ _13083_ VGND VGND VPWR VPWR _04341_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_706 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26347_ _10061_ _11507_ _11508_ net1344 VGND VGND VPWR VPWR _03128_ sky130_fd_sc_hd__a22o_1
XFILLER_0_181_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_182_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16100_ net2569 _13201_ _14385_ VGND VGND VPWR VPWR _14392_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17080_ _14135_ net2915 _04793_ VGND VGND VPWR VPWR _04796_ sky130_fd_sc_hd__mux2_1
X_29066_ _09287_ net2539 _13040_ VGND VGND VPWR VPWR _13047_ sky130_fd_sc_hd__mux2_1
X_26278_ _11471_ VGND VGND VPWR VPWR _03096_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28017_ _12470_ VGND VGND VPWR VPWR _03836_ sky130_fd_sc_hd__clkbuf_1
X_16031_ _14355_ VGND VGND VPWR VPWR _02006_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_161_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25229_ _10762_ net3059 _10848_ VGND VGND VPWR VPWR _10854_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_1292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26516__4 clknet_1_1__leaf__10080_ VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_204_5401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_272_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_272_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_202_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_176_Right_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17982_ _05176_ _05350_ _05351_ _05352_ VGND VGND VPWR VPWR rvcpu.dp.SrcBFW_Mux.y\[6\]
+ sky130_fd_sc_hd__a31o_1
X_29968_ net338 _01703_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[15\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19721_ _06799_ _06915_ _07016_ VGND VGND VPWR VPWR _07017_ sky130_fd_sc_hd__o21ba_1
X_16933_ net3265 _14484_ _04683_ VGND VGND VPWR VPWR _04717_ sky130_fd_sc_hd__mux2_1
X_28919_ _12698_ net4196 _12959_ VGND VGND VPWR VPWR _12965_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_196_5202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29899_ net277 _01634_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[17\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19652_ _06947_ VGND VGND VPWR VPWR _06948_ sky130_fd_sc_hd__buf_4
X_31930_ clknet_leaf_112_clk _03352_ VGND VGND VPWR VPWR datamem.data_ram\[60\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_16864_ _04680_ VGND VGND VPWR VPWR _01606_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_221_5792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18603_ _05799_ _05840_ VGND VGND VPWR VPWR _05961_ sky130_fd_sc_hd__nand2_1
X_15815_ net2039 _13187_ _14236_ VGND VGND VPWR VPWR _14239_ sky130_fd_sc_hd__mux2_1
X_31861_ clknet_leaf_124_clk _03315_ VGND VGND VPWR VPWR datamem.data_ram\[62\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_16795_ net4393 _14482_ _04634_ VGND VGND VPWR VPWR _04644_ sky130_fd_sc_hd__mux2_1
X_19583_ datamem.data_ram\[37\]\[8\] _06815_ _06877_ _06878_ VGND VGND VPWR VPWR _06879_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_189_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30812_ clknet_leaf_135_clk _02547_ VGND VGND VPWR VPWR datamem.data_ram\[45\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_18534_ _05349_ _05358_ _05684_ VGND VGND VPWR VPWR _05895_ sky130_fd_sc_hd__mux2_1
X_15746_ _14135_ net3322 _14199_ VGND VGND VPWR VPWR _14202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31792_ clknet_leaf_213_clk _03246_ VGND VGND VPWR VPWR datamem.data_ram\[2\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23345__983 clknet_1_1__leaf__10136_ VGND VGND VPWR VPWR net1109 sky130_fd_sc_hd__inv_2
XFILLER_0_88_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_213_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_201_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_4220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_213_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18465_ _05741_ _05826_ _05827_ _05667_ VGND VGND VPWR VPWR _05828_ sky130_fd_sc_hd__o22a_1
X_30743_ clknet_leaf_150_clk _02478_ VGND VGND VPWR VPWR datamem.data_ram\[48\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_23502__147 clknet_1_0__leaf__10161_ VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__inv_2
XFILLER_0_47_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15677_ _14155_ VGND VGND VPWR VPWR _02176_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_200_450 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_270 _13232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_201_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_281 _13260_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_201_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_292 _13350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17416_ _04973_ VGND VGND VPWR VPWR _04974_ sky130_fd_sc_hd__clkbuf_4
X_14628_ _13205_ VGND VGND VPWR VPWR _03196_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_185_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18396_ _05527_ _05533_ _05683_ VGND VGND VPWR VPWR _05760_ sky130_fd_sc_hd__mux2_1
X_30674_ clknet_leaf_190_clk _02409_ VGND VGND VPWR VPWR datamem.data_ram\[50\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_151_4117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_151_4128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32413_ clknet_leaf_246_clk _03835_ VGND VGND VPWR VPWR datamem.data_ram\[28\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17347_ _14128_ _04900_ VGND VGND VPWR VPWR _04937_ sky130_fd_sc_hd__nand2_2
XFILLER_0_172_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32344_ clknet_leaf_182_clk _03766_ VGND VGND VPWR VPWR datamem.data_ram\[30\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload201 clknet_leaf_209_clk VGND VGND VPWR VPWR clkload201/Y sky130_fd_sc_hd__clkinvlp_2
X_17278_ _13174_ rvcpu.dp.plmw.RdW\[3\] _13176_ VGND VGND VPWR VPWR _04900_ sky130_fd_sc_hd__and3b_1
Xclkload212 clknet_leaf_206_clk VGND VGND VPWR VPWR clkload212/Y sky130_fd_sc_hd__clkinvlp_2
Xclkload223 clknet_leaf_162_clk VGND VGND VPWR VPWR clkload223/Y sky130_fd_sc_hd__clkinv_1
XFILLER_0_130_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload234 clknet_leaf_113_clk VGND VGND VPWR VPWR clkload234/Y sky130_fd_sc_hd__clkinv_1
X_19017_ _06339_ _06340_ _06344_ _06350_ VGND VGND VPWR VPWR _06351_ sky130_fd_sc_hd__a211o_1
X_16229_ _14471_ VGND VGND VPWR VPWR _01924_ sky130_fd_sc_hd__clkbuf_1
Xclkload245 clknet_leaf_157_clk VGND VGND VPWR VPWR clkload245/Y sky130_fd_sc_hd__clkinvlp_2
X_32275_ clknet_leaf_167_clk _03697_ VGND VGND VPWR VPWR datamem.data_ram\[33\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload256 clknet_leaf_142_clk VGND VGND VPWR VPWR clkload256/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_12_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_228_5957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload267 clknet_leaf_126_clk VGND VGND VPWR VPWR clkload267/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_110_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_228_5968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31226_ clknet_leaf_50_clk _02929_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCD\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload278 clknet_1_1__leaf__10078_ VGND VGND VPWR VPWR clkload278/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_110_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_228_5979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload289 clknet_1_1__leaf__10239_ VGND VGND VPWR VPWR clkload289/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_110_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_4068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23845__409 clknet_1_1__leaf__10208_ VGND VGND VPWR VPWR net535 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_149_4079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_263_clk clknet_5_17__leaf_clk VGND VGND VPWR VPWR clknet_leaf_263_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_228_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31157_ clknet_leaf_46_clk rvcpu.ALUResultE\[16\] VGND VGND VPWR VPWR rvcpu.dp.plem.ALUResultM\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_181_4836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_181_4847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_143_Right_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2704 datamem.data_ram\[34\]\[14\] VGND VGND VPWR VPWR net3854 sky130_fd_sc_hd__dlygate4sd3_1
X_30108_ net470 _01843_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[11\]\[31\] sky130_fd_sc_hd__dfxtp_1
Xhold2715 datamem.data_ram\[56\]\[26\] VGND VGND VPWR VPWR net3865 sky130_fd_sc_hd__dlygate4sd3_1
X_19919_ datamem.data_ram\[63\]\[17\] _07020_ _06620_ datamem.data_ram\[60\]\[17\]
+ VGND VGND VPWR VPWR _07214_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_71_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2726 datamem.data_ram\[9\]\[26\] VGND VGND VPWR VPWR net3876 sky130_fd_sc_hd__dlygate4sd3_1
X_31088_ clknet_leaf_100_clk _02823_ VGND VGND VPWR VPWR datamem.data_ram\[21\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2737 datamem.data_ram\[21\]\[29\] VGND VGND VPWR VPWR net3887 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2748 rvcpu.dp.rf.reg_file_arr\[17\]\[11\] VGND VGND VPWR VPWR net3898 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2759 datamem.data_ram\[60\]\[30\] VGND VGND VPWR VPWR net3909 sky130_fd_sc_hd__dlygate4sd3_1
X_22930_ _10061_ _10053_ VGND VGND VPWR VPWR _10062_ sky130_fd_sc_hd__and2_1
X_30039_ net401 _01774_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[13\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_84_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22861_ _09433_ _09997_ _09789_ VGND VGND VPWR VPWR _09998_ sky130_fd_sc_hd__a21o_1
XFILLER_0_196_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_140_3854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24600_ _10209_ _10327_ _10501_ VGND VGND VPWR VPWR _10502_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_179_4787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21812_ rvcpu.dp.rf.reg_file_arr\[8\]\[22\] rvcpu.dp.rf.reg_file_arr\[10\]\[22\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[22\] rvcpu.dp.rf.reg_file_arr\[11\]\[22\] _08534_
+ _08818_ VGND VGND VPWR VPWR _09052_ sky130_fd_sc_hd__mux4_1
XFILLER_0_223_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25580_ _10076_ _11042_ VGND VGND VPWR VPWR _11051_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_179_4798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire42 _12841_ VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__buf_4
X_22792_ rvcpu.dp.rf.reg_file_arr\[0\]\[25\] rvcpu.dp.rf.reg_file_arr\[1\]\[25\] rvcpu.dp.rf.reg_file_arr\[2\]\[25\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[25\] _09477_ _09466_ VGND VGND VPWR VPWR _09933_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_78_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire53 _11066_ VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__buf_4
XFILLER_0_190_1288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24531_ _10394_ datamem.data_ram\[52\]\[12\] _10456_ VGND VGND VPWR VPWR _10461_
+ sky130_fd_sc_hd__mux2_1
X_21743_ rvcpu.dp.rf.reg_file_arr\[16\]\[19\] rvcpu.dp.rf.reg_file_arr\[17\]\[19\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[19\] rvcpu.dp.rf.reg_file_arr\[19\]\[19\] _08799_
+ _08800_ VGND VGND VPWR VPWR _08986_ sky130_fd_sc_hd__mux4_2
X_27250_ _11978_ _12031_ VGND VGND VPWR VPWR _12039_ sky130_fd_sc_hd__and2_1
XFILLER_0_148_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24462_ _10412_ net3744 _10404_ _10420_ VGND VGND VPWR VPWR _02331_ sky130_fd_sc_hd__a31o_1
XFILLER_0_175_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21674_ rvcpu.dp.rf.reg_file_arr\[28\]\[15\] rvcpu.dp.rf.reg_file_arr\[30\]\[15\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[15\] rvcpu.dp.rf.reg_file_arr\[31\]\[15\] _08559_
+ _08636_ VGND VGND VPWR VPWR _08921_ sky130_fd_sc_hd__mux4_1
XFILLER_0_176_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26201_ _11375_ _11438_ _11372_ VGND VGND VPWR VPWR _03052_ sky130_fd_sc_hd__o21a_1
XFILLER_0_149_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27181_ _11991_ net1516 _11995_ _11998_ VGND VGND VPWR VPWR _03472_ sky130_fd_sc_hd__a31o_1
XFILLER_0_11_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20625_ datamem.data_ram\[10\]\[13\] _06610_ _06781_ datamem.data_ram\[9\]\[13\]
+ _07915_ VGND VGND VPWR VPWR _07916_ sky130_fd_sc_hd__o221a_1
X_24393_ _10375_ VGND VGND VPWR VPWR _02307_ sky130_fd_sc_hd__clkbuf_1
X_26132_ net1858 _11397_ VGND VGND VPWR VPWR _11402_ sky130_fd_sc_hd__and2_1
X_23557__181 clknet_1_0__leaf__10174_ VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__inv_2
XFILLER_0_62_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20556_ datamem.data_ram\[14\]\[21\] _07028_ _06649_ datamem.data_ram\[8\]\[21\]
+ VGND VGND VPWR VPWR _07847_ sky130_fd_sc_hd__o22a_1
X_26063_ _11353_ net3462 _11350_ _11360_ VGND VGND VPWR VPWR _02992_ sky130_fd_sc_hd__a31o_1
XFILLER_0_81_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20487_ _06751_ _07773_ _07778_ _06594_ VGND VGND VPWR VPWR _07779_ sky130_fd_sc_hd__o31a_1
XFILLER_0_120_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25014_ _10729_ net3799 net100 VGND VGND VPWR VPWR _10730_ sky130_fd_sc_hd__mux2_1
X_22226_ _08592_ VGND VGND VPWR VPWR _09392_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_219_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_5_Left_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_254_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_254_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_203_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29822_ net200 _01557_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[1\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22157_ _09348_ VGND VGND VPWR VPWR _01098_ sky130_fd_sc_hd__clkbuf_1
X_24043__572 clknet_1_1__leaf__10245_ VGND VGND VPWR VPWR net698 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_110_Right_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21108_ _06640_ _08396_ VGND VGND VPWR VPWR _08397_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_7_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29753_ net1099 _01488_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[21\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_7_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26965_ _10402_ _10947_ VGND VGND VPWR VPWR _11866_ sky130_fd_sc_hd__nor2_1
X_22088_ _09299_ _09301_ _09231_ VGND VGND VPWR VPWR _09302_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_22_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28704_ _12687_ net3774 _12850_ VGND VGND VPWR VPWR _12851_ sky130_fd_sc_hd__mux2_1
X_25916_ net2062 _11275_ _11273_ _11277_ VGND VGND VPWR VPWR _02928_ sky130_fd_sc_hd__o211a_1
X_21039_ net122 datamem.data_ram\[14\]\[31\] datamem.data_ram\[15\]\[31\] _06639_
+ _06641_ VGND VGND VPWR VPWR _08328_ sky130_fd_sc_hd__o221a_1
X_26896_ _11820_ VGND VGND VPWR VPWR _11821_ sky130_fd_sc_hd__buf_2
X_29684_ net1030 _01419_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[23\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_214_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_195_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_195_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25847_ _11206_ _11207_ _11229_ VGND VGND VPWR VPWR _11230_ sky130_fd_sc_hd__and3_1
X_28635_ _10777_ _12622_ _12795_ VGND VGND VPWR VPWR _12814_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_92_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15600_ net3187 _13226_ _14103_ VGND VGND VPWR VPWR _14108_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_18_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16580_ _14181_ net4313 _04525_ VGND VGND VPWR VPWR _04530_ sky130_fd_sc_hd__mux2_1
X_25778_ rvcpu.dp.pcreg.q\[11\] _11171_ VGND VGND VPWR VPWR _11175_ sky130_fd_sc_hd__or2_1
XFILLER_0_186_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28566_ _10141_ _12612_ _12668_ VGND VGND VPWR VPWR _12777_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_9_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15531_ _13517_ _13302_ _13941_ _14056_ VGND VGND VPWR VPWR _14057_ sky130_fd_sc_hd__a211o_1
X_24729_ _10573_ VGND VGND VPWR VPWR _02445_ sky130_fd_sc_hd__clkbuf_1
X_27517_ _12190_ VGND VGND VPWR VPWR _03616_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28497_ _11980_ _12724_ VGND VGND VPWR VPWR _12733_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18250_ _05603_ _05314_ _05600_ _05609_ _05614_ VGND VGND VPWR VPWR _05615_ sky130_fd_sc_hd__o221a_1
XFILLER_0_127_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_831 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15462_ _13496_ _13990_ _13991_ VGND VGND VPWR VPWR _13992_ sky130_fd_sc_hd__a21oi_1
X_27448_ _09281_ VGND VGND VPWR VPWR _12151_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_56_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23950__504 clknet_1_0__leaf__10228_ VGND VGND VPWR VPWR net630 sky130_fd_sc_hd__inv_2
XFILLER_0_167_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17201_ _04859_ VGND VGND VPWR VPWR _01440_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18181_ rvcpu.dp.plde.ImmExtE\[26\] rvcpu.dp.SrcBFW_Mux.y\[26\] _05279_ VGND VGND
+ VPWR VPWR _05546_ sky130_fd_sc_hd__mux2_1
X_15393_ _13419_ _13603_ _13381_ _13599_ VGND VGND VPWR VPWR _13926_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_5_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27379_ _10727_ net3014 net86 VGND VGND VPWR VPWR _12109_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17132_ _14187_ net4348 _04815_ VGND VGND VPWR VPWR _04823_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29118_ _13074_ VGND VGND VPWR VPWR _04333_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_163_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30390_ net728 _02125_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[31\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29049_ _10072_ _13031_ VGND VGND VPWR VPWR _13038_ sky130_fd_sc_hd__and2_1
XFILLER_0_162_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17063_ _04786_ VGND VGND VPWR VPWR _01505_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16014_ net2429 _13278_ _14310_ VGND VGND VPWR VPWR _14345_ sky130_fd_sc_hd__mux2_1
X_32060_ clknet_leaf_119_clk _03482_ VGND VGND VPWR VPWR datamem.data_ram\[48\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31011_ clknet_leaf_158_clk _02746_ VGND VGND VPWR VPWR datamem.data_ram\[11\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_245_clk clknet_5_17__leaf_clk VGND VGND VPWR VPWR clknet_leaf_245_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_110_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_223_5843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_223_5854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17965_ _05335_ _05316_ _05315_ VGND VGND VPWR VPWR _05336_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_104_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_178_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19704_ _06932_ VGND VGND VPWR VPWR _07000_ sky130_fd_sc_hd__clkbuf_8
X_16916_ _04708_ VGND VGND VPWR VPWR _01582_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32962_ clknet_leaf_208_clk _04384_ VGND VGND VPWR VPWR datamem.data_ram\[63\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17896_ _05268_ _05263_ VGND VGND VPWR VPWR _05269_ sky130_fd_sc_hd__nor2_4
XFILLER_0_109_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19635_ _06930_ VGND VGND VPWR VPWR _06931_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_192_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31913_ _04424_ net121 VGND VGND VPWR VPWR datamem.rd_data_mem\[18\] sky130_fd_sc_hd__dlxtn_1
X_16847_ net2823 _14466_ _04670_ VGND VGND VPWR VPWR _04672_ sky130_fd_sc_hd__mux2_1
X_32893_ clknet_leaf_163_clk _04315_ VGND VGND VPWR VPWR datamem.data_ram\[10\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_178_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31844_ clknet_leaf_91_clk _03298_ VGND VGND VPWR VPWR datamem.data_ram\[8\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_69_Left_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19566_ _06836_ _06861_ VGND VGND VPWR VPWR _06862_ sky130_fd_sc_hd__nor2_4
X_16778_ _04635_ VGND VGND VPWR VPWR _01655_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_220_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_177_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18517_ _05704_ _05690_ VGND VGND VPWR VPWR _05878_ sky130_fd_sc_hd__and2_1
X_15729_ _14190_ VGND VGND VPWR VPWR _02159_ sky130_fd_sc_hd__clkbuf_1
X_19497_ datamem.data_ram\[29\]\[16\] _06664_ _06791_ _06792_ VGND VGND VPWR VPWR
+ _06793_ sky130_fd_sc_hd__o211a_1
X_31775_ clknet_leaf_250_clk _03229_ VGND VGND VPWR VPWR datamem.data_ram\[6\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_220_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_174_4662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_4673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18448_ _05810_ _05684_ _05771_ VGND VGND VPWR VPWR _05811_ sky130_fd_sc_hd__or3_1
XFILLER_0_34_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30726_ clknet_leaf_216_clk _02461_ VGND VGND VPWR VPWR datamem.data_ram\[48\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18379_ _05284_ _05290_ _05647_ _05656_ _05742_ VGND VGND VPWR VPWR _05743_ sky130_fd_sc_hd__a311o_1
XFILLER_0_12_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30657_ clknet_leaf_219_clk _02392_ VGND VGND VPWR VPWR datamem.data_ram\[50\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_209_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20410_ _06776_ _07694_ _07696_ _07701_ VGND VGND VPWR VPWR _07702_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_212_Right_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_209_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21390_ _08572_ _08650_ VGND VGND VPWR VPWR _08651_ sky130_fd_sc_hd__or2_1
X_30588_ clknet_leaf_192_clk _02323_ VGND VGND VPWR VPWR datamem.data_ram\[53\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_77_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20341_ datamem.data_ram\[61\]\[4\] _06970_ _06977_ datamem.data_ram\[60\]\[4\] _07632_
+ VGND VGND VPWR VPWR _07633_ sky130_fd_sc_hd__a221o_1
X_32327_ clknet_leaf_87_clk _03749_ VGND VGND VPWR VPWR datamem.data_ram\[31\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_133_3680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_133_3691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23428__80 clknet_1_1__leaf__10154_ VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__inv_2
X_20272_ datamem.data_ram\[34\]\[19\] _06728_ _06737_ datamem.data_ram\[35\]\[19\]
+ _06733_ VGND VGND VPWR VPWR _07565_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_73_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32258_ clknet_leaf_259_clk _03680_ VGND VGND VPWR VPWR datamem.data_ram\[34\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_73_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22011_ rvcpu.dp.plem.WriteDataM\[2\] _09215_ _09219_ _09238_ VGND VGND VPWR VPWR
+ _09239_ sky130_fd_sc_hd__a31o_4
Xclkbuf_leaf_236_clk clknet_5_20__leaf_clk VGND VGND VPWR VPWR clknet_leaf_236_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_101_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31209_ clknet_leaf_22_clk _02912_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCPlus4D\[30\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3202 datamem.data_ram\[2\]\[22\] VGND VGND VPWR VPWR net4352 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3213 rvcpu.dp.plde.ImmExtE\[18\] VGND VGND VPWR VPWR net4363 sky130_fd_sc_hd__dlygate4sd3_1
X_32189_ clknet_leaf_241_clk _03611_ VGND VGND VPWR VPWR datamem.data_ram\[37\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3224 datamem.data_ram\[58\]\[18\] VGND VGND VPWR VPWR net4374 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_228_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23443__94 clknet_1_0__leaf__10155_ VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__inv_2
Xhold3235 datamem.data_ram\[14\]\[14\] VGND VGND VPWR VPWR net4385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2501 datamem.data_ram\[1\]\[23\] VGND VGND VPWR VPWR net3651 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3246 datamem.data_ram\[52\]\[13\] VGND VGND VPWR VPWR net4396 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3257 datamem.data_ram\[16\]\[15\] VGND VGND VPWR VPWR net4407 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2512 datamem.data_ram\[50\]\[10\] VGND VGND VPWR VPWR net3662 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3268 datamem.data_ram\[53\]\[14\] VGND VGND VPWR VPWR net4418 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2523 datamem.data_ram\[9\]\[12\] VGND VGND VPWR VPWR net3673 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2534 datamem.data_ram\[8\]\[22\] VGND VGND VPWR VPWR net3684 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3279 rvcpu.dp.rf.reg_file_arr\[24\]\[19\] VGND VGND VPWR VPWR net4429 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1800 rvcpu.dp.rf.reg_file_arr\[11\]\[30\] VGND VGND VPWR VPWR net2950 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2545 datamem.data_ram\[10\]\[29\] VGND VGND VPWR VPWR net3695 sky130_fd_sc_hd__dlygate4sd3_1
X_26750_ _11689_ _11726_ VGND VGND VPWR VPWR _11733_ sky130_fd_sc_hd__and2_1
Xhold2556 datamem.data_ram\[24\]\[12\] VGND VGND VPWR VPWR net3706 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1811 rvcpu.dp.rf.reg_file_arr\[30\]\[6\] VGND VGND VPWR VPWR net2961 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1822 datamem.data_ram\[17\]\[21\] VGND VGND VPWR VPWR net2972 sky130_fd_sc_hd__dlygate4sd3_1
X_23962_ _09252_ net4350 _10229_ VGND VGND VPWR VPWR _10235_ sky130_fd_sc_hd__mux2_1
XFILLER_0_192_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2567 datamem.data_ram\[3\]\[20\] VGND VGND VPWR VPWR net3717 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2578 rvcpu.dp.rf.reg_file_arr\[11\]\[14\] VGND VGND VPWR VPWR net3728 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1833 datamem.data_ram\[61\]\[13\] VGND VGND VPWR VPWR net2983 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2589 datamem.data_ram\[43\]\[19\] VGND VGND VPWR VPWR net3739 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1844 rvcpu.dp.rf.reg_file_arr\[12\]\[7\] VGND VGND VPWR VPWR net2994 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25701_ _08144_ net109 VGND VGND VPWR VPWR _11123_ sky130_fd_sc_hd__nor2_8
X_22913_ rvcpu.dp.plem.WriteDataM\[0\] VGND VGND VPWR VPWR _10047_ sky130_fd_sc_hd__clkbuf_4
Xhold1855 rvcpu.dp.rf.reg_file_arr\[24\]\[21\] VGND VGND VPWR VPWR net3005 sky130_fd_sc_hd__dlygate4sd3_1
X_26681_ _10297_ _11054_ _11609_ VGND VGND VPWR VPWR _11694_ sky130_fd_sc_hd__and3_1
Xhold1866 datamem.data_ram\[18\]\[15\] VGND VGND VPWR VPWR net3016 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1877 rvcpu.dp.rf.reg_file_arr\[2\]\[30\] VGND VGND VPWR VPWR net3027 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1888 rvcpu.dp.rf.reg_file_arr\[13\]\[15\] VGND VGND VPWR VPWR net3038 sky130_fd_sc_hd__dlygate4sd3_1
X_25632_ _11083_ _11079_ VGND VGND VPWR VPWR _11084_ sky130_fd_sc_hd__and2_1
X_28420_ _09297_ VGND VGND VPWR VPWR _12687_ sky130_fd_sc_hd__clkbuf_2
Xhold1899 datamem.data_ram\[46\]\[13\] VGND VGND VPWR VPWR net3049 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22844_ _09415_ _09979_ _09981_ _09473_ VGND VGND VPWR VPWR _09982_ sky130_fd_sc_hd__o211a_1
XFILLER_0_195_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__10181_ clknet_0__10181_ VGND VGND VPWR VPWR clknet_1_1__leaf__10181_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28351_ _09225_ _12622_ _12573_ VGND VGND VPWR VPWR _12650_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25563_ _11040_ VGND VGND VPWR VPWR _11041_ sky130_fd_sc_hd__buf_2
XFILLER_0_6_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22775_ _09452_ _09914_ _09916_ _09795_ VGND VGND VPWR VPWR _09917_ sky130_fd_sc_hd__a211o_1
XFILLER_0_94_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27302_ _12064_ VGND VGND VPWR VPWR _12065_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_94_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24514_ _10450_ datamem.data_ram\[52\]\[21\] _10440_ VGND VGND VPWR VPWR _10451_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28282_ _12601_ _12612_ _12573_ VGND VGND VPWR VPWR _12613_ sky130_fd_sc_hd__a21oi_4
X_21726_ rvcpu.dp.rf.reg_file_arr\[20\]\[18\] rvcpu.dp.rf.reg_file_arr\[21\]\[18\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[18\] rvcpu.dp.rf.reg_file_arr\[23\]\[18\] _08778_
+ _08825_ VGND VGND VPWR VPWR _08970_ sky130_fd_sc_hd__mux4_1
XFILLER_0_66_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25494_ _10816_ net3876 _10999_ VGND VGND VPWR VPWR _11002_ sky130_fd_sc_hd__mux2_1
X_27233_ _12022_ net1399 _12018_ _12028_ VGND VGND VPWR VPWR _03494_ sky130_fd_sc_hd__a31o_1
XFILLER_0_136_335 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24445_ _10056_ net1829 _10404_ _10409_ VGND VGND VPWR VPWR _02325_ sky130_fd_sc_hd__a31o_1
XFILLER_0_93_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21657_ rvcpu.dp.rf.reg_file_arr\[20\]\[14\] rvcpu.dp.rf.reg_file_arr\[21\]\[14\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[14\] rvcpu.dp.rf.reg_file_arr\[23\]\[14\] _08524_
+ _08527_ VGND VGND VPWR VPWR _08905_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_62_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23713__306 clknet_1_0__leaf__10197_ VGND VGND VPWR VPWR net432 sky130_fd_sc_hd__inv_2
XFILLER_0_227_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27164_ _11972_ _11984_ VGND VGND VPWR VPWR _11988_ sky130_fd_sc_hd__and2_1
X_20608_ datamem.data_ram\[40\]\[13\] _06807_ _06731_ datamem.data_ram\[43\]\[13\]
+ VGND VGND VPWR VPWR _07899_ sky130_fd_sc_hd__o22a_1
XFILLER_0_145_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24376_ _09230_ VGND VGND VPWR VPWR _10366_ sky130_fd_sc_hd__buf_8
XFILLER_0_35_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21588_ _08569_ VGND VGND VPWR VPWR _08840_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_61_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26115_ net1675 _11386_ VGND VGND VPWR VPWR _11393_ sky130_fd_sc_hd__and2_1
X_27095_ _11827_ _11941_ VGND VGND VPWR VPWR _11944_ sky130_fd_sc_hd__and2_1
X_20539_ _07823_ datamem.data_ram\[6\]\[21\] datamem.data_ram\[7\]\[21\] _07829_ VGND
+ VGND VPWR VPWR _07830_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26046_ _10209_ _10921_ _10922_ VGND VGND VPWR VPWR _11351_ sky130_fd_sc_hd__and3_2
X_23258_ clknet_1_0__leaf__10108_ VGND VGND VPWR VPWR _10128_ sky130_fd_sc_hd__buf_1
Xclkbuf_leaf_227_clk clknet_5_21__leaf_clk VGND VGND VPWR VPWR clknet_leaf_227_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_63_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22209_ _09377_ VGND VGND VPWR VPWR _01121_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23189_ _10113_ _10114_ _09361_ VGND VGND VPWR VPWR _10115_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_197_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29805_ net1143 _01540_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[1\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_1184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27997_ _12458_ net2948 net76 VGND VGND VPWR VPWR _12459_ sky130_fd_sc_hd__mux2_1
XFILLER_0_218_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14962_ _13509_ _13510_ VGND VGND VPWR VPWR _13511_ sky130_fd_sc_hd__nor2_1
X_29736_ net1082 _01471_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[21\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_17750_ _05150_ VGND VGND VPWR VPWR _01166_ sky130_fd_sc_hd__clkbuf_1
Xhold7 rvcpu.dp.plde.PCPlus4E\[2\] VGND VGND VPWR VPWR net1157 sky130_fd_sc_hd__dlygate4sd3_1
X_26948_ _11825_ _11854_ VGND VGND VPWR VPWR _11856_ sky130_fd_sc_hd__and2_1
XFILLER_0_55_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16701_ _04594_ VGND VGND VPWR VPWR _01691_ sky130_fd_sc_hd__clkbuf_1
X_14893_ _13358_ _13443_ VGND VGND VPWR VPWR _13444_ sky130_fd_sc_hd__nand2_1
X_29667_ net1013 _01402_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[24\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_17681_ net2552 _13271_ _05104_ VGND VGND VPWR VPWR _05114_ sky130_fd_sc_hd__mux2_1
XFILLER_0_226_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26879_ _11795_ net1503 _11809_ _11811_ VGND VGND VPWR VPWR _03357_ sky130_fd_sc_hd__a31o_1
X_19420_ _06715_ VGND VGND VPWR VPWR _06716_ sky130_fd_sc_hd__clkbuf_8
X_28618_ _10777_ _12612_ _12795_ VGND VGND VPWR VPWR _12805_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_18_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16632_ _14164_ net2373 _04551_ VGND VGND VPWR VPWR _04558_ sky130_fd_sc_hd__mux2_1
XFILLER_0_226_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_394 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29598_ net952 _01333_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[25\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19351_ _06646_ VGND VGND VPWR VPWR _06647_ sky130_fd_sc_hd__buf_6
X_16563_ _14164_ net3038 _04514_ VGND VGND VPWR VPWR _04521_ sky130_fd_sc_hd__mux2_1
X_23874__435 clknet_1_0__leaf__10221_ VGND VGND VPWR VPWR net561 sky130_fd_sc_hd__inv_2
X_28549_ _10141_ _12602_ _12668_ VGND VGND VPWR VPWR _12768_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_57_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18302_ _05384_ _05385_ VGND VGND VPWR VPWR _05667_ sky130_fd_sc_hd__nand2_2
XFILLER_0_70_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15514_ _13409_ _13310_ _13617_ _14040_ VGND VGND VPWR VPWR _14041_ sky130_fd_sc_hd__a31o_1
XFILLER_0_169_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31560_ clknet_leaf_71_clk datamem.rd_data_mem\[10\] VGND VGND VPWR VPWR rvcpu.dp.plmw.ReadDataW\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_1319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19282_ _06579_ VGND VGND VPWR VPWR _04449_ sky130_fd_sc_hd__clkbuf_1
X_16494_ _04484_ VGND VGND VPWR VPWR _01796_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_216_5680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_216_5691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15445_ _13374_ _13974_ _13975_ _13412_ VGND VGND VPWR VPWR _13976_ sky130_fd_sc_hd__o211a_1
X_18233_ _05346_ _05595_ _05597_ VGND VGND VPWR VPWR _05598_ sky130_fd_sc_hd__o21a_1
XFILLER_0_154_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30511_ clknet_leaf_197_clk _02246_ VGND VGND VPWR VPWR datamem.data_ram\[56\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_31491_ clknet_leaf_46_clk rvcpu.dp.lAuiPCE\[17\] VGND VGND VPWR VPWR rvcpu.dp.plem.lAuiPCM\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_212_5577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30442_ net780 _02177_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[29\]\[21\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_212_5588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15376_ _13909_ _13471_ _13690_ VGND VGND VPWR VPWR _13910_ sky130_fd_sc_hd__or3_1
XFILLER_0_143_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18164_ _05527_ _05528_ VGND VGND VPWR VPWR _05529_ sky130_fd_sc_hd__and2_1
XFILLER_0_136_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23653__253 clknet_1_1__leaf__10181_ VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__inv_2
XFILLER_0_142_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17115_ _14170_ net2606 _04804_ VGND VGND VPWR VPWR _04814_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18095_ rvcpu.dp.plde.RD1E\[22\] _05292_ _05462_ VGND VGND VPWR VPWR _05463_ sky130_fd_sc_hd__o21a_2
X_30373_ net719 _02108_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[3\]\[24\] sky130_fd_sc_hd__dfxtp_1
Xmax_cap104 _09228_ VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__buf_8
Xhold407 datamem.data_ram\[35\]\[6\] VGND VGND VPWR VPWR net1557 sky130_fd_sc_hd__dlygate4sd3_1
Xhold418 datamem.data_ram\[56\]\[0\] VGND VGND VPWR VPWR net1568 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32112_ clknet_leaf_116_clk _03534_ VGND VGND VPWR VPWR datamem.data_ram\[58\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_17046_ _04777_ VGND VGND VPWR VPWR _01513_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_225_5905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold429 datamem.data_ram\[33\]\[5\] VGND VGND VPWR VPWR net1579 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_146_4005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_218_clk clknet_5_21__leaf_clk VGND VGND VPWR VPWR clknet_leaf_218_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_96_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32043_ clknet_leaf_130_clk _03465_ VGND VGND VPWR VPWR datamem.data_ram\[49\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18997_ _06313_ _06096_ _06331_ _05658_ VGND VGND VPWR VPWR _06332_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_225_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_163_4396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1107 datamem.data_ram\[57\]\[25\] VGND VGND VPWR VPWR net2257 sky130_fd_sc_hd__dlygate4sd3_1
X_17948_ rvcpu.dp.plde.RD1E\[13\] _05266_ _05270_ _13237_ _05319_ VGND VGND VPWR VPWR
+ _05320_ sky130_fd_sc_hd__a221o_2
Xhold1118 datamem.data_ram\[40\]\[26\] VGND VGND VPWR VPWR net2268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1129 rvcpu.dp.rf.reg_file_arr\[8\]\[9\] VGND VGND VPWR VPWR net2279 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_105_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_77_Left_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_105_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32945_ clknet_leaf_215_clk _04367_ VGND VGND VPWR VPWR datamem.data_ram\[6\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17879_ _05244_ _05247_ _05251_ VGND VGND VPWR VPWR _05252_ sky130_fd_sc_hd__nand3_2
XFILLER_0_221_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_176_4713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19618_ _06586_ _06580_ VGND VGND VPWR VPWR _06914_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_176_4724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32876_ clknet_leaf_56_clk _04298_ VGND VGND VPWR VPWR datamem.data_ram\[10\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20890_ _06753_ _08168_ _08172_ _08179_ VGND VGND VPWR VPWR _08180_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_66_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31827_ clknet_leaf_105_clk _03281_ VGND VGND VPWR VPWR datamem.data_ram\[16\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19549_ datamem.data_ram\[18\]\[24\] _06803_ _06731_ datamem.data_ram\[19\]\[24\]
+ _06733_ VGND VGND VPWR VPWR _06845_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_66_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22560_ _09412_ _09708_ _09710_ _09712_ _09413_ VGND VGND VPWR VPWR _09713_ sky130_fd_sc_hd__a221o_1
X_31758_ clknet_leaf_17_clk _03212_ VGND VGND VPWR VPWR rvcpu.dp.plde.ALUSrcE sky130_fd_sc_hd__dfxtp_2
XFILLER_0_119_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21511_ _08686_ _08765_ _08748_ VGND VGND VPWR VPWR _08766_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_174_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30709_ clknet_leaf_148_clk _02444_ VGND VGND VPWR VPWR datamem.data_ram\[49\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_683 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22491_ rvcpu.dp.rf.reg_file_arr\[4\]\[9\] rvcpu.dp.rf.reg_file_arr\[5\]\[9\] rvcpu.dp.rf.reg_file_arr\[6\]\[9\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[9\] _09478_ _09479_ VGND VGND VPWR VPWR _09648_ sky130_fd_sc_hd__mux4_1
X_31689_ clknet_leaf_37_clk _03147_ VGND VGND VPWR VPWR rvcpu.dp.pcreg.q\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_3731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_3742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24230_ _09256_ net4103 _10279_ VGND VGND VPWR VPWR _10286_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21442_ _08692_ _08694_ _08698_ _08700_ VGND VGND VPWR VPWR _08701_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_86_Left_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_131_3628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_3639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_226_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21373_ _08630_ _08633_ _08541_ VGND VGND VPWR VPWR _08634_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_872 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20324_ datamem.data_ram\[18\]\[4\] _06989_ _06921_ datamem.data_ram\[21\]\[4\] VGND
+ VGND VPWR VPWR _07616_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_9_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold930 rvcpu.dp.rf.reg_file_arr\[1\]\[31\] VGND VGND VPWR VPWR net2080 sky130_fd_sc_hd__dlygate4sd3_1
Xhold941 datamem.data_ram\[26\]\[23\] VGND VGND VPWR VPWR net2091 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold952 rvcpu.dp.rf.reg_file_arr\[11\]\[8\] VGND VGND VPWR VPWR net2102 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_209_clk clknet_5_22__leaf_clk VGND VGND VPWR VPWR clknet_leaf_209_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold963 datamem.data_ram\[35\]\[13\] VGND VGND VPWR VPWR net2113 sky130_fd_sc_hd__dlygate4sd3_1
X_27920_ _12411_ VGND VGND VPWR VPWR _03798_ sky130_fd_sc_hd__clkbuf_1
X_20255_ datamem.data_ram\[45\]\[3\] _06920_ _06961_ datamem.data_ram\[43\]\[3\] _07547_
+ VGND VGND VPWR VPWR _07548_ sky130_fd_sc_hd__a221o_1
Xhold3010 datamem.data_ram\[60\]\[16\] VGND VGND VPWR VPWR net4160 sky130_fd_sc_hd__dlygate4sd3_1
Xhold974 rvcpu.dp.rf.reg_file_arr\[4\]\[11\] VGND VGND VPWR VPWR net2124 sky130_fd_sc_hd__dlygate4sd3_1
Xhold985 rvcpu.dp.rf.reg_file_arr\[5\]\[1\] VGND VGND VPWR VPWR net2135 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold996 rvcpu.dp.rf.reg_file_arr\[18\]\[22\] VGND VGND VPWR VPWR net2146 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3021 datamem.data_ram\[45\]\[10\] VGND VGND VPWR VPWR net4171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3032 rvcpu.dp.rf.reg_file_arr\[12\]\[13\] VGND VGND VPWR VPWR net4182 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_34_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27851_ _12125_ net2385 _12373_ VGND VGND VPWR VPWR _12374_ sky130_fd_sc_hd__mux2_1
X_20186_ datamem.data_ram\[5\]\[11\] _06768_ _06760_ datamem.data_ram\[7\]\[11\] _07478_
+ VGND VGND VPWR VPWR _07479_ sky130_fd_sc_hd__o221a_1
Xhold3043 datamem.data_ram\[19\]\[31\] VGND VGND VPWR VPWR net4193 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3054 datamem.data_ram\[29\]\[18\] VGND VGND VPWR VPWR net4204 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2320 datamem.data_ram\[37\]\[28\] VGND VGND VPWR VPWR net3470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3065 datamem.data_ram\[7\]\[28\] VGND VGND VPWR VPWR net4215 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2331 datamem.data_ram\[19\]\[23\] VGND VGND VPWR VPWR net3481 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26802_ _11681_ _11762_ VGND VGND VPWR VPWR _11765_ sky130_fd_sc_hd__and2_1
Xhold3076 rvcpu.dp.rf.reg_file_arr\[20\]\[5\] VGND VGND VPWR VPWR net4226 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_95_Left_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2342 rvcpu.dp.rf.reg_file_arr\[15\]\[19\] VGND VGND VPWR VPWR net3492 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3087 rvcpu.dp.rf.reg_file_arr\[26\]\[19\] VGND VGND VPWR VPWR net4237 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3098 rvcpu.dp.rf.reg_file_arr\[24\]\[27\] VGND VGND VPWR VPWR net4248 sky130_fd_sc_hd__dlygate4sd3_1
X_24994_ _10444_ net3804 _10715_ VGND VGND VPWR VPWR _10718_ sky130_fd_sc_hd__mux2_1
X_27782_ _12091_ net4433 _12326_ VGND VGND VPWR VPWR _12332_ sky130_fd_sc_hd__mux2_1
Xhold2353 datamem.data_ram\[3\]\[30\] VGND VGND VPWR VPWR net3503 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2364 rvcpu.dp.rf.reg_file_arr\[25\]\[18\] VGND VGND VPWR VPWR net3514 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2375 datamem.data_ram\[30\]\[21\] VGND VGND VPWR VPWR net3525 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1630 datamem.data_ram\[22\]\[26\] VGND VGND VPWR VPWR net2780 sky130_fd_sc_hd__dlygate4sd3_1
X_29521_ net883 _01256_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[28\]\[28\] sky130_fd_sc_hd__dfxtp_1
Xhold1641 datamem.data_ram\[43\]\[29\] VGND VGND VPWR VPWR net2791 sky130_fd_sc_hd__dlygate4sd3_1
X_26733_ _11722_ VGND VGND VPWR VPWR _03300_ sky130_fd_sc_hd__clkbuf_1
Xhold2386 rvcpu.dp.rf.reg_file_arr\[27\]\[13\] VGND VGND VPWR VPWR net3536 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1652 datamem.data_ram\[37\]\[21\] VGND VGND VPWR VPWR net2802 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2397 datamem.data_ram\[32\]\[11\] VGND VGND VPWR VPWR net3547 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1663 datamem.data_ram\[4\]\[8\] VGND VGND VPWR VPWR net2813 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1674 rvcpu.dp.rf.reg_file_arr\[16\]\[20\] VGND VGND VPWR VPWR net2824 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1685 rvcpu.dp.rf.reg_file_arr\[0\]\[12\] VGND VGND VPWR VPWR net2835 sky130_fd_sc_hd__dlygate4sd3_1
X_26664_ _11665_ net1853 _11675_ _11682_ VGND VGND VPWR VPWR _03271_ sky130_fd_sc_hd__a31o_1
XFILLER_0_212_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_193_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1696 datamem.data_ram\[42\]\[27\] VGND VGND VPWR VPWR net2846 sky130_fd_sc_hd__dlygate4sd3_1
X_29452_ net814 _01187_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[30\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0__10264_ _10264_ VGND VGND VPWR VPWR clknet_0__10264_ sky130_fd_sc_hd__clkbuf_16
X_28403_ _12178_ _12622_ _12668_ VGND VGND VPWR VPWR _12678_ sky130_fd_sc_hd__a21oi_4
X_25615_ _10735_ net3459 net53 VGND VGND VPWR VPWR _11072_ sky130_fd_sc_hd__mux2_1
XFILLER_0_212_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22827_ rvcpu.dp.rf.reg_file_arr\[12\]\[27\] rvcpu.dp.rf.reg_file_arr\[13\]\[27\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[27\] rvcpu.dp.rf.reg_file_arr\[15\]\[27\] _09462_
+ _09721_ VGND VGND VPWR VPWR _09966_ sky130_fd_sc_hd__mux4_1
X_26595_ _11618_ net1763 _11639_ _11644_ VGND VGND VPWR VPWR _03240_ sky130_fd_sc_hd__a31o_1
X_29383_ clknet_leaf_267_clk _01118_ VGND VGND VPWR VPWR datamem.data_ram\[60\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25546_ _11031_ VGND VGND VPWR VPWR _02804_ sky130_fd_sc_hd__clkbuf_1
X_28334_ _10668_ _12612_ _12573_ VGND VGND VPWR VPWR _12641_ sky130_fd_sc_hd__a21oi_4
Xclkbuf_0__10195_ _10195_ VGND VGND VPWR VPWR clknet_0__10195_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22758_ _09705_ _09892_ _09896_ _09900_ VGND VGND VPWR VPWR _09901_ sky130_fd_sc_hd__and4_1
XFILLER_0_67_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21709_ _08952_ _08953_ _08743_ VGND VGND VPWR VPWR _08954_ sky130_fd_sc_hd__mux2_1
X_28265_ _12355_ net3226 _12603_ VGND VGND VPWR VPWR _12604_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25477_ _07808_ _10043_ _10600_ VGND VGND VPWR VPWR _10995_ sky130_fd_sc_hd__nor3_1
XFILLER_0_54_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22689_ _09398_ _09834_ VGND VGND VPWR VPWR _09835_ sky130_fd_sc_hd__or2_1
XFILLER_0_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_229_6005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_229_6016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15230_ _13767_ _13559_ VGND VGND VPWR VPWR _13771_ sky130_fd_sc_hd__or2_1
XFILLER_0_152_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27216_ _09299_ _11112_ _11898_ VGND VGND VPWR VPWR _12019_ sky130_fd_sc_hd__and3_1
X_24428_ _10396_ net4388 _10386_ VGND VGND VPWR VPWR _10397_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_229_6027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28196_ _12450_ net4072 net46 VGND VGND VPWR VPWR _12566_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15161_ _13429_ _13703_ _13541_ _13664_ _13704_ VGND VGND VPWR VPWR _13705_ sky130_fd_sc_hd__a311o_1
X_27147_ _11976_ _11966_ VGND VGND VPWR VPWR _11977_ sky130_fd_sc_hd__and2_1
XFILLER_0_152_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24359_ _09226_ _10327_ _10269_ VGND VGND VPWR VPWR _10357_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_105_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27078_ _11837_ _11924_ VGND VGND VPWR VPWR _11932_ sky130_fd_sc_hd__and2_1
X_15092_ _13618_ _13620_ _13624_ _13637_ VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__o31a_1
XFILLER_0_132_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26029_ _11121_ net1518 _11339_ _11341_ VGND VGND VPWR VPWR _02977_ sky130_fd_sc_hd__a31o_1
X_18920_ _05536_ _05785_ _05727_ _05537_ VGND VGND VPWR VPWR _06260_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_24_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18851_ _05481_ _06194_ VGND VGND VPWR VPWR _06195_ sky130_fd_sc_hd__xor2_1
X_17802_ _05194_ VGND VGND VPWR VPWR _05195_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_219_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18782_ _06122_ _06130_ VGND VGND VPWR VPWR _06131_ sky130_fd_sc_hd__or2_1
X_23683__279 clknet_1_0__leaf__10194_ VGND VGND VPWR VPWR net405 sky130_fd_sc_hd__inv_2
XFILLER_0_98_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15994_ net1978 _13248_ _14333_ VGND VGND VPWR VPWR _14335_ sky130_fd_sc_hd__mux2_1
XFILLER_0_174_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29719_ net1065 _01454_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[22\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_17733_ _13248_ net2711 _05140_ VGND VGND VPWR VPWR _05142_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14945_ _13297_ _13348_ VGND VGND VPWR VPWR _13494_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30991_ clknet_leaf_102_clk _02726_ VGND VGND VPWR VPWR datamem.data_ram\[13\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_215_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32730_ clknet_leaf_87_clk _04152_ VGND VGND VPWR VPWR datamem.data_ram\[16\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_17664_ _05105_ VGND VGND VPWR VPWR _01207_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_218_5720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14876_ _13313_ _13283_ VGND VGND VPWR VPWR _13428_ sky130_fd_sc_hd__nor2_2
XFILLER_0_106_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_218_5731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19403_ _06655_ VGND VGND VPWR VPWR _06699_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_58_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16615_ _14147_ net4044 _04540_ VGND VGND VPWR VPWR _04549_ sky130_fd_sc_hd__mux2_1
XFILLER_0_187_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32661_ clknet_leaf_79_clk _04083_ VGND VGND VPWR VPWR datamem.data_ram\[19\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17595_ _13244_ net4150 _05068_ VGND VGND VPWR VPWR _05069_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_214_5628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31612_ clknet_leaf_25_clk net1171 VGND VGND VPWR VPWR rvcpu.dp.plmw.PCPlus4W\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19334_ _06629_ VGND VGND VPWR VPWR _06630_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_214_5639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_171_4610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16546_ _14147_ net4153 _04503_ VGND VGND VPWR VPWR _04512_ sky130_fd_sc_hd__mux2_1
XFILLER_0_174_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32592_ clknet_leaf_171_clk _04014_ VGND VGND VPWR VPWR datamem.data_ram\[21\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_23123__800 clknet_1_1__leaf__10105_ VGND VGND VPWR VPWR net926 sky130_fd_sc_hd__inv_2
XFILLER_0_174_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19265_ _05655_ _05743_ _06565_ _05281_ VGND VGND VPWR VPWR _00002_ sky130_fd_sc_hd__a2bb2o_1
X_31543_ clknet_leaf_15_clk net1273 VGND VGND VPWR VPWR rvcpu.dp.plem.RdM\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16477_ _04475_ VGND VGND VPWR VPWR _01804_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_171_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_215_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18216_ _05579_ _05580_ VGND VGND VPWR VPWR _05581_ sky130_fd_sc_hd__nand2_1
X_15428_ _13303_ _13321_ _13454_ VGND VGND VPWR VPWR _13959_ sky130_fd_sc_hd__or3_1
XFILLER_0_128_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31474_ clknet_leaf_66_clk rvcpu.dp.lAuiPCE\[0\] VGND VGND VPWR VPWR rvcpu.dp.plem.lAuiPCM\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_19196_ _06506_ VGND VGND VPWR VPWR rvcpu.dp.lAuiPCE\[22\] sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_198_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15359_ _13358_ _13545_ _13758_ _13893_ _13441_ VGND VGND VPWR VPWR _13894_ sky130_fd_sc_hd__a311o_1
X_18147_ _05510_ _05511_ VGND VGND VPWR VPWR _05512_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30425_ net763 _02160_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[29\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_223_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold204 datamem.data_ram\[28\]\[6\] VGND VGND VPWR VPWR net1354 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_169_4550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold215 _02915_ VGND VGND VPWR VPWR net1365 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_169_4561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold226 rvcpu.dp.plfd.PCPlus4D\[11\] VGND VGND VPWR VPWR net1376 sky130_fd_sc_hd__dlygate4sd3_1
X_18078_ rvcpu.dp.plde.RD1E\[11\] _05266_ _05270_ _13243_ _05407_ VGND VGND VPWR VPWR
+ _05446_ sky130_fd_sc_hd__a221o_2
X_30356_ net702 _02091_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[3\]\[7\] sky130_fd_sc_hd__dfxtp_1
Xhold237 datamem.data_ram\[19\]\[7\] VGND VGND VPWR VPWR net1387 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_223_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold248 datamem.data_ram\[38\]\[3\] VGND VGND VPWR VPWR net1398 sky130_fd_sc_hd__dlygate4sd3_1
Xhold259 datamem.data_ram\[39\]\[4\] VGND VGND VPWR VPWR net1409 sky130_fd_sc_hd__dlygate4sd3_1
X_17029_ net2839 _14442_ _04768_ VGND VGND VPWR VPWR _04769_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_165_4447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30287_ net633 _02022_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[5\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_165_4458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20040_ datamem.data_ram\[6\]\[26\] _06744_ _06765_ datamem.data_ram\[4\]\[26\] VGND
+ VGND VPWR VPWR _07334_ sky130_fd_sc_hd__o22a_1
X_32026_ clknet_leaf_128_clk _03448_ VGND VGND VPWR VPWR datamem.data_ram\[26\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21991_ _09220_ VGND VGND VPWR VPWR _09221_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_68_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23210__861 clknet_1_0__leaf__10112_ VGND VGND VPWR VPWR net987 sky130_fd_sc_hd__inv_2
XFILLER_0_212_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_124_3465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_3476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20942_ datamem.data_ram\[59\]\[22\] _07851_ _06934_ datamem.data_ram\[57\]\[22\]
+ VGND VGND VPWR VPWR _08232_ sky130_fd_sc_hd__o22a_1
X_32928_ clknet_leaf_3_clk _04350_ VGND VGND VPWR VPWR datamem.data_ram\[0\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32859_ clknet_leaf_55_clk _04281_ VGND VGND VPWR VPWR datamem.data_ram\[11\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_20873_ datamem.data_ram\[54\]\[14\] _06683_ _08160_ _08162_ VGND VGND VPWR VPWR
+ _08163_ sky130_fd_sc_hd__o211a_1
XFILLER_0_49_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25400_ _10413_ _10950_ VGND VGND VPWR VPWR _10955_ sky130_fd_sc_hd__and2_1
XFILLER_0_166_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22612_ rvcpu.dp.rf.reg_file_arr\[20\]\[16\] rvcpu.dp.rf.reg_file_arr\[21\]\[16\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[16\] rvcpu.dp.rf.reg_file_arr\[23\]\[16\] _09517_
+ _09577_ VGND VGND VPWR VPWR _09762_ sky130_fd_sc_hd__mux4_2
XFILLER_0_7_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26380_ _13328_ _11268_ _11523_ _11527_ _10041_ VGND VGND VPWR VPWR _03142_ sky130_fd_sc_hd__o221a_1
XFILLER_0_152_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_220_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25331_ _10911_ VGND VGND VPWR VPWR _02709_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_27_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_1302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22543_ rvcpu.dp.rf.reg_file_arr\[4\]\[12\] rvcpu.dp.rf.reg_file_arr\[5\]\[12\] rvcpu.dp.rf.reg_file_arr\[6\]\[12\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[12\] _09604_ _09424_ VGND VGND VPWR VPWR _09697_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_107_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28050_ _12488_ VGND VGND VPWR VPWR _03851_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_98_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25262_ _10538_ net1404 _10867_ _10872_ VGND VGND VPWR VPWR _02679_ sky130_fd_sc_hd__a31o_1
XFILLER_0_9_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22474_ _09389_ _09621_ _09626_ _09631_ VGND VGND VPWR VPWR _09632_ sky130_fd_sc_hd__and4_1
XFILLER_0_161_422 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27001_ _09299_ _10921_ _10922_ VGND VGND VPWR VPWR _11886_ sky130_fd_sc_hd__and3_1
XFILLER_0_173_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24213_ _09326_ net4029 _10270_ VGND VGND VPWR VPWR _10277_ sky130_fd_sc_hd__mux2_1
X_21425_ _08560_ VGND VGND VPWR VPWR _08684_ sky130_fd_sc_hd__buf_4
XFILLER_0_17_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25193_ _10834_ VGND VGND VPWR VPWR _02648_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21356_ _08615_ _08616_ rvcpu.ALUResultE\[31\] _08617_ VGND VGND VPWR VPWR _08618_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_142_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_188_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20307_ _07599_ VGND VGND VPWR VPWR _04440_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_198_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24075_ _10209_ _09269_ _09361_ VGND VGND VPWR VPWR _10249_ sky130_fd_sc_hd__a21oi_4
X_28952_ _12743_ net3691 net67 VGND VGND VPWR VPWR _12983_ sky130_fd_sc_hd__mux2_1
X_21287_ _08548_ VGND VGND VPWR VPWR _08549_ sky130_fd_sc_hd__buf_6
Xhold760 rvcpu.dp.rf.reg_file_arr\[19\]\[4\] VGND VGND VPWR VPWR net1910 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold771 datamem.data_ram\[59\]\[26\] VGND VGND VPWR VPWR net1921 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold782 rvcpu.dp.rf.reg_file_arr\[12\]\[2\] VGND VGND VPWR VPWR net1932 sky130_fd_sc_hd__dlygate4sd3_1
X_27903_ _12391_ net1384 _12393_ _12402_ VGND VGND VPWR VPWR _03790_ sky130_fd_sc_hd__a31o_1
X_23825__407 clknet_1_0__leaf__10208_ VGND VGND VPWR VPWR net533 sky130_fd_sc_hd__inv_2
XFILLER_0_229_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20238_ datamem.data_ram\[52\]\[3\] _06954_ _06947_ datamem.data_ram\[49\]\[3\] VGND
+ VGND VPWR VPWR _07531_ sky130_fd_sc_hd__a22o_1
Xhold793 rvcpu.dp.rf.reg_file_arr\[1\]\[7\] VGND VGND VPWR VPWR net1943 sky130_fd_sc_hd__dlygate4sd3_1
X_28883_ _12760_ net2797 _12941_ VGND VGND VPWR VPWR _12946_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27834_ _12362_ VGND VGND VPWR VPWR _03761_ sky130_fd_sc_hd__clkbuf_1
X_20169_ datamem.data_ram\[26\]\[11\] _06754_ _06697_ datamem.data_ram\[24\]\[11\]
+ VGND VGND VPWR VPWR _07462_ sky130_fd_sc_hd__o22a_1
XFILLER_0_200_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2150 datamem.data_ram\[18\]\[25\] VGND VGND VPWR VPWR net3300 sky130_fd_sc_hd__dlygate4sd3_1
X_23905__464 clknet_1_1__leaf__10223_ VGND VGND VPWR VPWR net590 sky130_fd_sc_hd__inv_2
XFILLER_0_217_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_607 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2161 datamem.data_ram\[54\]\[29\] VGND VGND VPWR VPWR net3311 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2172 rvcpu.dp.rf.reg_file_arr\[31\]\[29\] VGND VGND VPWR VPWR net3322 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2183 datamem.data_ram\[34\]\[25\] VGND VGND VPWR VPWR net3333 sky130_fd_sc_hd__dlygate4sd3_1
X_27765_ _12322_ VGND VGND VPWR VPWR _03732_ sky130_fd_sc_hd__clkbuf_1
Xhold2194 datamem.data_ram\[15\]\[8\] VGND VGND VPWR VPWR net3344 sky130_fd_sc_hd__dlygate4sd3_1
X_24977_ _10470_ net2670 net101 VGND VGND VPWR VPWR _10709_ sky130_fd_sc_hd__mux2_1
Xhold1460 datamem.data_ram\[9\]\[19\] VGND VGND VPWR VPWR net2610 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29504_ net866 _01239_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[28\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14730_ rvcpu.dp.pcreg.q\[6\] VGND VGND VPWR VPWR _13283_ sky130_fd_sc_hd__inv_2
X_26716_ _10500_ VGND VGND VPWR VPWR _11713_ sky130_fd_sc_hd__buf_8
Xhold1471 rvcpu.dp.rf.reg_file_arr\[31\]\[4\] VGND VGND VPWR VPWR net2621 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1482 rvcpu.dp.rf.reg_file_arr\[20\]\[1\] VGND VGND VPWR VPWR net2632 sky130_fd_sc_hd__dlygate4sd3_1
X_27696_ _12136_ net3573 _12280_ VGND VGND VPWR VPWR _12286_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1493 rvcpu.dp.rf.reg_file_arr\[4\]\[30\] VGND VGND VPWR VPWR net2643 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14661_ _13230_ VGND VGND VPWR VPWR _03188_ sky130_fd_sc_hd__clkbuf_1
X_29435_ net797 _01170_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[30\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_26647_ _11665_ net1743 _11662_ _11670_ VGND VGND VPWR VPWR _03266_ sky130_fd_sc_hd__a31o_1
XFILLER_0_196_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_211_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16400_ net1912 _14430_ _14561_ VGND VGND VPWR VPWR _14566_ sky130_fd_sc_hd__mux2_1
Xclkbuf_0__10247_ _10247_ VGND VGND VPWR VPWR clknet_0__10247_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_131_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23719__312 clknet_1_0__leaf__10197_ VGND VGND VPWR VPWR net438 sky130_fd_sc_hd__inv_2
X_14592_ _13174_ _13175_ _13176_ VGND VGND VPWR VPWR _13177_ sky130_fd_sc_hd__or3_4
X_17380_ _14162_ net2435 _04949_ VGND VGND VPWR VPWR _04955_ sky130_fd_sc_hd__mux2_1
X_29366_ clknet_leaf_208_clk _01101_ VGND VGND VPWR VPWR datamem.data_ram\[60\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_26578_ _11634_ VGND VGND VPWR VPWR _03233_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_211_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16331_ _14529_ VGND VGND VPWR VPWR _01872_ sky130_fd_sc_hd__clkbuf_1
X_28317_ _10668_ _12602_ _12573_ VGND VGND VPWR VPWR _12632_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_95_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__10178_ _10178_ VGND VGND VPWR VPWR clknet_0__10178_ sky130_fd_sc_hd__clkbuf_16
X_25529_ _11022_ VGND VGND VPWR VPWR _02796_ sky130_fd_sc_hd__clkbuf_1
X_29297_ clknet_leaf_6_clk _01032_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD1E\[4\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__10078_ clknet_0__10078_ VGND VGND VPWR VPWR clknet_1_1__leaf__10078_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_125_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19050_ _06378_ VGND VGND VPWR VPWR rvcpu.dp.lAuiPCE\[4\] sky130_fd_sc_hd__clkbuf_1
X_16262_ net4276 _14428_ _14489_ VGND VGND VPWR VPWR _14493_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28248_ _12450_ net2844 net44 VGND VGND VPWR VPWR _12594_ sky130_fd_sc_hd__mux2_1
X_15213_ _13290_ _13444_ VGND VGND VPWR VPWR _13755_ sky130_fd_sc_hd__nand2_1
X_18001_ rvcpu.dp.plem.ALUResultM\[3\] VGND VGND VPWR VPWR _05371_ sky130_fd_sc_hd__inv_4
XFILLER_0_36_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16193_ _13219_ VGND VGND VPWR VPWR _14447_ sky130_fd_sc_hd__buf_4
X_28179_ _12433_ net3388 _12555_ VGND VGND VPWR VPWR _12557_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15144_ _13683_ _13684_ _13686_ _13687_ _13439_ VGND VGND VPWR VPWR _13688_ sky130_fd_sc_hd__a41o_1
X_30210_ net564 _01945_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[8\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_31190_ clknet_leaf_38_clk _02893_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCPlus4D\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_205_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30141_ net503 _01876_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[0\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_15075_ _13301_ _13562_ _13359_ VGND VGND VPWR VPWR _13621_ sky130_fd_sc_hd__a21o_1
X_19952_ datamem.data_ram\[50\]\[18\] _06692_ _07240_ _07245_ VGND VGND VPWR VPWR
+ _07246_ sky130_fd_sc_hd__o211a_1
XFILLER_0_26_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23153__826 clknet_1_0__leaf__10109_ VGND VGND VPWR VPWR net952 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_207_5454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_207_5465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18903_ _05459_ _05732_ _05730_ _05458_ VGND VGND VPWR VPWR _06244_ sky130_fd_sc_hd__a2bb2o_1
X_30072_ net434 _01807_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[12\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19883_ _07170_ _07175_ _07177_ VGND VGND VPWR VPWR _07178_ sky130_fd_sc_hd__a21o_1
X_23765__354 clknet_1_1__leaf__10201_ VGND VGND VPWR VPWR net480 sky130_fd_sc_hd__inv_2
XFILLER_0_207_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_208_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_5_27__f_clk clknet_2_3_0_clk VGND VGND VPWR VPWR clknet_5_27__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_18834_ _05866_ _05864_ _06179_ VGND VGND VPWR VPWR _06180_ sky130_fd_sc_hd__o21a_1
XFILLER_0_207_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_160_4333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_160_4344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_5266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_5277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18765_ _05698_ _05967_ _06114_ VGND VGND VPWR VPWR _06115_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_175_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15977_ net2123 _13223_ _14322_ VGND VGND VPWR VPWR _14326_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17716_ _13223_ net2158 _05129_ VGND VGND VPWR VPWR _05133_ sky130_fd_sc_hd__mux2_1
X_14928_ _13284_ _13346_ VGND VGND VPWR VPWR _13477_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18696_ _05419_ _05727_ _05974_ _05416_ _06049_ VGND VGND VPWR VPWR _06050_ sky130_fd_sc_hd__a221o_1
X_30974_ clknet_leaf_160_clk _02709_ VGND VGND VPWR VPWR datamem.data_ram\[39\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32713_ clknet_leaf_252_clk _04135_ VGND VGND VPWR VPWR datamem.data_ram\[17\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_63_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17647_ _05096_ VGND VGND VPWR VPWR _01215_ sky130_fd_sc_hd__clkbuf_1
X_14859_ _13407_ _13410_ VGND VGND VPWR VPWR _13411_ sky130_fd_sc_hd__nor2_1
XFILLER_0_175_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_158_4284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32644_ clknet_leaf_153_clk _04066_ VGND VGND VPWR VPWR datamem.data_ram\[1\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_158_4295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17578_ _13220_ net2749 _05057_ VGND VGND VPWR VPWR _05060_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19317_ _06612_ VGND VGND VPWR VPWR _06613_ sky130_fd_sc_hd__buf_6
X_16529_ _04502_ VGND VGND VPWR VPWR _04503_ sky130_fd_sc_hd__clkbuf_4
X_32575_ clknet_leaf_274_clk _03997_ VGND VGND VPWR VPWR datamem.data_ram\[22\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_190_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31526_ clknet_leaf_45_clk net1162 VGND VGND VPWR VPWR rvcpu.dp.plem.PCPlus4M\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_19248_ _06551_ rvcpu.dp.plde.ImmExtE\[29\] _06493_ VGND VGND VPWR VPWR _06552_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19179_ _06490_ _06491_ VGND VGND VPWR VPWR _06492_ sky130_fd_sc_hd__and2_1
X_31457_ clknet_leaf_5_clk rvcpu.dp.SrcBFW_Mux.y\[15\] VGND VGND VPWR VPWR rvcpu.dp.plem.WriteDataM\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_23471__119 clknet_1_0__leaf__10158_ VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__inv_2
XFILLER_0_83_1210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_4509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21210_ _08354_ _08488_ _08471_ VGND VGND VPWR VPWR _08489_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_143_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_93_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30408_ net746 _02143_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[31\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22190_ _09367_ VGND VGND VPWR VPWR _01112_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_112_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31388_ clknet_leaf_37_clk _03091_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCE\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21141_ datamem.data_ram\[58\]\[23\] _06689_ _06729_ datamem.data_ram\[59\]\[23\]
+ _08429_ VGND VGND VPWR VPWR _08430_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_113_3199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30339_ net685 _02074_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[4\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23093__773 clknet_1_0__leaf__10102_ VGND VGND VPWR VPWR net899 sky130_fd_sc_hd__inv_2
X_21072_ datamem.data_ram\[56\]\[7\] _06935_ _06941_ datamem.data_ram\[59\]\[7\] _08360_
+ VGND VGND VPWR VPWR _08361_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23015__719 clknet_1_0__leaf__10086_ VGND VGND VPWR VPWR net845 sky130_fd_sc_hd__inv_2
X_32009_ clknet_leaf_127_clk _03431_ VGND VGND VPWR VPWR datamem.data_ram\[27\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_20023_ datamem.data_ram\[42\]\[2\] _06930_ _06924_ datamem.data_ram\[47\]\[2\] VGND
+ VGND VPWR VPWR _07317_ sky130_fd_sc_hd__a22o_1
X_24900_ _10454_ net4045 _10659_ VGND VGND VPWR VPWR _10667_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_126_3516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25880_ _11153_ VGND VGND VPWR VPWR _11256_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_126_3527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24831_ _10629_ VGND VGND VPWR VPWR _02491_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_198_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24762_ _10468_ net3692 _10589_ VGND VGND VPWR VPWR _10591_ sky130_fd_sc_hd__mux2_1
X_27550_ _12145_ net2936 _12206_ VGND VGND VPWR VPWR _12208_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_87_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21974_ _08540_ _09204_ VGND VGND VPWR VPWR _09205_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_87_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20925_ datamem.data_ram\[44\]\[22\] datamem.data_ram\[45\]\[22\] _07849_ VGND VGND
+ VPWR VPWR _08215_ sky130_fd_sc_hd__mux2_1
X_27481_ _12128_ net2465 _12169_ VGND VGND VPWR VPWR _12171_ sky130_fd_sc_hd__mux2_1
X_24693_ _10442_ net3867 _10552_ VGND VGND VPWR VPWR _10554_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29220_ _11533_ net1458 _13122_ _13129_ VGND VGND VPWR VPWR _04380_ sky130_fd_sc_hd__a31o_1
X_26432_ net1362 _11268_ _11564_ _11565_ _10041_ VGND VGND VPWR VPWR _03156_ sky130_fd_sc_hd__o221a_1
XFILLER_0_178_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23644_ _10188_ VGND VGND VPWR VPWR _01745_ sky130_fd_sc_hd__clkbuf_1
X_20856_ _07635_ datamem.data_ram\[15\]\[14\] _07832_ datamem.data_ram\[14\]\[14\]
+ _07845_ VGND VGND VPWR VPWR _08146_ sky130_fd_sc_hd__a221o_1
XFILLER_0_3_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26363_ _11501_ net1710 _11510_ _11515_ VGND VGND VPWR VPWR _03137_ sky130_fd_sc_hd__a31o_1
XFILLER_0_194_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29151_ _09287_ net3984 _13085_ VGND VGND VPWR VPWR _13092_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20787_ datamem.data_ram\[18\]\[30\] datamem.data_ram\[19\]\[30\] _07835_ VGND VGND
+ VPWR VPWR _08077_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_46_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28102_ _12458_ net3962 net75 VGND VGND VPWR VPWR _12516_ sky130_fd_sc_hd__mux2_1
X_25314_ _10816_ net2984 _10899_ VGND VGND VPWR VPWR _10902_ sky130_fd_sc_hd__mux2_1
X_22526_ rvcpu.dp.rf.reg_file_arr\[0\]\[11\] rvcpu.dp.rf.reg_file_arr\[1\]\[11\] rvcpu.dp.rf.reg_file_arr\[2\]\[11\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[11\] _09463_ _09466_ VGND VGND VPWR VPWR _09681_
+ sky130_fd_sc_hd__mux4_1
X_26294_ net2115 _11478_ VGND VGND VPWR VPWR _11480_ sky130_fd_sc_hd__and2_1
X_29082_ _13055_ VGND VGND VPWR VPWR _04316_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28033_ _12441_ net3064 _12473_ VGND VGND VPWR VPWR _12479_ sky130_fd_sc_hd__mux2_1
X_25245_ _10862_ VGND VGND VPWR VPWR _02672_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22457_ _09511_ _09614_ VGND VGND VPWR VPWR _09615_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_157_Right_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21408_ rvcpu.dp.rf.reg_file_arr\[4\]\[2\] rvcpu.dp.rf.reg_file_arr\[5\]\[2\] rvcpu.dp.rf.reg_file_arr\[6\]\[2\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[2\] _08567_ _08570_ VGND VGND VPWR VPWR _08668_ sky130_fd_sc_hd__mux4_1
X_25176_ _09325_ VGND VGND VPWR VPWR _10824_ sky130_fd_sc_hd__buf_2
X_22388_ _09415_ _09547_ _09549_ VGND VGND VPWR VPWR _09550_ sky130_fd_sc_hd__a21o_1
XFILLER_0_206_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21339_ rvcpu.ALUResultE\[5\] rvcpu.ALUResultE\[6\] rvcpu.ALUResultE\[7\] _08600_
+ VGND VGND VPWR VPWR _08601_ sky130_fd_sc_hd__or4_1
XFILLER_0_124_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29984_ net354 _01719_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[14\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_23217__867 clknet_1_1__leaf__10124_ VGND VGND VPWR VPWR net993 sky130_fd_sc_hd__inv_2
X_28935_ _12973_ VGND VGND VPWR VPWR _04251_ sky130_fd_sc_hd__clkbuf_1
Xhold590 datamem.data_ram\[61\]\[1\] VGND VGND VPWR VPWR net1740 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15900_ net2329 _13210_ _14275_ VGND VGND VPWR VPWR _14285_ sky130_fd_sc_hd__mux2_1
XFILLER_0_194_1006 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28866_ _12696_ net3370 _12932_ VGND VGND VPWR VPWR _12937_ sky130_fd_sc_hd__mux2_1
X_16880_ _04689_ VGND VGND VPWR VPWR _01599_ sky130_fd_sc_hd__clkbuf_1
X_24196__35 clknet_1_0__leaf__10267_ VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__inv_2
XFILLER_0_216_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_202_5340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_218_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_205_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_202_5351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27817_ _12351_ VGND VGND VPWR VPWR _03755_ sky130_fd_sc_hd__clkbuf_1
X_15831_ _14235_ VGND VGND VPWR VPWR _14247_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_204_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_216_275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28797_ _12900_ VGND VGND VPWR VPWR _04186_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18550_ _05585_ _05586_ _05368_ VGND VGND VPWR VPWR _05910_ sky130_fd_sc_hd__a21o_1
X_27748_ _12313_ VGND VGND VPWR VPWR _03724_ sky130_fd_sc_hd__clkbuf_1
X_15762_ _14198_ VGND VGND VPWR VPWR _14210_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_194_5141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_194_5152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_194_5163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1290 rvcpu.dp.rf.reg_file_arr\[28\]\[24\] VGND VGND VPWR VPWR net2440 sky130_fd_sc_hd__dlygate4sd3_1
X_17501_ _13207_ net4299 _05010_ VGND VGND VPWR VPWR _05019_ sky130_fd_sc_hd__mux2_1
XFILLER_0_213_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14713_ net1991 _13269_ _13245_ VGND VGND VPWR VPWR _13270_ sky130_fd_sc_hd__mux2_1
X_18481_ _05768_ _05756_ _05842_ VGND VGND VPWR VPWR _05843_ sky130_fd_sc_hd__o21a_1
XANTENNA_430 _06790_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27679_ _12276_ VGND VGND VPWR VPWR _03692_ sky130_fd_sc_hd__clkbuf_1
X_15693_ _13234_ VGND VGND VPWR VPWR _14166_ sky130_fd_sc_hd__buf_4
XFILLER_0_157_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_441 _07023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_213_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_190_5049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_452 _07860_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29418_ clknet_leaf_12_clk _01153_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD2E\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17432_ _04982_ VGND VGND VPWR VPWR _01324_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_200_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14644_ net2231 _13217_ _13214_ VGND VGND VPWR VPWR _13218_ sky130_fd_sc_hd__mux2_1
XANTENNA_463 _08744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_170_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_474 _09281_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_30690_ clknet_leaf_174_clk _02425_ VGND VGND VPWR VPWR datamem.data_ram\[4\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_485 _09478_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_496 _10044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_184_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29349_ clknet_leaf_144_clk _01084_ VGND VGND VPWR VPWR datamem.data_ram\[61\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_17363_ _14145_ net3878 _04938_ VGND VGND VPWR VPWR _04946_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19102_ _06413_ _06417_ _06414_ VGND VGND VPWR VPWR _06424_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16314_ net2235 _14480_ _14511_ VGND VGND VPWR VPWR _14520_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_153_4170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32360_ clknet_leaf_275_clk _03782_ VGND VGND VPWR VPWR datamem.data_ram\[30\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17294_ _04909_ VGND VGND VPWR VPWR _01397_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31311_ clknet_leaf_46_clk _03014_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCPlus4E\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_19033_ rvcpu.dp.plde.ImmExtE\[0\] rvcpu.dp.plde.PCE\[0\] _06357_ _06363_ VGND VGND
+ VPWR VPWR _06364_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_126_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16245_ _13271_ VGND VGND VPWR VPWR _14482_ sky130_fd_sc_hd__buf_4
X_32291_ clknet_leaf_211_clk _03713_ VGND VGND VPWR VPWR datamem.data_ram\[32\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_124_Right_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_209_5505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_209_5516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31242_ clknet_leaf_34_clk _02945_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCD\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16176_ _14435_ VGND VGND VPWR VPWR _01941_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_112_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15127_ rvcpu.dp.pcreg.q\[6\] _13389_ VGND VGND VPWR VPWR _13672_ sky130_fd_sc_hd__nand2_2
X_31173_ clknet_leaf_228_clk _02876_ VGND VGND VPWR VPWR datamem.data_ram\[5\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_15058_ _13292_ _13604_ _13329_ VGND VGND VPWR VPWR _13605_ sky130_fd_sc_hd__o21a_1
X_19935_ datamem.data_ram\[37\]\[18\] _06703_ _06648_ datamem.data_ram\[32\]\[18\]
+ VGND VGND VPWR VPWR _07229_ sky130_fd_sc_hd__o22a_1
X_30124_ net486 _01859_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[10\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2908 datamem.data_ram\[49\]\[18\] VGND VGND VPWR VPWR net4058 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2919 datamem.data_ram\[11\]\[23\] VGND VGND VPWR VPWR net4069 sky130_fd_sc_hd__dlygate4sd3_1
X_30055_ net417 _01790_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[12\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_19866_ datamem.data_ram\[13\]\[1\] _06969_ _06926_ datamem.data_ram\[15\]\[1\] VGND
+ VGND VPWR VPWR _07161_ sky130_fd_sc_hd__a22o_1
XFILLER_0_177_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18817_ _06155_ _06160_ _06163_ VGND VGND VPWR VPWR _06164_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_128_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19797_ datamem.data_ram\[58\]\[9\] _06611_ _06647_ datamem.data_ram\[56\]\[9\] _06601_
+ VGND VGND VPWR VPWR _07092_ sky130_fd_sc_hd__o221a_1
XFILLER_0_179_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_218_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_121_3402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18748_ _06085_ _05786_ _05784_ _05324_ _06098_ VGND VGND VPWR VPWR _06099_ sky130_fd_sc_hd__o221a_1
XFILLER_0_222_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18679_ _06018_ _05786_ _05784_ _05442_ _06033_ VGND VGND VPWR VPWR _06034_ sky130_fd_sc_hd__o221a_1
X_30957_ clknet_leaf_154_clk _02692_ VGND VGND VPWR VPWR datamem.data_ram\[3\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20710_ datamem.data_ram\[30\]\[5\] _06952_ _06925_ datamem.data_ram\[31\]\[5\] _06679_
+ VGND VGND VPWR VPWR _08001_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_82_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_82_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21690_ rvcpu.dp.rf.reg_file_arr\[20\]\[16\] rvcpu.dp.rf.reg_file_arr\[21\]\[16\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[16\] rvcpu.dp.rf.reg_file_arr\[23\]\[16\] _08778_
+ _08825_ VGND VGND VPWR VPWR _08936_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_82_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30888_ clknet_leaf_223_clk _02623_ VGND VGND VPWR VPWR datamem.data_ram\[42\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32627_ clknet_leaf_93_clk _04049_ VGND VGND VPWR VPWR datamem.data_ram\[1\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_20641_ datamem.data_ram\[16\]\[29\] _06807_ _06789_ datamem.data_ram\[17\]\[29\]
+ VGND VGND VPWR VPWR _07932_ sky130_fd_sc_hd__o22a_1
XFILLER_0_176_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_3342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23322__962 clknet_1_0__leaf__10134_ VGND VGND VPWR VPWR net1088 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_119_3353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32558_ clknet_leaf_244_clk _03980_ VGND VGND VPWR VPWR datamem.data_ram\[22\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_20572_ _07862_ VGND VGND VPWR VPWR _07863_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_190_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22311_ _09452_ VGND VGND VPWR VPWR _09476_ sky130_fd_sc_hd__clkbuf_8
X_31509_ clknet_leaf_52_clk net1174 VGND VGND VPWR VPWR rvcpu.dp.plem.PCPlus4M\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_225_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32489_ clknet_leaf_77_clk _03911_ VGND VGND VPWR VPWR datamem.data_ram\[25\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25030_ _10740_ VGND VGND VPWR VPWR _02579_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22242_ _09394_ VGND VGND VPWR VPWR _09408_ sky130_fd_sc_hd__buf_4
XFILLER_0_104_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_200_Left_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23101__780 clknet_1_0__leaf__10103_ VGND VGND VPWR VPWR net906 sky130_fd_sc_hd__inv_2
XFILLER_0_103_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22173_ _09322_ net2482 _09352_ VGND VGND VPWR VPWR _09358_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__10219_ clknet_0__10219_ VGND VGND VPWR VPWR clknet_1_0__leaf__10219_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_140_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21124_ datamem.data_ram\[40\]\[23\] datamem.data_ram\[41\]\[23\] _07874_ VGND VGND
+ VPWR VPWR _08413_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26981_ _11863_ net1758 _11865_ _11874_ VGND VGND VPWR VPWR _03396_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28720_ _10979_ _12612_ _12795_ VGND VGND VPWR VPWR _12859_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_10_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25932_ _11146_ VGND VGND VPWR VPWR _11286_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21055_ _07866_ _08342_ _08343_ _07862_ VGND VGND VPWR VPWR _08344_ sky130_fd_sc_hd__o22a_1
XFILLER_0_201_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20006_ datamem.data_ram\[58\]\[2\] _06930_ _06924_ datamem.data_ram\[63\]\[2\] VGND
+ VGND VPWR VPWR _07300_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_145_3969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_10__f_clk clknet_2_1_0_clk VGND VGND VPWR VPWR clknet_5_10__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_28651_ _12822_ VGND VGND VPWR VPWR _04118_ sky130_fd_sc_hd__clkbuf_1
X_25863_ _11206_ _11207_ _11242_ VGND VGND VPWR VPWR _11243_ sky130_fd_sc_hd__and3_1
XFILLER_0_213_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27602_ _12235_ VGND VGND VPWR VPWR _03656_ sky130_fd_sc_hd__clkbuf_1
X_24814_ _10620_ VGND VGND VPWR VPWR _02483_ sky130_fd_sc_hd__clkbuf_1
X_28582_ _12785_ VGND VGND VPWR VPWR _04086_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_2_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25794_ net1675 _11181_ _11177_ _11187_ VGND VGND VPWR VPWR _02896_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_2_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27533_ _12128_ net2467 _12197_ VGND VGND VPWR VPWR _12199_ sky130_fd_sc_hd__mux2_1
X_24745_ _10388_ net3565 _10580_ VGND VGND VPWR VPWR _10582_ sky130_fd_sc_hd__mux2_1
X_21957_ _08692_ _09186_ _09188_ VGND VGND VPWR VPWR _09189_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_48_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_226_Right_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20908_ datamem.data_ram\[23\]\[22\] _07021_ _07182_ datamem.data_ram\[20\]\[22\]
+ _06681_ VGND VGND VPWR VPWR _08198_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_48_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_189_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27464_ _12161_ VGND VGND VPWR VPWR _03592_ sky130_fd_sc_hd__clkbuf_1
X_24676_ _10388_ datamem.data_ram\[4\]\[9\] _10543_ VGND VGND VPWR VPWR _10545_ sky130_fd_sc_hd__mux2_1
XFILLER_0_194_631 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21888_ _08842_ _09123_ VGND VGND VPWR VPWR _09124_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_104_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_104_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29203_ _13119_ VGND VGND VPWR VPWR _04373_ sky130_fd_sc_hd__clkbuf_1
X_26415_ _11545_ rvcpu.ALUResultE\[11\] VGND VGND VPWR VPWR _11554_ sky130_fd_sc_hd__and2_1
X_23627_ clknet_1_1__leaf__10172_ VGND VGND VPWR VPWR _10181_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_13_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20839_ _07840_ _08126_ _08128_ _07845_ VGND VGND VPWR VPWR _08129_ sky130_fd_sc_hd__a211o_1
X_27395_ _12117_ VGND VGND VPWR VPWR _03567_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_13_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_182_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29134_ _09255_ net3945 _13076_ VGND VGND VPWR VPWR _13083_ sky130_fd_sc_hd__mux2_1
X_26346_ _10058_ _11507_ _11508_ net1335 VGND VGND VPWR VPWR _03127_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22509_ _09469_ _09664_ VGND VGND VPWR VPWR _09665_ sky130_fd_sc_hd__or2_1
X_26277_ net1852 _11467_ VGND VGND VPWR VPWR _11471_ sky130_fd_sc_hd__and2_1
X_29065_ _13046_ VGND VGND VPWR VPWR _04308_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_712 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1114 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28016_ _12367_ net2899 net97 VGND VGND VPWR VPWR _12470_ sky130_fd_sc_hd__mux2_1
X_16030_ net1907 _13198_ _14349_ VGND VGND VPWR VPWR _14355_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25228_ _10853_ VGND VGND VPWR VPWR _02664_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_220_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25159_ _10811_ net3321 net58 VGND VGND VPWR VPWR _10813_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_204_5402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17981_ _05347_ _05176_ VGND VGND VPWR VPWR _05352_ sky130_fd_sc_hd__nor2_1
X_29967_ net337 _01702_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[15\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19720_ _06986_ _06988_ _07015_ VGND VGND VPWR VPWR _07016_ sky130_fd_sc_hd__and3_1
X_16932_ _04716_ VGND VGND VPWR VPWR _01574_ sky130_fd_sc_hd__clkbuf_1
X_28918_ _12964_ VGND VGND VPWR VPWR _04243_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_229_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29898_ net276 _01633_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[17\]\[29\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_196_5203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19651_ _06946_ VGND VGND VPWR VPWR _06947_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_217_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16863_ net2871 _14482_ _04670_ VGND VGND VPWR VPWR _04680_ sky130_fd_sc_hd__mux2_1
X_28849_ _12743_ net4190 net69 VGND VGND VPWR VPWR _12928_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_221_5793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18602_ _05676_ _05669_ _05758_ VGND VGND VPWR VPWR _05960_ sky130_fd_sc_hd__or3_2
X_15814_ _14238_ VGND VGND VPWR VPWR _02114_ sky130_fd_sc_hd__clkbuf_1
X_31860_ clknet_leaf_124_clk _03314_ VGND VGND VPWR VPWR datamem.data_ram\[62\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19582_ datamem.data_ram\[34\]\[8\] _06609_ _06780_ datamem.data_ram\[33\]\[8\] _06677_
+ VGND VGND VPWR VPWR _06878_ sky130_fd_sc_hd__o221a_1
X_16794_ _04643_ VGND VGND VPWR VPWR _01647_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_172_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_177_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30811_ clknet_leaf_135_clk _02546_ VGND VGND VPWR VPWR datamem.data_ram\[45\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_18533_ _05692_ _05893_ VGND VGND VPWR VPWR _05894_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23803__387 clknet_1_1__leaf__10206_ VGND VGND VPWR VPWR net513 sky130_fd_sc_hd__inv_2
X_15745_ _14201_ VGND VGND VPWR VPWR _02154_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_220_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31791_ clknet_leaf_234_clk _03245_ VGND VGND VPWR VPWR datamem.data_ram\[2\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_4210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30742_ clknet_leaf_148_clk _02477_ VGND VGND VPWR VPWR datamem.data_ram\[48\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_18464_ _05648_ _05642_ _05682_ VGND VGND VPWR VPWR _05827_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_155_4221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15676_ _14154_ net2602 _14152_ VGND VGND VPWR VPWR _14155_ sky130_fd_sc_hd__mux2_1
XANTENNA_260 _13209_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_271 _13235_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_200_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_282 _13260_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17415_ _04538_ _04900_ VGND VGND VPWR VPWR _04973_ sky130_fd_sc_hd__nand2_2
XANTENNA_293 _13350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_184_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14627_ net2064 _13204_ _13181_ VGND VGND VPWR VPWR _13205_ sky130_fd_sc_hd__mux2_1
X_18395_ _05756_ _05758_ _05668_ VGND VGND VPWR VPWR _05759_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30673_ clknet_leaf_179_clk _02408_ VGND VGND VPWR VPWR datamem.data_ram\[50\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_151_4118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_151_4129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32412_ clknet_leaf_231_clk _03834_ VGND VGND VPWR VPWR datamem.data_ram\[28\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17346_ _04936_ VGND VGND VPWR VPWR _01372_ sky130_fd_sc_hd__clkbuf_1
X_23617__235 clknet_1_0__leaf__10180_ VGND VGND VPWR VPWR net361 sky130_fd_sc_hd__inv_2
X_32343_ clknet_leaf_184_clk _03765_ VGND VGND VPWR VPWR datamem.data_ram\[30\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_17277_ _04899_ VGND VGND VPWR VPWR _01404_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload202 clknet_leaf_210_clk VGND VGND VPWR VPWR clkload202/Y sky130_fd_sc_hd__clkinvlp_2
X_23159__832 clknet_1_1__leaf__10109_ VGND VGND VPWR VPWR net958 sky130_fd_sc_hd__inv_2
Xclkload213 clknet_leaf_207_clk VGND VGND VPWR VPWR clkload213/Y sky130_fd_sc_hd__clkinv_1
XFILLER_0_144_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload224 clknet_leaf_163_clk VGND VGND VPWR VPWR clkload224/Y sky130_fd_sc_hd__clkinv_1
X_19016_ _05694_ _06348_ _06349_ _05703_ VGND VGND VPWR VPWR _06350_ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16228_ net2141 _14470_ _14464_ VGND VGND VPWR VPWR _14471_ sky130_fd_sc_hd__mux2_1
Xclkload235 clknet_leaf_115_clk VGND VGND VPWR VPWR clkload235/Y sky130_fd_sc_hd__clkinv_4
X_32274_ clknet_leaf_88_clk _03696_ VGND VGND VPWR VPWR datamem.data_ram\[33\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload246 clknet_leaf_149_clk VGND VGND VPWR VPWR clkload246/Y sky130_fd_sc_hd__inv_6
XFILLER_0_113_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload257 clknet_leaf_143_clk VGND VGND VPWR VPWR clkload257/Y sky130_fd_sc_hd__inv_8
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_228_5958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload268 clknet_leaf_131_clk VGND VGND VPWR VPWR clkload268/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_110_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_228_5969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31225_ clknet_leaf_39_clk _02928_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCD\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_185_4940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload279 clknet_1_1__leaf__10244_ VGND VGND VPWR VPWR clkload279/X sky130_fd_sc_hd__clkbuf_8
X_16159_ _13183_ VGND VGND VPWR VPWR _14424_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_110_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_110_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_4069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31156_ clknet_leaf_69_clk rvcpu.ALUResultE\[15\] VGND VGND VPWR VPWR rvcpu.dp.plem.ALUResultM\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_181_4837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_181_4848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2705 datamem.data_ram\[24\]\[25\] VGND VGND VPWR VPWR net3855 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30107_ net469 _01842_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[11\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_19918_ datamem.data_ram\[32\]\[17\] _07191_ _07209_ _07212_ VGND VGND VPWR VPWR
+ _07213_ sky130_fd_sc_hd__o211a_1
Xhold2716 rvcpu.dp.rf.reg_file_arr\[26\]\[18\] VGND VGND VPWR VPWR net3866 sky130_fd_sc_hd__dlygate4sd3_1
X_31087_ clknet_leaf_107_clk _02822_ VGND VGND VPWR VPWR datamem.data_ram\[21\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2727 datamem.data_ram\[30\]\[8\] VGND VGND VPWR VPWR net3877 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_71_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2738 datamem.data_ram\[45\]\[29\] VGND VGND VPWR VPWR net3888 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2749 rvcpu.dp.rf.reg_file_arr\[15\]\[1\] VGND VGND VPWR VPWR net3899 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19849_ datamem.data_ram\[50\]\[1\] _06932_ _06958_ datamem.data_ram\[49\]\[1\] _06742_
+ VGND VGND VPWR VPWR _07144_ sky130_fd_sc_hd__a221o_1
X_30038_ net400 _01773_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[13\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_24175__16 clknet_1_1__leaf__10265_ VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_108_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22860_ rvcpu.dp.rf.reg_file_arr\[4\]\[29\] rvcpu.dp.rf.reg_file_arr\[5\]\[29\] rvcpu.dp.rf.reg_file_arr\[6\]\[29\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[29\] _09416_ _09418_ VGND VGND VPWR VPWR _09997_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_84_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_140_3844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21811_ _08692_ _09048_ _09050_ VGND VGND VPWR VPWR _09051_ sky130_fd_sc_hd__a21o_1
XFILLER_0_218_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_3866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_179_4788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22791_ rvcpu.dp.rf.reg_file_arr\[4\]\[25\] rvcpu.dp.rf.reg_file_arr\[5\]\[25\] rvcpu.dp.rf.reg_file_arr\[6\]\[25\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[25\] _09464_ _09467_ VGND VGND VPWR VPWR _09932_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_179_4799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31989_ clknet_leaf_92_clk _03411_ VGND VGND VPWR VPWR datamem.data_ram\[37\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24530_ _10460_ VGND VGND VPWR VPWR _02359_ sky130_fd_sc_hd__clkbuf_1
X_21742_ _08977_ _08981_ _08985_ _08624_ VGND VGND VPWR VPWR _01046_ sky130_fd_sc_hd__o31a_1
XFILLER_0_210_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_878 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24461_ _10076_ _10406_ VGND VGND VPWR VPWR _10420_ sky130_fd_sc_hd__and2_1
X_21673_ _08798_ _08919_ VGND VGND VPWR VPWR _08920_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_43_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26200_ net116 VGND VGND VPWR VPWR _11438_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_43_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27180_ _11968_ _11996_ VGND VGND VPWR VPWR _11998_ sky130_fd_sc_hd__and2_1
X_20624_ _07839_ _07910_ _07914_ _07844_ VGND VGND VPWR VPWR _07915_ sky130_fd_sc_hd__a211o_1
X_24392_ _09260_ net4263 _10367_ VGND VGND VPWR VPWR _10375_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26131_ _11401_ VGND VGND VPWR VPWR _03018_ sky130_fd_sc_hd__clkbuf_1
X_20555_ _07842_ _07843_ _07845_ VGND VGND VPWR VPWR _07846_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_225_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26062_ _11064_ _11351_ VGND VGND VPWR VPWR _11360_ sky130_fd_sc_hd__and2_1
XFILLER_0_225_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20486_ datamem.data_ram\[59\]\[20\] _06634_ _07774_ _07777_ VGND VGND VPWR VPWR
+ _07778_ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25013_ _09275_ VGND VGND VPWR VPWR _10729_ sky130_fd_sc_hd__buf_2
X_22225_ _09390_ VGND VGND VPWR VPWR _09391_ sky130_fd_sc_hd__clkbuf_4
X_29821_ net199 _01556_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[1\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_22156_ _09288_ net2709 net62 VGND VGND VPWR VPWR _09348_ sky130_fd_sc_hd__mux2_1
X_21107_ datamem.data_ram\[16\]\[7\] datamem.data_ram\[17\]\[7\] _06651_ VGND VGND
+ VPWR VPWR _08396_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29752_ net1098 _01487_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[21\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_7_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26964_ _11864_ VGND VGND VPWR VPWR _11865_ sky130_fd_sc_hd__clkbuf_2
X_22087_ _09227_ net108 VGND VGND VPWR VPWR _09301_ sky130_fd_sc_hd__nor2_8
XTAP_TAPCELL_ROW_7_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28703_ _10979_ _12602_ _12795_ VGND VGND VPWR VPWR _12850_ sky130_fd_sc_hd__a21oi_4
X_25915_ net1783 _11263_ VGND VGND VPWR VPWR _11277_ sky130_fd_sc_hd__or2_1
X_21038_ _06605_ datamem.data_ram\[11\]\[31\] _06933_ datamem.data_ram\[10\]\[31\]
+ _07844_ VGND VGND VPWR VPWR _08327_ sky130_fd_sc_hd__o221a_1
XFILLER_0_22_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29683_ net1029 _01418_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[23\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_26895_ _07191_ _10918_ _10897_ VGND VGND VPWR VPWR _11820_ sky130_fd_sc_hd__or3_1
X_28634_ _12813_ VGND VGND VPWR VPWR _04110_ sky130_fd_sc_hd__clkbuf_1
X_25846_ rvcpu.dp.plfd.PCPlus4D\[25\] _11228_ _11142_ VGND VGND VPWR VPWR _11229_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_214_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_202_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23329__968 clknet_1_1__leaf__10135_ VGND VGND VPWR VPWR net1094 sky130_fd_sc_hd__inv_2
XFILLER_0_214_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28565_ _12776_ VGND VGND VPWR VPWR _04078_ sky130_fd_sc_hd__clkbuf_1
X_25777_ rvcpu.dp.pcreg.q\[11\] _11171_ VGND VGND VPWR VPWR _11174_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15530_ _13542_ _13604_ _13721_ VGND VGND VPWR VPWR _14056_ sky130_fd_sc_hd__and3_1
X_27516_ _12083_ net3452 net99 VGND VGND VPWR VPWR _12190_ sky130_fd_sc_hd__mux2_1
X_24728_ _10442_ net3188 _10571_ VGND VGND VPWR VPWR _10573_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28496_ _12727_ net1544 _12723_ _12732_ VGND VGND VPWR VPWR _04053_ sky130_fd_sc_hd__a31o_1
XFILLER_0_210_1304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_106_Left_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15461_ _13559_ _13351_ _13533_ VGND VGND VPWR VPWR _13991_ sky130_fd_sc_hd__a21oi_1
X_27447_ _12150_ VGND VGND VPWR VPWR _03586_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24659_ _10410_ _10532_ VGND VGND VPWR VPWR _10535_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_190_clk clknet_5_28__leaf_clk VGND VGND VPWR VPWR clknet_leaf_190_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_38_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_182_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17200_ _14187_ net4377 _04851_ VGND VGND VPWR VPWR _04859_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23108__786 clknet_1_0__leaf__10104_ VGND VGND VPWR VPWR net912 sky130_fd_sc_hd__inv_2
XFILLER_0_182_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18180_ rvcpu.dp.plde.RD1E\[26\] _05291_ _05544_ VGND VGND VPWR VPWR _05545_ sky130_fd_sc_hd__o21a_1
XFILLER_0_53_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15392_ _13919_ _13920_ _13921_ _13924_ VGND VGND VPWR VPWR _13925_ sky130_fd_sc_hd__a31o_1
X_27378_ _12108_ VGND VGND VPWR VPWR _03559_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_189_5040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17131_ _04822_ VGND VGND VPWR VPWR _01473_ sky130_fd_sc_hd__clkbuf_1
X_29117_ _09287_ net4011 _13067_ VGND VGND VPWR VPWR _13074_ sky130_fd_sc_hd__mux2_1
X_26329_ _11353_ net1731 _11496_ _11499_ VGND VGND VPWR VPWR _03119_ sky130_fd_sc_hd__a31o_1
XFILLER_0_135_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29048_ _13018_ net1703 _13030_ _13037_ VGND VGND VPWR VPWR _04300_ sky130_fd_sc_hd__a31o_1
X_17062_ net4226 _14476_ _04779_ VGND VGND VPWR VPWR _04786_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16013_ _14344_ VGND VGND VPWR VPWR _02021_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_115_Left_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31010_ clknet_leaf_157_clk _02745_ VGND VGND VPWR VPWR datamem.data_ram\[11\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_78_Right_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_223_5844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_223_5855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17964_ _05334_ _05310_ VGND VGND VPWR VPWR _05335_ sky130_fd_sc_hd__and2_1
XFILLER_0_224_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19703_ datamem.data_ram\[5\]\[0\] _06970_ _06967_ _06998_ VGND VGND VPWR VPWR _06999_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_109_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16915_ net2389 _14466_ _04706_ VGND VGND VPWR VPWR _04708_ sky130_fd_sc_hd__mux2_1
X_32961_ clknet_leaf_206_clk _04383_ VGND VGND VPWR VPWR datamem.data_ram\[63\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_17895_ _05244_ _05247_ _05251_ VGND VGND VPWR VPWR _05268_ sky130_fd_sc_hd__and3_4
XFILLER_0_139_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19634_ _06929_ VGND VGND VPWR VPWR _06930_ sky130_fd_sc_hd__clkbuf_8
X_31912_ _04423_ net120 VGND VGND VPWR VPWR datamem.rd_data_mem\[17\] sky130_fd_sc_hd__dlxtn_1
XFILLER_0_75_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16846_ _04671_ VGND VGND VPWR VPWR _01615_ sky130_fd_sc_hd__clkbuf_1
X_32892_ clknet_leaf_163_clk _04314_ VGND VGND VPWR VPWR datamem.data_ram\[10\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31843_ clknet_leaf_164_clk _03297_ VGND VGND VPWR VPWR datamem.data_ram\[8\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_19565_ _06752_ _06842_ _06847_ _06859_ _06860_ VGND VGND VPWR VPWR _06861_ sky130_fd_sc_hd__o311a_1
X_16777_ net3864 _14463_ _04634_ VGND VGND VPWR VPWR _04635_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_124_Left_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_87_Right_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18516_ _05837_ _05846_ _05859_ _05877_ VGND VGND VPWR VPWR rvcpu.ALUResultE\[2\]
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_125_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_220_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15728_ _14189_ net4013 _14173_ VGND VGND VPWR VPWR _14190_ sky130_fd_sc_hd__mux2_1
XFILLER_0_186_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19496_ datamem.data_ram\[26\]\[16\] _06611_ _06784_ datamem.data_ram\[31\]\[16\]
+ _06601_ VGND VGND VPWR VPWR _06792_ sky130_fd_sc_hd__o221a_1
XFILLER_0_73_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31774_ clknet_leaf_208_clk _03228_ VGND VGND VPWR VPWR datamem.data_ram\[1\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_174_4663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18447_ _05575_ _05389_ VGND VGND VPWR VPWR _05810_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_506 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30725_ clknet_leaf_217_clk _02460_ VGND VGND VPWR VPWR datamem.data_ram\[48\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_174_4674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15659_ _13200_ VGND VGND VPWR VPWR _14143_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_34_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_181_clk clknet_5_19__leaf_clk VGND VGND VPWR VPWR clknet_leaf_181_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_200_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18378_ _05741_ _05280_ VGND VGND VPWR VPWR _05742_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30656_ clknet_leaf_219_clk _02391_ VGND VGND VPWR VPWR datamem.data_ram\[50\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17329_ net4213 _13253_ _04924_ VGND VGND VPWR VPWR _04928_ sky130_fd_sc_hd__mux2_1
X_30587_ clknet_leaf_177_clk _02322_ VGND VGND VPWR VPWR datamem.data_ram\[53\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20340_ datamem.data_ram\[58\]\[4\] _06989_ _06990_ datamem.data_ram\[56\]\[4\] VGND
+ VGND VPWR VPWR _07632_ sky130_fd_sc_hd__a22o_1
X_32326_ clknet_leaf_82_clk _03748_ VGND VGND VPWR VPWR datamem.data_ram\[31\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_133_3681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_3692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_133_Left_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_96_Right_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20271_ datamem.data_ram\[39\]\[19\] _06760_ _06699_ datamem.data_ram\[33\]\[19\]
+ VGND VGND VPWR VPWR _07564_ sky130_fd_sc_hd__o22a_1
XFILLER_0_3_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32257_ clknet_leaf_242_clk _03679_ VGND VGND VPWR VPWR datamem.data_ram\[34\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22010_ rvcpu.dp.plem.WriteDataM\[18\] _09221_ VGND VGND VPWR VPWR _09238_ sky130_fd_sc_hd__and2_1
X_31208_ clknet_leaf_34_clk _02911_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCPlus4D\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_228_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3203 datamem.data_ram\[58\]\[17\] VGND VGND VPWR VPWR net4353 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold3214 datamem.data_ram\[62\]\[23\] VGND VGND VPWR VPWR net4364 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32188_ clknet_leaf_256_clk _03610_ VGND VGND VPWR VPWR datamem.data_ram\[37\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3225 datamem.data_ram\[25\]\[18\] VGND VGND VPWR VPWR net4375 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3236 datamem.data_ram\[55\]\[23\] VGND VGND VPWR VPWR net4386 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3247 datamem.data_ram\[25\]\[22\] VGND VGND VPWR VPWR net4397 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2502 datamem.data_ram\[27\]\[25\] VGND VGND VPWR VPWR net3652 sky130_fd_sc_hd__dlygate4sd3_1
X_31139_ clknet_leaf_187_clk _02874_ VGND VGND VPWR VPWR datamem.data_ram\[4\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2513 datamem.data_ram\[42\]\[20\] VGND VGND VPWR VPWR net3663 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3258 rvcpu.dp.rf.reg_file_arr\[23\]\[24\] VGND VGND VPWR VPWR net4408 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2524 rvcpu.dp.rf.reg_file_arr\[18\]\[17\] VGND VGND VPWR VPWR net3674 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3269 datamem.data_ram\[52\]\[14\] VGND VGND VPWR VPWR net4419 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2535 rvcpu.dp.rf.reg_file_arr\[14\]\[26\] VGND VGND VPWR VPWR net3685 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2546 rvcpu.dp.rf.reg_file_arr\[27\]\[31\] VGND VGND VPWR VPWR net3696 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1801 datamem.data_ram\[34\]\[10\] VGND VGND VPWR VPWR net2951 sky130_fd_sc_hd__dlygate4sd3_1
X_23961_ _10234_ VGND VGND VPWR VPWR _02016_ sky130_fd_sc_hd__clkbuf_1
Xhold2557 rvcpu.dp.rf.reg_file_arr\[15\]\[26\] VGND VGND VPWR VPWR net3707 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1812 datamem.data_ram\[2\]\[8\] VGND VGND VPWR VPWR net2962 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1823 datamem.data_ram\[45\]\[20\] VGND VGND VPWR VPWR net2973 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2568 datamem.data_ram\[25\]\[13\] VGND VGND VPWR VPWR net3718 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1834 datamem.data_ram\[39\]\[26\] VGND VGND VPWR VPWR net2984 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2579 datamem.data_ram\[23\]\[31\] VGND VGND VPWR VPWR net3729 sky130_fd_sc_hd__dlygate4sd3_1
X_25700_ _11121_ net1846 _11111_ _11122_ VGND VGND VPWR VPWR _02867_ sky130_fd_sc_hd__a31o_1
XFILLER_0_192_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1845 datamem.data_ram\[16\]\[10\] VGND VGND VPWR VPWR net2995 sky130_fd_sc_hd__dlygate4sd3_1
X_22912_ _10045_ VGND VGND VPWR VPWR _10046_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_32_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26680_ _11692_ VGND VGND VPWR VPWR _11693_ sky130_fd_sc_hd__clkbuf_2
Xhold1856 datamem.data_ram\[20\]\[16\] VGND VGND VPWR VPWR net3006 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1867 rvcpu.dp.rf.reg_file_arr\[1\]\[13\] VGND VGND VPWR VPWR net3017 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1878 rvcpu.dp.rf.reg_file_arr\[22\]\[13\] VGND VGND VPWR VPWR net3028 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_142_Left_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1889 datamem.data_ram\[19\]\[18\] VGND VGND VPWR VPWR net3039 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25631_ _10060_ VGND VGND VPWR VPWR _11083_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_211_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22843_ _09636_ _09980_ VGND VGND VPWR VPWR _09981_ sky130_fd_sc_hd__or2_1
Xclkbuf_1_1__f__10180_ clknet_0__10180_ VGND VGND VPWR VPWR clknet_1_1__leaf__10180_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_190_1053 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28350_ _12649_ VGND VGND VPWR VPWR _03990_ sky130_fd_sc_hd__clkbuf_1
X_25562_ _10946_ _11039_ VGND VGND VPWR VPWR _11040_ sky130_fd_sc_hd__or2_1
X_22774_ _09481_ _09915_ VGND VGND VPWR VPWR _09916_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_101_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27301_ _07203_ _09227_ _11839_ VGND VGND VPWR VPWR _12064_ sky130_fd_sc_hd__or3_1
XFILLER_0_78_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24513_ _09251_ VGND VGND VPWR VPWR _10450_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_148_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21725_ rvcpu.dp.rf.reg_file_arr\[16\]\[18\] rvcpu.dp.rf.reg_file_arr\[17\]\[18\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[18\] rvcpu.dp.rf.reg_file_arr\[19\]\[18\] _08703_
+ _08721_ VGND VGND VPWR VPWR _08969_ sky130_fd_sc_hd__mux4_1
X_24073__599 clknet_1_1__leaf__10248_ VGND VGND VPWR VPWR net725 sky130_fd_sc_hd__inv_2
X_28281_ _08133_ _09228_ VGND VGND VPWR VPWR _12612_ sky130_fd_sc_hd__nor2_8
X_25493_ _11001_ VGND VGND VPWR VPWR _02781_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_172_clk clknet_5_24__leaf_clk VGND VGND VPWR VPWR clknet_leaf_172_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_17_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27232_ _11980_ _12019_ VGND VGND VPWR VPWR _12028_ sky130_fd_sc_hd__and2_1
XFILLER_0_191_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24444_ _10408_ _10406_ VGND VGND VPWR VPWR _10409_ sky130_fd_sc_hd__and2_1
X_21656_ rvcpu.dp.rf.reg_file_arr\[16\]\[14\] rvcpu.dp.rf.reg_file_arr\[17\]\[14\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[14\] rvcpu.dp.rf.reg_file_arr\[19\]\[14\] _08524_
+ _08527_ VGND VGND VPWR VPWR _08904_ sky130_fd_sc_hd__mux4_1
XFILLER_0_53_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20607_ _07895_ _07897_ _07872_ VGND VGND VPWR VPWR _07898_ sky130_fd_sc_hd__a21o_1
X_27163_ _11974_ net1590 _11983_ _11987_ VGND VGND VPWR VPWR _03465_ sky130_fd_sc_hd__a31o_1
XFILLER_0_117_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24375_ _10365_ VGND VGND VPWR VPWR _02299_ sky130_fd_sc_hd__clkbuf_1
X_21587_ _08566_ VGND VGND VPWR VPWR _08839_ sky130_fd_sc_hd__buf_6
XPHY_EDGE_ROW_151_Left_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26114_ _11392_ VGND VGND VPWR VPWR _03010_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_163_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20538_ _07828_ VGND VGND VPWR VPWR _07829_ sky130_fd_sc_hd__buf_6
X_27094_ _11938_ net1797 _11940_ _11943_ VGND VGND VPWR VPWR _03440_ sky130_fd_sc_hd__a31o_1
XFILLER_0_144_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26045_ _11349_ VGND VGND VPWR VPWR _11350_ sky130_fd_sc_hd__clkbuf_2
X_20469_ datamem.data_ram\[46\]\[20\] _06744_ _06725_ datamem.data_ram\[47\]\[20\]
+ _07760_ VGND VGND VPWR VPWR _07761_ sky130_fd_sc_hd__o221a_1
XFILLER_0_104_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22208_ _09285_ net3637 _09371_ VGND VGND VPWR VPWR _09377_ sky130_fd_sc_hd__mux2_1
X_23188_ _08144_ net104 VGND VGND VPWR VPWR _10114_ sky130_fd_sc_hd__nor2_8
Xclkbuf_5_8__f_clk clknet_2_1_0_clk VGND VGND VPWR VPWR clknet_5_8__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_30_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29804_ clknet_leaf_202_clk _01539_ VGND VGND VPWR VPWR datamem.data_ram\[59\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_973 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22139_ _09256_ net3924 _09332_ VGND VGND VPWR VPWR _09339_ sky130_fd_sc_hd__mux2_1
XFILLER_0_207_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27996_ _09284_ VGND VGND VPWR VPWR _12458_ sky130_fd_sc_hd__buf_2
XFILLER_0_203_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_218_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29735_ net1081 _01470_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[21\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_14961_ _13397_ _13307_ VGND VGND VPWR VPWR _13510_ sky130_fd_sc_hd__nand2_4
X_26947_ _11849_ net1422 _11853_ _11855_ VGND VGND VPWR VPWR _03381_ sky130_fd_sc_hd__a31o_1
Xhold8 rvcpu.dp.plem.PCPlus4M\[24\] VGND VGND VPWR VPWR net1158 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_160_Left_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16700_ _14164_ net2919 _04587_ VGND VGND VPWR VPWR _04594_ sky130_fd_sc_hd__mux2_1
X_29666_ net1012 _01401_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[24\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_17680_ _05113_ VGND VGND VPWR VPWR _01199_ sky130_fd_sc_hd__clkbuf_1
X_26878_ _11676_ _11810_ VGND VGND VPWR VPWR _11811_ sky130_fd_sc_hd__and2_1
X_14892_ _13337_ _13435_ VGND VGND VPWR VPWR _13443_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_226_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16631_ _04557_ VGND VGND VPWR VPWR _01724_ sky130_fd_sc_hd__clkbuf_1
X_28617_ _12804_ VGND VGND VPWR VPWR _04102_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25829_ _11213_ _11214_ VGND VGND VPWR VPWR _11215_ sky130_fd_sc_hd__nor2_1
X_29597_ net951 _01332_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[25\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23262__908 clknet_1_0__leaf__10128_ VGND VGND VPWR VPWR net1034 sky130_fd_sc_hd__inv_2
XFILLER_0_69_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19350_ _06645_ VGND VGND VPWR VPWR _06646_ sky130_fd_sc_hd__buf_8
X_28548_ _12767_ VGND VGND VPWR VPWR _04070_ sky130_fd_sc_hd__clkbuf_1
X_16562_ _04520_ VGND VGND VPWR VPWR _01764_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18301_ _05665_ VGND VGND VPWR VPWR _05666_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_210_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15513_ _13326_ _13585_ _14037_ _14039_ VGND VGND VPWR VPWR _14040_ sky130_fd_sc_hd__a31o_1
XFILLER_0_183_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19281_ _06567_ _06578_ VGND VGND VPWR VPWR _06579_ sky130_fd_sc_hd__and2_1
X_28479_ _07808_ _10042_ _10044_ VGND VGND VPWR VPWR _12722_ sky130_fd_sc_hd__or3_1
Xclkbuf_leaf_163_clk clknet_5_25__leaf_clk VGND VGND VPWR VPWR clknet_leaf_163_clk
+ sky130_fd_sc_hd__clkbuf_8
X_16493_ net2760 _14453_ _04478_ VGND VGND VPWR VPWR _04484_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_216_5670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_216_5681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18232_ _05596_ _05343_ VGND VGND VPWR VPWR _05597_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30510_ clknet_leaf_208_clk _02245_ VGND VGND VPWR VPWR datamem.data_ram\[56\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_15444_ _13472_ _13565_ _13482_ VGND VGND VPWR VPWR _13975_ sky130_fd_sc_hd__a21o_1
X_31490_ clknet_leaf_47_clk rvcpu.dp.lAuiPCE\[16\] VGND VGND VPWR VPWR rvcpu.dp.plem.lAuiPCM\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_212_5578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18163_ rvcpu.dp.plde.ImmExtE\[25\] rvcpu.dp.SrcBFW_Mux.y\[25\] _05279_ VGND VGND
+ VPWR VPWR _05528_ sky130_fd_sc_hd__mux2_1
X_30441_ net779 _02176_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[29\]\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_212_5589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15375_ _13304_ _13425_ VGND VGND VPWR VPWR _13909_ sky130_fd_sc_hd__nor2_1
XFILLER_0_182_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17114_ _04813_ VGND VGND VPWR VPWR _01481_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18094_ rvcpu.dp.plem.ALUResultM\[22\] _05339_ _05340_ _13209_ VGND VGND VPWR VPWR
+ _05462_ sky130_fd_sc_hd__o22a_1
XFILLER_0_20_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30372_ net718 _02107_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[3\]\[23\] sky130_fd_sc_hd__dfxtp_1
Xmax_cap105 _05307_ VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_111_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold408 datamem.data_ram\[21\]\[4\] VGND VGND VPWR VPWR net1558 sky130_fd_sc_hd__dlygate4sd3_1
X_32111_ clknet_leaf_119_clk _03533_ VGND VGND VPWR VPWR datamem.data_ram\[58\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xmax_cap116 _11377_ VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__buf_1
Xhold419 datamem.data_ram\[5\]\[2\] VGND VGND VPWR VPWR net1569 sky130_fd_sc_hd__dlygate4sd3_1
X_17045_ net2827 _14459_ _04768_ VGND VGND VPWR VPWR _04777_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_225_5906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_180_1266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_4006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32042_ clknet_leaf_132_clk _03464_ VGND VGND VPWR VPWR datamem.data_ram\[49\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18996_ _06004_ _06330_ _06097_ VGND VGND VPWR VPWR _06331_ sky130_fd_sc_hd__a21bo_1
X_17947_ rvcpu.dp.plem.ALUResultM\[13\] _05268_ VGND VGND VPWR VPWR _05319_ sky130_fd_sc_hd__and2_1
Xhold1108 rvcpu.dp.rf.reg_file_arr\[8\]\[29\] VGND VGND VPWR VPWR net2258 sky130_fd_sc_hd__dlygate4sd3_1
X_23809__393 clknet_1_1__leaf__10206_ VGND VGND VPWR VPWR net519 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_163_4397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1119 datamem.data_ram\[31\]\[22\] VGND VGND VPWR VPWR net2269 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32944_ clknet_leaf_146_clk _04366_ VGND VGND VPWR VPWR datamem.data_ram\[6\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_105_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17878_ _05248_ rvcpu.dp.plem.RdM\[3\] _05249_ _05250_ rvcpu.dp.plem.RegWriteM VGND
+ VGND VPWR VPWR _05251_ sky130_fd_sc_hd__o221a_1
XFILLER_0_174_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19617_ _06799_ _06910_ _06912_ VGND VGND VPWR VPWR _06913_ sky130_fd_sc_hd__mux2_1
X_16829_ _04662_ VGND VGND VPWR VPWR _01623_ sky130_fd_sc_hd__clkbuf_1
X_32875_ clknet_leaf_56_clk _04297_ VGND VGND VPWR VPWR datamem.data_ram\[10\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_176_4714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_176_4725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_220_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31826_ clknet_leaf_105_clk _03280_ VGND VGND VPWR VPWR datamem.data_ram\[16\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_19548_ datamem.data_ram\[22\]\[24\] _06718_ _06696_ datamem.data_ram\[16\]\[24\]
+ VGND VGND VPWR VPWR _06844_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_66_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_193_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31757_ clknet_leaf_72_clk _03211_ VGND VGND VPWR VPWR datamem.data_ram\[45\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_19479_ datamem.data_ram\[21\]\[16\] _06665_ _06621_ datamem.data_ram\[20\]\[16\]
+ VGND VGND VPWR VPWR _06775_ sky130_fd_sc_hd__o22a_1
XFILLER_0_152_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_154_clk clknet_5_28__leaf_clk VGND VGND VPWR VPWR clknet_leaf_154_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_146_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21510_ rvcpu.dp.rf.reg_file_arr\[24\]\[7\] rvcpu.dp.rf.reg_file_arr\[25\]\[7\] rvcpu.dp.rf.reg_file_arr\[26\]\[7\]
+ rvcpu.dp.rf.reg_file_arr\[27\]\[7\] _08517_ _08519_ VGND VGND VPWR VPWR _08765_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_145_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30708_ clknet_leaf_199_clk _02443_ VGND VGND VPWR VPWR datamem.data_ram\[49\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22490_ _09461_ _09644_ _09646_ _09489_ VGND VGND VPWR VPWR _09647_ sky130_fd_sc_hd__o211a_1
X_31688_ clknet_leaf_33_clk _03146_ VGND VGND VPWR VPWR rvcpu.dp.pcreg.q\[6\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_79_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_3732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_695 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_3743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21441_ _08699_ VGND VGND VPWR VPWR _08700_ sky130_fd_sc_hd__clkbuf_4
X_30639_ clknet_leaf_192_clk _02374_ VGND VGND VPWR VPWR datamem.data_ram\[51\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_3629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21372_ rvcpu.dp.rf.reg_file_arr\[20\]\[1\] rvcpu.dp.rf.reg_file_arr\[21\]\[1\] rvcpu.dp.rf.reg_file_arr\[22\]\[1\]
+ rvcpu.dp.rf.reg_file_arr\[23\]\[1\] _08631_ _08632_ VGND VGND VPWR VPWR _08633_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_160_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20323_ datamem.data_ram\[28\]\[4\] _07123_ _07611_ _07614_ VGND VGND VPWR VPWR _07615_
+ sky130_fd_sc_hd__a211o_1
X_32309_ clknet_leaf_263_clk _03731_ VGND VGND VPWR VPWR datamem.data_ram\[32\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_96_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24091_ _10257_ VGND VGND VPWR VPWR _02123_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_9_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold920 rvcpu.dp.rf.reg_file_arr\[7\]\[3\] VGND VGND VPWR VPWR net2070 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold931 rvcpu.dp.rf.reg_file_arr\[1\]\[22\] VGND VGND VPWR VPWR net2081 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold942 rvcpu.dp.rf.reg_file_arr\[18\]\[7\] VGND VGND VPWR VPWR net2092 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20254_ datamem.data_ram\[42\]\[3\] _06931_ _06924_ datamem.data_ram\[47\]\[3\] VGND
+ VGND VPWR VPWR _07547_ sky130_fd_sc_hd__a22o_1
Xhold953 rvcpu.dp.rf.reg_file_arr\[4\]\[10\] VGND VGND VPWR VPWR net2103 sky130_fd_sc_hd__dlygate4sd3_1
Xhold964 datamem.data_ram\[49\]\[23\] VGND VGND VPWR VPWR net2114 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold3000 rvcpu.dp.rf.reg_file_arr\[28\]\[11\] VGND VGND VPWR VPWR net4150 sky130_fd_sc_hd__dlygate4sd3_1
Xhold975 datamem.data_ram\[38\]\[30\] VGND VGND VPWR VPWR net2125 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3011 rvcpu.dp.rf.reg_file_arr\[29\]\[30\] VGND VGND VPWR VPWR net4161 sky130_fd_sc_hd__dlygate4sd3_1
Xhold986 rvcpu.dp.rf.reg_file_arr\[5\]\[8\] VGND VGND VPWR VPWR net2136 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3022 datamem.data_ram\[9\]\[18\] VGND VGND VPWR VPWR net4172 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_34_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27850_ _10668_ _12335_ _12356_ VGND VGND VPWR VPWR _12373_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_34_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold997 datamem.data_ram\[62\]\[29\] VGND VGND VPWR VPWR net2147 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3033 datamem.data_ram\[15\]\[14\] VGND VGND VPWR VPWR net4183 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20185_ datamem.data_ram\[6\]\[11\] _07085_ _07243_ datamem.data_ram\[1\]\[11\] VGND
+ VGND VPWR VPWR _07478_ sky130_fd_sc_hd__o22a_1
Xhold3044 datamem.data_ram\[3\]\[28\] VGND VGND VPWR VPWR net4194 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3055 rvcpu.dp.rf.reg_file_arr\[2\]\[6\] VGND VGND VPWR VPWR net4205 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2310 rvcpu.dp.rf.reg_file_arr\[4\]\[31\] VGND VGND VPWR VPWR net3460 sky130_fd_sc_hd__dlygate4sd3_1
X_26801_ _11753_ net1426 _11761_ _11764_ VGND VGND VPWR VPWR _03326_ sky130_fd_sc_hd__a31o_1
Xhold2321 rvcpu.dp.rf.reg_file_arr\[12\]\[20\] VGND VGND VPWR VPWR net3471 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3066 datamem.data_ram\[30\]\[27\] VGND VGND VPWR VPWR net4216 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3077 datamem.data_ram\[53\]\[26\] VGND VGND VPWR VPWR net4227 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2332 datamem.data_ram\[23\]\[15\] VGND VGND VPWR VPWR net3482 sky130_fd_sc_hd__dlygate4sd3_1
X_27781_ _12331_ VGND VGND VPWR VPWR _03739_ sky130_fd_sc_hd__clkbuf_1
Xhold3088 rvcpu.dp.rf.reg_file_arr\[16\]\[31\] VGND VGND VPWR VPWR net4238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2343 datamem.data_ram\[20\]\[15\] VGND VGND VPWR VPWR net3493 sky130_fd_sc_hd__dlygate4sd3_1
X_24993_ _10717_ VGND VGND VPWR VPWR _02565_ sky130_fd_sc_hd__clkbuf_1
Xhold2354 datamem.data_ram\[58\]\[22\] VGND VGND VPWR VPWR net3504 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3099 rvcpu.dp.rf.reg_file_arr\[15\]\[18\] VGND VGND VPWR VPWR net4249 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1620 datamem.data_ram\[12\]\[18\] VGND VGND VPWR VPWR net2770 sky130_fd_sc_hd__dlygate4sd3_1
X_29520_ net882 _01255_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[28\]\[27\] sky130_fd_sc_hd__dfxtp_1
Xhold2365 rvcpu.dp.rf.reg_file_arr\[28\]\[10\] VGND VGND VPWR VPWR net3515 sky130_fd_sc_hd__dlygate4sd3_1
X_26732_ _10766_ net3327 _11714_ VGND VGND VPWR VPWR _11722_ sky130_fd_sc_hd__mux2_1
Xhold2376 datamem.data_ram\[31\]\[25\] VGND VGND VPWR VPWR net3526 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1631 datamem.data_ram\[43\]\[8\] VGND VGND VPWR VPWR net2781 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2387 datamem.data_ram\[48\]\[19\] VGND VGND VPWR VPWR net3537 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1642 datamem.data_ram\[31\]\[30\] VGND VGND VPWR VPWR net2792 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_192_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1653 datamem.data_ram\[39\]\[25\] VGND VGND VPWR VPWR net2803 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2398 datamem.data_ram\[17\]\[26\] VGND VGND VPWR VPWR net3548 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1664 rvcpu.dp.rf.reg_file_arr\[20\]\[6\] VGND VGND VPWR VPWR net2814 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1675 datamem.data_ram\[18\]\[23\] VGND VGND VPWR VPWR net2825 sky130_fd_sc_hd__dlygate4sd3_1
X_29451_ net813 _01186_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[30\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_26663_ _11681_ _11677_ VGND VGND VPWR VPWR _11682_ sky130_fd_sc_hd__and2_1
XFILLER_0_169_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1686 rvcpu.dp.rf.reg_file_arr\[5\]\[27\] VGND VGND VPWR VPWR net2836 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1697 rvcpu.dp.rf.reg_file_arr\[31\]\[15\] VGND VGND VPWR VPWR net2847 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28402_ _12677_ VGND VGND VPWR VPWR _04014_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_212_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25614_ _11071_ VGND VGND VPWR VPWR _02832_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0__10263_ _10263_ VGND VGND VPWR VPWR clknet_0__10263_ sky130_fd_sc_hd__clkbuf_16
X_29382_ clknet_leaf_176_clk _01117_ VGND VGND VPWR VPWR datamem.data_ram\[60\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22826_ rvcpu.dp.rf.reg_file_arr\[8\]\[27\] rvcpu.dp.rf.reg_file_arr\[10\]\[27\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[27\] rvcpu.dp.rf.reg_file_arr\[11\]\[27\] _09483_
+ _09656_ VGND VGND VPWR VPWR _09965_ sky130_fd_sc_hd__mux4_1
X_26594_ _11086_ _11640_ VGND VGND VPWR VPWR _11644_ sky130_fd_sc_hd__and2_1
XFILLER_0_196_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28333_ _12640_ VGND VGND VPWR VPWR _03982_ sky130_fd_sc_hd__clkbuf_1
X_25545_ _10751_ net2315 _11030_ VGND VGND VPWR VPWR _11031_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__10194_ _10194_ VGND VGND VPWR VPWR clknet_0__10194_ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_145_clk clknet_5_29__leaf_clk VGND VGND VPWR VPWR clknet_leaf_145_clk
+ sky130_fd_sc_hd__clkbuf_8
X_22757_ _09627_ _09897_ _09899_ _09795_ VGND VGND VPWR VPWR _09900_ sky130_fd_sc_hd__a211o_1
XFILLER_0_149_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21708_ rvcpu.dp.rf.reg_file_arr\[20\]\[17\] rvcpu.dp.rf.reg_file_arr\[21\]\[17\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[17\] rvcpu.dp.rf.reg_file_arr\[23\]\[17\] _08778_
+ _08825_ VGND VGND VPWR VPWR _08953_ sky130_fd_sc_hd__mux4_1
X_28264_ _12601_ _12602_ _12573_ VGND VGND VPWR VPWR _12603_ sky130_fd_sc_hd__a21oi_4
X_25476_ _10991_ net1442 _10984_ _10994_ VGND VGND VPWR VPWR _02771_ sky130_fd_sc_hd__a31o_1
X_22688_ rvcpu.dp.rf.reg_file_arr\[20\]\[20\] rvcpu.dp.rf.reg_file_arr\[21\]\[20\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[20\] rvcpu.dp.rf.reg_file_arr\[23\]\[20\] _09517_
+ _09577_ VGND VGND VPWR VPWR _09834_ sky130_fd_sc_hd__mux4_2
XFILLER_0_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_229_6006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27215_ _12017_ VGND VGND VPWR VPWR _12018_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_229_6017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21639_ _08742_ _08887_ VGND VGND VPWR VPWR _08888_ sky130_fd_sc_hd__or2_1
XFILLER_0_81_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24427_ _09284_ VGND VGND VPWR VPWR _10396_ sky130_fd_sc_hd__buf_2
X_28195_ _12565_ VGND VGND VPWR VPWR _03919_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_229_Left_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_212_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15160_ _13475_ _13290_ VGND VGND VPWR VPWR _13704_ sky130_fd_sc_hd__nor2_1
X_27146_ _10069_ VGND VGND VPWR VPWR _11976_ sky130_fd_sc_hd__buf_2
XFILLER_0_180_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24358_ _10356_ VGND VGND VPWR VPWR _02291_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15091_ _13627_ _13633_ _13636_ VGND VGND VPWR VPWR _13637_ sky130_fd_sc_hd__or3b_1
XFILLER_0_120_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27077_ _11919_ net1397 _11923_ _11931_ VGND VGND VPWR VPWR _03435_ sky130_fd_sc_hd__a31o_1
XFILLER_0_127_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24289_ _09273_ net4202 _10316_ VGND VGND VPWR VPWR _10318_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26028_ _11078_ _11340_ VGND VGND VPWR VPWR _11341_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24123__629 clknet_1_0__leaf__10260_ VGND VGND VPWR VPWR net755 sky130_fd_sc_hd__inv_2
X_18850_ _05454_ _05498_ _05504_ _05513_ _05519_ VGND VGND VPWR VPWR _06194_ sky130_fd_sc_hd__a41o_1
XFILLER_0_197_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17801_ _05154_ _05161_ VGND VGND VPWR VPWR _05194_ sky130_fd_sc_hd__nand2_2
X_18781_ _05239_ _06124_ _06126_ _06129_ VGND VGND VPWR VPWR _06130_ sky130_fd_sc_hd__a211o_1
X_27979_ _12446_ VGND VGND VPWR VPWR _03822_ sky130_fd_sc_hd__clkbuf_1
X_15993_ _14334_ VGND VGND VPWR VPWR _02031_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_206_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29718_ net1064 _01453_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[22\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_17732_ _05141_ VGND VGND VPWR VPWR _01175_ sky130_fd_sc_hd__clkbuf_1
X_14944_ _13415_ _13492_ VGND VGND VPWR VPWR _13493_ sky130_fd_sc_hd__nor2_2
XFILLER_0_101_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30990_ clknet_leaf_102_clk _02725_ VGND VGND VPWR VPWR datamem.data_ram\[13\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_26506__58 clknet_1_1__leaf__11602_ VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__inv_2
XFILLER_0_175_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29649_ net995 _01384_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[24\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_17663_ net2314 _13243_ _05104_ VGND VGND VPWR VPWR _05105_ sky130_fd_sc_hd__mux2_1
X_14875_ _13424_ _13426_ VGND VGND VPWR VPWR _13427_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_218_5721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19402_ _06697_ VGND VGND VPWR VPWR _06698_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_218_5732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_203_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16614_ _04548_ VGND VGND VPWR VPWR _01732_ sky130_fd_sc_hd__clkbuf_1
X_32660_ clknet_leaf_79_clk _04082_ VGND VGND VPWR VPWR datamem.data_ram\[19\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_17594_ _05045_ VGND VGND VPWR VPWR _05068_ sky130_fd_sc_hd__buf_4
XFILLER_0_159_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31611_ clknet_leaf_18_clk net1177 VGND VGND VPWR VPWR rvcpu.dp.plmw.PCPlus4W\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_19333_ _06628_ VGND VGND VPWR VPWR _06629_ sky130_fd_sc_hd__buf_8
XFILLER_0_175_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16545_ _04511_ VGND VGND VPWR VPWR _01772_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_214_5629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_171_4600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_136_clk clknet_5_30__leaf_clk VGND VGND VPWR VPWR clknet_leaf_136_clk
+ sky130_fd_sc_hd__clkbuf_8
X_32591_ clknet_leaf_73_clk _04013_ VGND VGND VPWR VPWR datamem.data_ram\[21\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_171_4611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19264_ _06564_ _05559_ _05655_ VGND VGND VPWR VPWR _06565_ sky130_fd_sc_hd__o21a_1
X_31542_ clknet_leaf_16_clk net1283 VGND VGND VPWR VPWR rvcpu.dp.plem.RdM\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22984__691 clknet_1_1__leaf__10083_ VGND VGND VPWR VPWR net817 sky130_fd_sc_hd__inv_2
X_16476_ net3108 _14436_ _04467_ VGND VGND VPWR VPWR _04475_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18215_ rvcpu.dp.plde.RD1E\[1\] _05266_ _05270_ _13274_ _05387_ VGND VGND VPWR VPWR
+ _05580_ sky130_fd_sc_hd__a221o_1
XFILLER_0_128_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15427_ _13542_ _13473_ _13853_ _13957_ _13475_ VGND VGND VPWR VPWR _13958_ sky130_fd_sc_hd__o311a_1
XFILLER_0_115_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19195_ _06505_ rvcpu.dp.plde.ImmExtE\[22\] _06493_ VGND VGND VPWR VPWR _06506_ sky130_fd_sc_hd__mux2_1
X_31473_ clknet_leaf_5_clk rvcpu.dp.SrcBFW_Mux.y\[31\] VGND VGND VPWR VPWR rvcpu.dp.plem.WriteDataM\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_182_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_182_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_208_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18146_ _05506_ _05509_ VGND VGND VPWR VPWR _05511_ sky130_fd_sc_hd__nor2_1
X_30424_ net762 _02159_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[29\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15358_ _13332_ _13634_ VGND VGND VPWR VPWR _13893_ sky130_fd_sc_hd__nor2_2
XFILLER_0_54_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_4540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold205 datamem.data_ram\[4\]\[6\] VGND VGND VPWR VPWR net1355 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_169_4551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18077_ _05442_ _05443_ _05444_ VGND VGND VPWR VPWR _05445_ sky130_fd_sc_hd__o21bai_1
X_30355_ net701 _02090_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[3\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_223_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15289_ _13682_ _13780_ _13805_ VGND VGND VPWR VPWR _13827_ sky130_fd_sc_hd__o21ai_1
Xhold216 datamem.data_ram\[47\]\[5\] VGND VGND VPWR VPWR net1366 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_169_4562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold227 rvcpu.dp.plfd.PCD\[1\] VGND VGND VPWR VPWR net1377 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold238 datamem.data_ram\[12\]\[2\] VGND VGND VPWR VPWR net1388 sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 datamem.data_ram\[29\]\[7\] VGND VGND VPWR VPWR net1399 sky130_fd_sc_hd__dlygate4sd3_1
X_17028_ _04756_ VGND VGND VPWR VPWR _04768_ sky130_fd_sc_hd__buf_4
X_30286_ net632 _02021_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[5\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_165_4448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_165_4459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32025_ clknet_leaf_127_clk _03447_ VGND VGND VPWR VPWR datamem.data_ram\[26\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24098__606 clknet_1_1__leaf__10258_ VGND VGND VPWR VPWR net732 sky130_fd_sc_hd__inv_2
XFILLER_0_226_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18979_ _05694_ _05819_ _05944_ _06137_ VGND VGND VPWR VPWR _06315_ sky130_fd_sc_hd__o31a_1
X_23742__333 clknet_1_0__leaf__10199_ VGND VGND VPWR VPWR net459 sky130_fd_sc_hd__inv_2
X_21990_ _06582_ _09213_ VGND VGND VPWR VPWR _09220_ sky130_fd_sc_hd__nor2_8
XTAP_TAPCELL_ROW_68_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_3466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20941_ datamem.data_ram\[55\]\[22\] _07021_ _06621_ datamem.data_ram\[52\]\[22\]
+ _08230_ VGND VGND VPWR VPWR _08231_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_124_3477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32927_ clknet_leaf_173_clk _04349_ VGND VGND VPWR VPWR datamem.data_ram\[0\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23857__420 clknet_1_1__leaf__10219_ VGND VGND VPWR VPWR net546 sky130_fd_sc_hd__inv_2
X_20872_ datamem.data_ram\[51\]\[14\] _07849_ _08161_ _07851_ VGND VGND VPWR VPWR
+ _08162_ sky130_fd_sc_hd__a211o_1
X_32858_ clknet_leaf_54_clk _04280_ VGND VGND VPWR VPWR datamem.data_ram\[11\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22611_ _09511_ _09760_ VGND VGND VPWR VPWR _09761_ sky130_fd_sc_hd__or2_1
X_31809_ clknet_leaf_109_clk _03263_ VGND VGND VPWR VPWR datamem.data_ram\[17\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_127_clk clknet_5_31__leaf_clk VGND VGND VPWR VPWR clknet_leaf_127_clk
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_138_Right_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32789_ clknet_leaf_287_clk _04211_ VGND VGND VPWR VPWR datamem.data_ram\[14\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25330_ _10754_ net4165 _10909_ VGND VGND VPWR VPWR _10911_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22542_ rvcpu.dp.rf.reg_file_arr\[0\]\[12\] rvcpu.dp.rf.reg_file_arr\[1\]\[12\] rvcpu.dp.rf.reg_file_arr\[2\]\[12\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[12\] _09417_ _09585_ VGND VGND VPWR VPWR _09696_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_187_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25261_ _10413_ _10868_ VGND VGND VPWR VPWR _10872_ sky130_fd_sc_hd__and2_1
X_22473_ _09627_ _09628_ _09630_ _09438_ VGND VGND VPWR VPWR _09631_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_98_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_98_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27000_ _11884_ VGND VGND VPWR VPWR _11885_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_17_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24212_ _10276_ VGND VGND VPWR VPWR _02225_ sky130_fd_sc_hd__clkbuf_1
X_21424_ _08628_ VGND VGND VPWR VPWR _08683_ sky130_fd_sc_hd__buf_4
XFILLER_0_60_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25192_ _10733_ net3656 net57 VGND VGND VPWR VPWR _10834_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21355_ rvcpu.dp.plde.funct3E\[1\] rvcpu.dp.plde.funct3E\[0\] rvcpu.dp.plde.funct3E\[2\]
+ VGND VGND VPWR VPWR _08617_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_86_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23291__934 clknet_1_0__leaf__10131_ VGND VGND VPWR VPWR net1060 sky130_fd_sc_hd__inv_2
XFILLER_0_188_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20306_ _07507_ _07552_ _07598_ VGND VGND VPWR VPWR _07599_ sky130_fd_sc_hd__or3_1
XFILLER_0_130_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28951_ _12982_ VGND VGND VPWR VPWR _04258_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold750 rvcpu.dp.pcreg.q\[25\] VGND VGND VPWR VPWR net1900 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21286_ rvcpu.dp.plfd.InstrD\[15\] VGND VGND VPWR VPWR _08548_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_57_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold761 datamem.data_ram\[46\]\[22\] VGND VGND VPWR VPWR net1911 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27902_ _11980_ _12394_ VGND VGND VPWR VPWR _12402_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_57_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold772 rvcpu.dp.rf.reg_file_arr\[5\]\[23\] VGND VGND VPWR VPWR net1922 sky130_fd_sc_hd__dlygate4sd3_1
X_20237_ datamem.data_ram\[54\]\[3\] _07127_ _06966_ datamem.data_ram\[51\]\[3\] VGND
+ VGND VPWR VPWR _07530_ sky130_fd_sc_hd__a22o_1
Xhold783 datamem.data_ram\[46\]\[30\] VGND VGND VPWR VPWR net1933 sky130_fd_sc_hd__dlygate4sd3_1
X_28882_ _12945_ VGND VGND VPWR VPWR _04226_ sky130_fd_sc_hd__clkbuf_1
Xhold794 rvcpu.dp.rf.reg_file_arr\[8\]\[20\] VGND VGND VPWR VPWR net1944 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27833_ _12361_ net3304 _12357_ VGND VGND VPWR VPWR _12362_ sky130_fd_sc_hd__mux2_1
X_20168_ _06596_ _07426_ _07460_ VGND VGND VPWR VPWR _07461_ sky130_fd_sc_hd__a21oi_4
Xhold2140 datamem.data_ram\[13\]\[21\] VGND VGND VPWR VPWR net3290 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2151 rvcpu.dp.rf.reg_file_arr\[31\]\[13\] VGND VGND VPWR VPWR net3301 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2162 datamem.data_ram\[59\]\[14\] VGND VGND VPWR VPWR net3312 sky130_fd_sc_hd__dlygate4sd3_1
X_27764_ _12153_ net2278 _12316_ VGND VGND VPWR VPWR _12322_ sky130_fd_sc_hd__mux2_1
Xhold2173 datamem.data_ram\[63\]\[30\] VGND VGND VPWR VPWR net3323 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_619 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24976_ _10708_ VGND VGND VPWR VPWR _02557_ sky130_fd_sc_hd__clkbuf_1
X_20099_ datamem.data_ram\[5\]\[10\] _06723_ _06828_ datamem.data_ram\[3\]\[10\] _06733_
+ VGND VGND VPWR VPWR _07393_ sky130_fd_sc_hd__o221a_1
XFILLER_0_118_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2184 rvcpu.dp.rf.reg_file_arr\[31\]\[21\] VGND VGND VPWR VPWR net3334 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1450 rvcpu.dp.rf.reg_file_arr\[15\]\[6\] VGND VGND VPWR VPWR net2600 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2195 datamem.data_ram\[34\]\[13\] VGND VGND VPWR VPWR net3345 sky130_fd_sc_hd__dlygate4sd3_1
X_29503_ net865 _01238_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[28\]\[10\] sky130_fd_sc_hd__dfxtp_1
Xhold1461 datamem.data_ram\[41\]\[17\] VGND VGND VPWR VPWR net2611 sky130_fd_sc_hd__dlygate4sd3_1
X_26715_ _11712_ VGND VGND VPWR VPWR _03292_ sky130_fd_sc_hd__clkbuf_1
Xhold1472 rvcpu.dp.rf.reg_file_arr\[27\]\[6\] VGND VGND VPWR VPWR net2622 sky130_fd_sc_hd__dlygate4sd3_1
X_27695_ _12285_ VGND VGND VPWR VPWR _03699_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1483 datamem.data_ram\[5\]\[14\] VGND VGND VPWR VPWR net2633 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_200_5290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1494 datamem.data_ram\[55\]\[28\] VGND VGND VPWR VPWR net2644 sky130_fd_sc_hd__dlygate4sd3_1
X_29434_ net796 _01169_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[30\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_26646_ _11089_ _11663_ VGND VGND VPWR VPWR _11670_ sky130_fd_sc_hd__and2_1
XFILLER_0_169_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14660_ net2947 _13229_ _13214_ VGND VGND VPWR VPWR _13230_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_197_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_211_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0__10246_ _10246_ VGND VGND VPWR VPWR clknet_0__10246_ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_0_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22809_ rvcpu.dp.rf.reg_file_arr\[12\]\[26\] rvcpu.dp.rf.reg_file_arr\[13\]\[26\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[26\] rvcpu.dp.rf.reg_file_arr\[15\]\[26\] _09464_
+ _09467_ VGND VGND VPWR VPWR _09949_ sky130_fd_sc_hd__mux4_1
X_29365_ clknet_leaf_206_clk _01100_ VGND VGND VPWR VPWR datamem.data_ram\[60\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_118_clk clknet_5_27__leaf_clk VGND VGND VPWR VPWR clknet_leaf_118_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_156_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14591_ rvcpu.dp.plmw.RdW\[4\] VGND VGND VPWR VPWR _13176_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_0_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26577_ _10733_ net2924 _11629_ VGND VGND VPWR VPWR _11634_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_105_Right_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23789_ clknet_1_0__leaf__10203_ VGND VGND VPWR VPWR _10205_ sky130_fd_sc_hd__buf_1
XFILLER_0_223_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16330_ net1965 _14428_ _14525_ VGND VGND VPWR VPWR _14529_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28316_ _12631_ VGND VGND VPWR VPWR _03974_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__10177_ _10177_ VGND VGND VPWR VPWR clknet_0__10177_ sky130_fd_sc_hd__clkbuf_16
X_25528_ _10724_ net3375 net54 VGND VGND VPWR VPWR _11022_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29296_ clknet_leaf_1_clk _01031_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD1E\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28247_ _12593_ VGND VGND VPWR VPWR _03943_ sky130_fd_sc_hd__clkbuf_1
X_16261_ _14492_ VGND VGND VPWR VPWR _01905_ sky130_fd_sc_hd__clkbuf_1
X_25459_ _09351_ _10935_ _10052_ VGND VGND VPWR VPWR _10985_ sky130_fd_sc_hd__and3_2
XFILLER_0_125_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18000_ _05321_ rvcpu.dp.SrcBFW_Mux.y\[3\] _05369_ VGND VGND VPWR VPWR _05370_ sky130_fd_sc_hd__o21a_2
X_15212_ _13304_ _13546_ _13465_ _13607_ VGND VGND VPWR VPWR _13754_ sky130_fd_sc_hd__a211o_1
X_23912__469 clknet_1_1__leaf__10225_ VGND VGND VPWR VPWR net595 sky130_fd_sc_hd__inv_2
X_28178_ _12556_ VGND VGND VPWR VPWR _03911_ sky130_fd_sc_hd__clkbuf_1
X_16192_ _14446_ VGND VGND VPWR VPWR _01936_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_11_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15143_ _13524_ _13642_ _13423_ VGND VGND VPWR VPWR _13687_ sky130_fd_sc_hd__a21o_1
X_27129_ _11963_ VGND VGND VPWR VPWR _11964_ sky130_fd_sc_hd__buf_2
XFILLER_0_209_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30140_ net502 _01875_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[10\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_15074_ _13504_ _13619_ _13515_ _13521_ VGND VGND VPWR VPWR _13620_ sky130_fd_sc_hd__a211o_1
X_19951_ datamem.data_ram\[52\]\[18\] _06619_ _07241_ _07244_ VGND VGND VPWR VPWR
+ _07245_ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_207_5455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18902_ _05701_ _05678_ _05694_ VGND VGND VPWR VPWR _06243_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_207_5466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30071_ net433 _01806_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[12\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_19882_ _07176_ VGND VGND VPWR VPWR _07177_ sky130_fd_sc_hd__clkbuf_8
X_18833_ _05658_ _06030_ _05734_ VGND VGND VPWR VPWR _06179_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_184_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_4334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_160_4345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_5267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23268__914 clknet_1_1__leaf__10128_ VGND VGND VPWR VPWR net1040 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_199_5278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18764_ _05693_ _06113_ VGND VGND VPWR VPWR _06114_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15976_ _14325_ VGND VGND VPWR VPWR _02039_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17715_ _05132_ VGND VGND VPWR VPWR _01183_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14927_ _13470_ _13471_ _13473_ _13474_ _13475_ VGND VGND VPWR VPWR _13476_ sky130_fd_sc_hd__o221a_1
X_18695_ _05417_ _05784_ VGND VGND VPWR VPWR _06049_ sky130_fd_sc_hd__nor2_1
X_30973_ clknet_leaf_162_clk _02708_ VGND VGND VPWR VPWR datamem.data_ram\[39\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_78 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32712_ clknet_leaf_171_clk _04134_ VGND VGND VPWR VPWR datamem.data_ram\[17\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_63_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17646_ net2014 _13219_ _05093_ VGND VGND VPWR VPWR _05096_ sky130_fd_sc_hd__mux2_1
X_14858_ _13291_ _13409_ VGND VGND VPWR VPWR _13410_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_63_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32643_ clknet_leaf_164_clk _04065_ VGND VGND VPWR VPWR datamem.data_ram\[1\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_109_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_109_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_202_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_4285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17577_ _05059_ VGND VGND VPWR VPWR _01248_ sky130_fd_sc_hd__clkbuf_1
X_14789_ _13296_ _13281_ VGND VGND VPWR VPWR _13342_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_158_4296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19316_ _06611_ VGND VGND VPWR VPWR _06612_ sky130_fd_sc_hd__buf_8
XFILLER_0_175_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16528_ _14128_ _04465_ VGND VGND VPWR VPWR _04502_ sky130_fd_sc_hd__nand2_4
XFILLER_0_45_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32574_ clknet_leaf_271_clk _03996_ VGND VGND VPWR VPWR datamem.data_ram\[22\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31525_ clknet_leaf_68_clk net1153 VGND VGND VPWR VPWR rvcpu.dp.plem.PCPlus4M\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_19247_ _06547_ _06550_ VGND VGND VPWR VPWR _06551_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16459_ _13176_ rvcpu.dp.plmw.RdW\[3\] _13174_ VGND VGND VPWR VPWR _04465_ sky130_fd_sc_hd__and3b_2
XFILLER_0_128_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23240__888 clknet_1_1__leaf__10126_ VGND VGND VPWR VPWR net1014 sky130_fd_sc_hd__inv_2
XFILLER_0_186_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19178_ _06473_ _06476_ _06481_ _06488_ _06480_ VGND VGND VPWR VPWR _06491_ sky130_fd_sc_hd__a311o_1
X_31456_ clknet_leaf_5_clk rvcpu.dp.SrcBFW_Mux.y\[14\] VGND VGND VPWR VPWR rvcpu.dp.plem.WriteDataM\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_3292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18129_ _05490_ _05493_ VGND VGND VPWR VPWR _05495_ sky130_fd_sc_hd__or2_1
X_30407_ net745 _02142_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[31\]\[18\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_93_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31387_ clknet_leaf_40_clk _03090_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCE\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21140_ datamem.data_ram\[56\]\[23\] _06644_ VGND VGND VPWR VPWR _08429_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30338_ net684 _02073_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[4\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_23586__207 clknet_1_0__leaf__10177_ VGND VGND VPWR VPWR net333 sky130_fd_sc_hd__inv_2
XFILLER_0_223_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21071_ datamem.data_ram\[58\]\[7\] _06930_ _06946_ datamem.data_ram\[57\]\[7\] _08359_
+ VGND VGND VPWR VPWR _08360_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30269_ net623 _02004_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[6\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_32008_ clknet_leaf_128_clk _03430_ VGND VGND VPWR VPWR datamem.data_ram\[27\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_20022_ datamem.data_ram\[40\]\[2\] _06935_ _06946_ datamem.data_ram\[41\]\[2\] _07315_
+ VGND VGND VPWR VPWR _07316_ sky130_fd_sc_hd__a221o_1
XFILLER_0_158_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_3517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_3528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_207_Right_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24830_ _10400_ net3540 _10621_ VGND VGND VPWR VPWR _10629_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24761_ _10590_ VGND VGND VPWR VPWR _02460_ sky130_fd_sc_hd__clkbuf_1
X_21973_ rvcpu.dp.rf.reg_file_arr\[0\]\[31\] rvcpu.dp.rf.reg_file_arr\[1\]\[31\] rvcpu.dp.rf.reg_file_arr\[2\]\[31\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[31\] _08535_ _08552_ VGND VGND VPWR VPWR _09204_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_87_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20924_ _08212_ _08213_ _07821_ VGND VGND VPWR VPWR _08214_ sky130_fd_sc_hd__mux2_1
X_27480_ _12170_ VGND VGND VPWR VPWR _03599_ sky130_fd_sc_hd__clkbuf_1
X_24692_ _10553_ VGND VGND VPWR VPWR _02428_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_179_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26431_ _11524_ rvcpu.ALUResultE\[16\] _11193_ _11526_ VGND VGND VPWR VPWR _11565_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_193_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23643_ _09285_ net4112 _10182_ VGND VGND VPWR VPWR _10188_ sky130_fd_sc_hd__mux2_1
X_24152__655 clknet_1_0__leaf__10263_ VGND VGND VPWR VPWR net781 sky130_fd_sc_hd__inv_2
X_20855_ _08139_ _08143_ _08144_ VGND VGND VPWR VPWR _08145_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29150_ _13091_ VGND VGND VPWR VPWR _04348_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26362_ _11086_ _11511_ VGND VGND VPWR VPWR _11515_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20786_ datamem.data_ram\[16\]\[30\] _07828_ _07839_ VGND VGND VPWR VPWR _08076_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_147_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28101_ _12515_ VGND VGND VPWR VPWR _03875_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_46_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25313_ _10901_ VGND VGND VPWR VPWR _02701_ sky130_fd_sc_hd__clkbuf_1
X_29081_ _12762_ net2433 _13049_ VGND VGND VPWR VPWR _13055_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_475 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22525_ rvcpu.dp.rf.reg_file_arr\[4\]\[11\] rvcpu.dp.rf.reg_file_arr\[5\]\[11\] rvcpu.dp.rf.reg_file_arr\[6\]\[11\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[11\] _09386_ _09419_ VGND VGND VPWR VPWR _09680_
+ sky130_fd_sc_hd__mux4_1
X_26293_ _11479_ VGND VGND VPWR VPWR _03103_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_228_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28032_ _12478_ VGND VGND VPWR VPWR _03843_ sky130_fd_sc_hd__clkbuf_1
X_25244_ _10733_ net3129 net55 VGND VGND VPWR VPWR _10862_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22456_ rvcpu.dp.rf.reg_file_arr\[24\]\[8\] rvcpu.dp.rf.reg_file_arr\[25\]\[8\] rvcpu.dp.rf.reg_file_arr\[26\]\[8\]
+ rvcpu.dp.rf.reg_file_arr\[27\]\[8\] _09393_ _09395_ VGND VGND VPWR VPWR _09614_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_165_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_798 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21407_ _08663_ _08664_ _08666_ _08652_ VGND VGND VPWR VPWR _08667_ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25175_ _10823_ VGND VGND VPWR VPWR _02641_ sky130_fd_sc_hd__clkbuf_1
X_22387_ _09528_ _09548_ _09426_ VGND VGND VPWR VPWR _09549_ sky130_fd_sc_hd__a21o_1
XFILLER_0_206_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21338_ rvcpu.ALUResultE\[1\] rvcpu.ALUResultE\[2\] rvcpu.ALUResultE\[3\] rvcpu.ALUResultE\[4\]
+ VGND VGND VPWR VPWR _08600_ sky130_fd_sc_hd__or4_1
X_29983_ net353 _01718_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[14\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_23749__339 clknet_1_1__leaf__10200_ VGND VGND VPWR VPWR net465 sky130_fd_sc_hd__inv_2
XFILLER_0_124_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28934_ _12760_ net3454 _12968_ VGND VGND VPWR VPWR _12973_ sky130_fd_sc_hd__mux2_1
X_21269_ _08522_ VGND VGND VPWR VPWR _08531_ sky130_fd_sc_hd__clkbuf_4
X_24057_ clknet_1_1__leaf__10244_ VGND VGND VPWR VPWR _10247_ sky130_fd_sc_hd__buf_1
Xhold580 datamem.data_ram\[10\]\[6\] VGND VGND VPWR VPWR net1730 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold591 datamem.data_ram\[14\]\[0\] VGND VGND VPWR VPWR net1741 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28865_ _12936_ VGND VGND VPWR VPWR _04218_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_216_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_194_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_202_5341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27816_ _12151_ net3171 net78 VGND VGND VPWR VPWR _12351_ sky130_fd_sc_hd__mux2_1
X_15830_ _14246_ VGND VGND VPWR VPWR _02106_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_202_5352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28796_ _12741_ net2776 net70 VGND VGND VPWR VPWR _12900_ sky130_fd_sc_hd__mux2_1
XFILLER_0_218_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27747_ _12136_ net3816 _12307_ VGND VGND VPWR VPWR _12313_ sky130_fd_sc_hd__mux2_1
X_15761_ _14209_ VGND VGND VPWR VPWR _02146_ sky130_fd_sc_hd__clkbuf_1
X_24959_ _10390_ net4171 _10696_ VGND VGND VPWR VPWR _10699_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_194_5142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17500_ _05018_ VGND VGND VPWR VPWR _01292_ sky130_fd_sc_hd__clkbuf_1
Xhold1280 rvcpu.dp.rf.reg_file_arr\[4\]\[15\] VGND VGND VPWR VPWR net2430 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_194_5153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14712_ _13268_ VGND VGND VPWR VPWR _13269_ sky130_fd_sc_hd__clkbuf_8
Xhold1291 datamem.data_ram\[16\]\[13\] VGND VGND VPWR VPWR net2441 sky130_fd_sc_hd__dlygate4sd3_1
X_18480_ _05768_ _05761_ VGND VGND VPWR VPWR _05842_ sky130_fd_sc_hd__nand2_1
X_27678_ _12091_ net2927 net51 VGND VGND VPWR VPWR _12276_ sky130_fd_sc_hd__mux2_1
X_15692_ _14165_ VGND VGND VPWR VPWR _02171_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_213_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_420 _06769_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_431 _06790_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_197_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29417_ clknet_leaf_12_clk _01152_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD2E\[28\] sky130_fd_sc_hd__dfxtp_1
X_17431_ _14145_ net4118 _04974_ VGND VGND VPWR VPWR _04982_ sky130_fd_sc_hd__mux2_1
XANTENNA_442 _07023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26629_ _10070_ _11659_ _11660_ net1336 VGND VGND VPWR VPWR _03258_ sky130_fd_sc_hd__a22o_1
X_14643_ _13216_ VGND VGND VPWR VPWR _13217_ sky130_fd_sc_hd__clkbuf_8
XANTENNA_453 _08124_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_170_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_464 _08744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_475 _09313_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_196_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_184_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_486 _09478_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_497 _10297_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17362_ _04945_ VGND VGND VPWR VPWR _01357_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_16_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__10129_ clknet_0__10129_ VGND VGND VPWR VPWR clknet_1_1__leaf__10129_
+ sky130_fd_sc_hd__clkbuf_16
X_29348_ clknet_leaf_199_clk _01083_ VGND VGND VPWR VPWR datamem.data_ram\[61\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19101_ _06421_ _06422_ VGND VGND VPWR VPWR _06423_ sky130_fd_sc_hd__nand2_1
X_16313_ _14519_ VGND VGND VPWR VPWR _01880_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_153_4160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_211_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17293_ net4330 _13200_ _04902_ VGND VGND VPWR VPWR _04909_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29279_ _09305_ net2550 _13159_ VGND VGND VPWR VPWR _13161_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_153_4171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31310_ clknet_leaf_47_clk _03013_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCPlus4E\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_19032_ rvcpu.dp.plde.ImmExtE\[1\] rvcpu.dp.plde.PCE\[1\] VGND VGND VPWR VPWR _06363_
+ sky130_fd_sc_hd__and2_1
X_16244_ _14481_ VGND VGND VPWR VPWR _01919_ sky130_fd_sc_hd__clkbuf_1
X_32290_ clknet_leaf_229_clk _03712_ VGND VGND VPWR VPWR datamem.data_ram\[32\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_551 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_209_5506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31241_ clknet_leaf_35_clk net1824 VGND VGND VPWR VPWR rvcpu.dp.plfd.PCD\[30\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_209_5517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16175_ net2533 _14434_ _14422_ VGND VGND VPWR VPWR _14435_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15126_ _13296_ _13347_ VGND VGND VPWR VPWR _13671_ sky130_fd_sc_hd__nor2_2
X_31172_ clknet_leaf_25_clk rvcpu.ALUResultE\[31\] VGND VGND VPWR VPWR rvcpu.dp.plem.ALUResultM\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30123_ net485 _01858_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[10\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_15057_ _13328_ _13447_ VGND VGND VPWR VPWR _13604_ sky130_fd_sc_hd__nand2_2
X_19934_ _06583_ _07121_ _07228_ VGND VGND VPWR VPWR _04426_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_120_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2909 datamem.data_ram\[50\]\[29\] VGND VGND VPWR VPWR net4059 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_43_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_183_4890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30054_ net416 _01789_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[12\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_19865_ datamem.data_ram\[14\]\[1\] _07159_ _06949_ datamem.data_ram\[9\]\[1\] VGND
+ VGND VPWR VPWR _07160_ sky130_fd_sc_hd__a22o_1
XFILLER_0_207_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18816_ _06136_ _05830_ _06140_ _06162_ VGND VGND VPWR VPWR _06163_ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19796_ datamem.data_ram\[61\]\[9\] _06663_ _06706_ datamem.data_ram\[63\]\[9\] VGND
+ VGND VPWR VPWR _07091_ sky130_fd_sc_hd__o22a_1
XFILLER_0_208_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_121_3403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18747_ _05332_ _05974_ VGND VGND VPWR VPWR _06098_ sky130_fd_sc_hd__nand2_1
X_15959_ _14316_ VGND VGND VPWR VPWR _02047_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_218_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_179_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18678_ _05444_ _05974_ VGND VGND VPWR VPWR _06033_ sky130_fd_sc_hd__nand2_1
X_30956_ clknet_leaf_279_clk _02691_ VGND VGND VPWR VPWR datamem.data_ram\[3\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_994 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_82_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17629_ net2683 _13194_ _05082_ VGND VGND VPWR VPWR _05087_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_82_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30887_ clknet_leaf_203_clk _02622_ VGND VGND VPWR VPWR datamem.data_ram\[42\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20640_ datamem.data_ram\[22\]\[29\] _06682_ _06806_ datamem.data_ram\[20\]\[29\]
+ VGND VGND VPWR VPWR _07931_ sky130_fd_sc_hd__o22a_1
XFILLER_0_74_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32626_ clknet_leaf_93_clk _04048_ VGND VGND VPWR VPWR datamem.data_ram\[1\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_3343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_190_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32557_ clknet_leaf_237_clk _03979_ VGND VGND VPWR VPWR datamem.data_ram\[22\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_20571_ _06917_ VGND VGND VPWR VPWR _07862_ sky130_fd_sc_hd__buf_4
XFILLER_0_160_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31508_ clknet_leaf_51_clk net1157 VGND VGND VPWR VPWR rvcpu.dp.plem.PCPlus4M\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22310_ _09461_ _09468_ _09471_ _09474_ VGND VGND VPWR VPWR _09475_ sky130_fd_sc_hd__o211a_1
XFILLER_0_160_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32488_ clknet_leaf_183_clk _03910_ VGND VGND VPWR VPWR datamem.data_ram\[25\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22241_ rvcpu.dp.rf.reg_file_arr\[16\]\[0\] rvcpu.dp.rf.reg_file_arr\[17\]\[0\] rvcpu.dp.rf.reg_file_arr\[18\]\[0\]
+ rvcpu.dp.rf.reg_file_arr\[19\]\[0\] _09406_ _09395_ VGND VGND VPWR VPWR _09407_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31439_ _00002_ _00003_ VGND VGND VPWR VPWR rvcpu.dp.Cout sky130_fd_sc_hd__dlxtn_1
XFILLER_0_131_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22172_ _09357_ VGND VGND VPWR VPWR _01104_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21123_ _07820_ _08409_ _08411_ _07867_ VGND VGND VPWR VPWR _08412_ sky130_fd_sc_hd__o211a_1
XFILLER_0_160_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26980_ _11837_ _11866_ VGND VGND VPWR VPWR _11874_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25931_ net1867 _11275_ _11273_ _11285_ VGND VGND VPWR VPWR _02935_ sky130_fd_sc_hd__o211a_1
X_21054_ datamem.data_ram\[36\]\[31\] datamem.data_ram\[37\]\[31\] _07825_ VGND VGND
+ VPWR VPWR _08343_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20005_ _06752_ _07282_ _07287_ _07298_ VGND VGND VPWR VPWR _07299_ sky130_fd_sc_hd__a31o_1
X_28650_ _12749_ net3016 _12814_ VGND VGND VPWR VPWR _12822_ sky130_fd_sc_hd__mux2_1
XFILLER_0_199_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25862_ rvcpu.dp.plfd.PCPlus4D\[28\] _11241_ _08598_ VGND VGND VPWR VPWR _11242_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27601_ _12145_ net3488 net81 VGND VGND VPWR VPWR _12235_ sky130_fd_sc_hd__mux2_1
X_23941__495 clknet_1_0__leaf__10228_ VGND VGND VPWR VPWR net621 sky130_fd_sc_hd__inv_2
X_24813_ _10454_ net2544 _10612_ VGND VGND VPWR VPWR _10620_ sky130_fd_sc_hd__mux2_1
X_28581_ _12766_ net3481 _12777_ VGND VGND VPWR VPWR _12785_ sky130_fd_sc_hd__mux2_1
X_25793_ _11185_ _11186_ _11157_ VGND VGND VPWR VPWR _11187_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27532_ _12198_ VGND VGND VPWR VPWR _03623_ sky130_fd_sc_hd__clkbuf_1
X_24744_ _10581_ VGND VGND VPWR VPWR _02452_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_190_Right_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21956_ _08695_ _09187_ _08579_ VGND VGND VPWR VPWR _09188_ sky130_fd_sc_hd__a21o_1
XFILLER_0_179_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20907_ _08185_ _08189_ _07071_ _08196_ VGND VGND VPWR VPWR _08197_ sky130_fd_sc_hd__a211o_1
X_27463_ _12083_ net3664 net83 VGND VGND VPWR VPWR _12161_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24675_ _10544_ VGND VGND VPWR VPWR _02420_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21887_ rvcpu.dp.rf.reg_file_arr\[0\]\[26\] rvcpu.dp.rf.reg_file_arr\[1\]\[26\] rvcpu.dp.rf.reg_file_arr\[2\]\[26\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[26\] _08550_ _08554_ VGND VGND VPWR VPWR _09123_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_104_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23182__853 clknet_1_0__leaf__10111_ VGND VGND VPWR VPWR net979 sky130_fd_sc_hd__inv_2
XFILLER_0_204_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_194_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29202_ _09325_ net2004 _13112_ VGND VGND VPWR VPWR _13119_ sky130_fd_sc_hd__mux2_1
X_26414_ net1690 _11268_ _11552_ _11553_ _10041_ VGND VGND VPWR VPWR _03150_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_104_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27394_ _12080_ net2893 net85 VGND VGND VPWR VPWR _12117_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20838_ datamem.data_ram\[31\]\[14\] _07832_ _08127_ _07821_ VGND VGND VPWR VPWR
+ _08128_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_13_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29133_ _13082_ VGND VGND VPWR VPWR _04340_ sky130_fd_sc_hd__clkbuf_1
X_26345_ _10048_ _11507_ _11508_ net1310 VGND VGND VPWR VPWR _03126_ sky130_fd_sc_hd__a22o_1
XFILLER_0_182_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20769_ _06604_ _07872_ VGND VGND VPWR VPWR _08059_ sky130_fd_sc_hd__nor2_1
XFILLER_0_181_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23454__104 clknet_1_0__leaf__10156_ VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__inv_2
X_22508_ rvcpu.dp.rf.reg_file_arr\[8\]\[10\] rvcpu.dp.rf.reg_file_arr\[10\]\[10\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[10\] rvcpu.dp.rf.reg_file_arr\[11\]\[10\] _09418_
+ _09485_ VGND VGND VPWR VPWR _09664_ sky130_fd_sc_hd__mux4_1
X_29064_ _09284_ net3392 net65 VGND VGND VPWR VPWR _13046_ sky130_fd_sc_hd__mux2_1
X_26276_ _11470_ VGND VGND VPWR VPWR _03095_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23488_ clknet_1_0__leaf__10152_ VGND VGND VPWR VPWR _10160_ sky130_fd_sc_hd__buf_1
XFILLER_0_18_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28015_ _12469_ VGND VGND VPWR VPWR _03835_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_220_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25227_ _10760_ net3852 _10848_ VGND VGND VPWR VPWR _10853_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22439_ _09451_ _09597_ _09404_ VGND VGND VPWR VPWR _09598_ sky130_fd_sc_hd__o21a_1
XFILLER_0_150_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23983__518 clknet_1_0__leaf__10239_ VGND VGND VPWR VPWR net644 sky130_fd_sc_hd__inv_2
X_23534__161 clknet_1_0__leaf__10171_ VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__inv_2
XFILLER_0_60_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25158_ _10570_ _10601_ _10705_ VGND VGND VPWR VPWR _10812_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_131_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17980_ _05179_ _05180_ rvcpu.dp.plde.RD2E\[6\] VGND VGND VPWR VPWR _05351_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_204_5403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25089_ _10739_ net3054 _10768_ VGND VGND VPWR VPWR _10776_ sky130_fd_sc_hd__mux2_1
X_29966_ net336 _01701_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[15\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_179_Left_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16931_ net4290 _14482_ _04706_ VGND VGND VPWR VPWR _04716_ sky130_fd_sc_hd__mux2_1
X_28917_ _12696_ net3838 _12959_ VGND VGND VPWR VPWR _12964_ sky130_fd_sc_hd__mux2_1
X_29897_ net275 _01632_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[17\]\[28\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_196_5204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19650_ _06945_ VGND VGND VPWR VPWR _06946_ sky130_fd_sc_hd__buf_4
X_16862_ _04679_ VGND VGND VPWR VPWR _01607_ sky130_fd_sc_hd__clkbuf_1
X_28848_ _12927_ VGND VGND VPWR VPWR _04210_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_217_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_204_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24020__552 clknet_1_0__leaf__10242_ VGND VGND VPWR VPWR net678 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_221_5794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18601_ _05956_ _05809_ _05958_ VGND VGND VPWR VPWR _05959_ sky130_fd_sc_hd__and3_1
X_15813_ net2024 _13184_ _14236_ VGND VGND VPWR VPWR _14238_ sky130_fd_sc_hd__mux2_1
X_19581_ datamem.data_ram\[35\]\[8\] _06632_ _06669_ datamem.data_ram\[39\]\[8\] VGND
+ VGND VPWR VPWR _06877_ sky130_fd_sc_hd__o22a_1
X_28779_ _12758_ net2654 _12887_ VGND VGND VPWR VPWR _12891_ sky130_fd_sc_hd__mux2_1
X_16793_ net4199 _14480_ _04634_ VGND VGND VPWR VPWR _04643_ sky130_fd_sc_hd__mux2_1
XFILLER_0_176_1282 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30810_ clknet_leaf_136_clk _02545_ VGND VGND VPWR VPWR datamem.data_ram\[45\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_18532_ _05891_ _05892_ _05674_ VGND VGND VPWR VPWR _05893_ sky130_fd_sc_hd__mux2_1
XFILLER_0_220_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15744_ _14133_ net3964 _14199_ VGND VGND VPWR VPWR _14201_ sky130_fd_sc_hd__mux2_1
X_31790_ clknet_leaf_103_clk _03244_ VGND VGND VPWR VPWR datamem.data_ram\[8\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30741_ clknet_leaf_148_clk _02476_ VGND VGND VPWR VPWR datamem.data_ram\[48\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_18463_ _05667_ _05683_ VGND VGND VPWR VPWR _05826_ sky130_fd_sc_hd__nand2_1
XFILLER_0_169_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_155_4211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15675_ _13216_ VGND VGND VPWR VPWR _14154_ sky130_fd_sc_hd__buf_4
XFILLER_0_75_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_201_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_155_4222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23306__947 clknet_1_0__leaf__10133_ VGND VGND VPWR VPWR net1073 sky130_fd_sc_hd__inv_2
XANTENNA_250 _13195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_261 _13213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17414_ _04972_ VGND VGND VPWR VPWR _01332_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_272 _13235_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_188_Left_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_184_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14626_ _13203_ VGND VGND VPWR VPWR _13204_ sky130_fd_sc_hd__buf_4
X_18394_ _05741_ _05662_ _05757_ VGND VGND VPWR VPWR _05758_ sky130_fd_sc_hd__a21o_1
XANTENNA_283 _13260_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_30672_ clknet_leaf_189_clk _02407_ VGND VGND VPWR VPWR datamem.data_ram\[50\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_294 _13493_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_151_4108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_151_4119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32411_ clknet_leaf_240_clk _03833_ VGND VGND VPWR VPWR datamem.data_ram\[28\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_17345_ net4444 _13277_ _04901_ VGND VGND VPWR VPWR _04936_ sky130_fd_sc_hd__mux2_1
X_23695__290 clknet_1_1__leaf__10195_ VGND VGND VPWR VPWR net416 sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_40_clk clknet_5_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_40_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_184_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32342_ clknet_leaf_246_clk _03764_ VGND VGND VPWR VPWR datamem.data_ram\[30\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17276_ _14195_ net3946 _04864_ VGND VGND VPWR VPWR _04899_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19015_ _05698_ _06231_ VGND VGND VPWR VPWR _06349_ sky130_fd_sc_hd__or2_1
Xclkload203 clknet_leaf_211_clk VGND VGND VPWR VPWR clkload203/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_181_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_3240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16227_ _13253_ VGND VGND VPWR VPWR _14470_ sky130_fd_sc_hd__buf_4
Xclkload214 clknet_leaf_208_clk VGND VGND VPWR VPWR clkload214/X sky130_fd_sc_hd__clkbuf_4
X_32273_ clknet_leaf_168_clk _03695_ VGND VGND VPWR VPWR datamem.data_ram\[33\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload225 clknet_leaf_164_clk VGND VGND VPWR VPWR clkload225/X sky130_fd_sc_hd__clkbuf_4
Xclkload236 clknet_leaf_116_clk VGND VGND VPWR VPWR clkload236/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_70_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload247 clknet_leaf_150_clk VGND VGND VPWR VPWR clkload247/Y sky130_fd_sc_hd__inv_6
XFILLER_0_12_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31224_ clknet_leaf_39_clk _02927_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCD\[13\] sky130_fd_sc_hd__dfxtp_1
Xclkload258 clknet_leaf_145_clk VGND VGND VPWR VPWR clkload258/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_228_5959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload269 clknet_leaf_132_clk VGND VGND VPWR VPWR clkload269/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_185_4930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16158_ _14423_ VGND VGND VPWR VPWR _01947_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_110_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_185_4941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_110_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15109_ _13387_ _13389_ _13390_ VGND VGND VPWR VPWR _13654_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_75_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_197_Left_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31155_ clknet_leaf_47_clk rvcpu.ALUResultE\[14\] VGND VGND VPWR VPWR rvcpu.dp.plem.ALUResultM\[14\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16089_ _14386_ VGND VGND VPWR VPWR _01979_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_227_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_181_4838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23352__989 clknet_1_0__leaf__10137_ VGND VGND VPWR VPWR net1115 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_181_4849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30106_ net468 _01841_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[11\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_19917_ datamem.data_ram\[39\]\[17\] _07021_ _07210_ _07211_ VGND VGND VPWR VPWR
+ _07212_ sky130_fd_sc_hd__o211a_1
Xhold2706 rvcpu.dp.rf.reg_file_arr\[22\]\[16\] VGND VGND VPWR VPWR net3856 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31086_ clknet_leaf_107_clk _02821_ VGND VGND VPWR VPWR datamem.data_ram\[21\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2717 datamem.data_ram\[4\]\[17\] VGND VGND VPWR VPWR net3867 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_71_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2728 rvcpu.dp.rf.reg_file_arr\[25\]\[24\] VGND VGND VPWR VPWR net3878 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_71_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2739 datamem.data_ram\[13\]\[22\] VGND VGND VPWR VPWR net3889 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30037_ net399 _01772_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[13\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_19848_ datamem.data_ram\[48\]\[1\] _07138_ _06977_ datamem.data_ram\[52\]\[1\] _07142_
+ VGND VGND VPWR VPWR _07143_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_108_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19779_ datamem.data_ram\[34\]\[9\] _06754_ _06738_ datamem.data_ram\[35\]\[9\] _07031_
+ VGND VGND VPWR VPWR _07074_ sky130_fd_sc_hd__o221a_1
XFILLER_0_74_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_108_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21810_ _08813_ _09049_ _08689_ VGND VGND VPWR VPWR _09050_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_140_3856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22790_ _09415_ _09928_ _09930_ _09488_ VGND VGND VPWR VPWR _09931_ sky130_fd_sc_hd__o211a_1
X_31988_ clknet_leaf_119_clk _03410_ VGND VGND VPWR VPWR datamem.data_ram\[37\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_179_4789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_982 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21741_ _08547_ _08982_ _08984_ _08576_ VGND VGND VPWR VPWR _08985_ sky130_fd_sc_hd__o211a_1
X_30939_ clknet_leaf_172_clk _02674_ VGND VGND VPWR VPWR datamem.data_ram\[40\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23246__894 clknet_1_0__leaf__10126_ VGND VGND VPWR VPWR net1020 sky130_fd_sc_hd__inv_2
X_24460_ _10412_ net4094 _10404_ _10419_ VGND VGND VPWR VPWR _02330_ sky130_fd_sc_hd__a31o_1
XFILLER_0_87_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21672_ rvcpu.dp.rf.reg_file_arr\[20\]\[15\] rvcpu.dp.rf.reg_file_arr\[21\]\[15\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[15\] rvcpu.dp.rf.reg_file_arr\[23\]\[15\] _08799_
+ _08800_ VGND VGND VPWR VPWR _08919_ sky130_fd_sc_hd__mux4_2
XFILLER_0_59_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23411_ clknet_1_1__leaf__10152_ VGND VGND VPWR VPWR _10153_ sky130_fd_sc_hd__buf_1
XFILLER_0_191_635 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32609_ clknet_leaf_82_clk _04031_ VGND VGND VPWR VPWR datamem.data_ram\[20\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_20623_ datamem.data_ram\[15\]\[13\] _06944_ _07913_ rvcpu.dp.plem.ALUResultM\[3\]
+ VGND VGND VPWR VPWR _07914_ sky130_fd_sc_hd__o211a_1
XFILLER_0_190_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24391_ _10374_ VGND VGND VPWR VPWR _02306_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_31_clk clknet_5_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_31_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_163_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26130_ net2037 _11397_ VGND VGND VPWR VPWR _11401_ sky130_fd_sc_hd__and2_1
X_20554_ _07844_ VGND VGND VPWR VPWR _07845_ sky130_fd_sc_hd__buf_6
XFILLER_0_11_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26490__44 clknet_1_1__leaf__10267_ VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__inv_2
XFILLER_0_229_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26061_ _11353_ net1351 _11350_ _11359_ VGND VGND VPWR VPWR _02991_ sky130_fd_sc_hd__a31o_1
X_20485_ datamem.data_ram\[58\]\[20\] _06610_ _06600_ _07776_ VGND VGND VPWR VPWR
+ _07777_ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25012_ _10728_ VGND VGND VPWR VPWR _02573_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22224_ rvcpu.dp.plfd.InstrD\[22\] VGND VGND VPWR VPWR _09390_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_203_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29820_ net198 _01555_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[1\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_22155_ _09347_ VGND VGND VPWR VPWR _01097_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_203_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21106_ datamem.data_ram\[18\]\[7\] datamem.data_ram\[19\]\[7\] _06651_ VGND VGND
+ VPWR VPWR _08395_ sky130_fd_sc_hd__mux2_1
XFILLER_0_199_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26963_ _10402_ _10947_ VGND VGND VPWR VPWR _11864_ sky130_fd_sc_hd__or2_1
X_22086_ _09220_ _09293_ _09295_ VGND VGND VPWR VPWR _09300_ sky130_fd_sc_hd__nor3_4
X_29751_ net1097 _01486_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[21\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout120 _00000_ VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_7_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_98_clk clknet_5_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_98_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25914_ net1830 _11275_ _11273_ _11276_ VGND VGND VPWR VPWR _02927_ sky130_fd_sc_hd__o211a_1
XFILLER_0_195_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28702_ _12849_ VGND VGND VPWR VPWR _04142_ sky130_fd_sc_hd__clkbuf_1
X_21037_ datamem.data_ram\[12\]\[31\] datamem.data_ram\[13\]\[31\] _07824_ VGND VGND
+ VPWR VPWR _08326_ sky130_fd_sc_hd__mux2_1
X_29682_ net1028 _01417_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[23\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_26894_ _11813_ net1462 _11809_ _11819_ VGND VGND VPWR VPWR _03364_ sky130_fd_sc_hd__a31o_1
XFILLER_0_22_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28633_ _12766_ net2825 _12805_ VGND VGND VPWR VPWR _12813_ sky130_fd_sc_hd__mux2_1
XFILLER_0_214_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25845_ _11226_ _11227_ VGND VGND VPWR VPWR _11228_ sky130_fd_sc_hd__nor2_1
X_24158__661 clknet_1_1__leaf__10263_ VGND VGND VPWR VPWR net787 sky130_fd_sc_hd__inv_2
X_23564__187 clknet_1_1__leaf__10175_ VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__inv_2
XFILLER_0_97_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28564_ _12702_ net4193 _12768_ VGND VGND VPWR VPWR _12776_ sky130_fd_sc_hd__mux2_1
X_25776_ net1455 _11144_ _11147_ _11173_ VGND VGND VPWR VPWR _02892_ sky130_fd_sc_hd__o211a_1
X_22988_ clknet_1_0__leaf__10080_ VGND VGND VPWR VPWR _10084_ sky130_fd_sc_hd__buf_1
XFILLER_0_158_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27515_ _12189_ VGND VGND VPWR VPWR _03615_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_201_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24727_ _10572_ VGND VGND VPWR VPWR _02444_ sky130_fd_sc_hd__clkbuf_1
X_28495_ _11978_ _12724_ VGND VGND VPWR VPWR _12732_ sky130_fd_sc_hd__and2_1
X_21939_ _08835_ _09171_ VGND VGND VPWR VPWR _09172_ sky130_fd_sc_hd__or2_1
XFILLER_0_179_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_800 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15460_ _13607_ _13465_ _13781_ VGND VGND VPWR VPWR _13990_ sky130_fd_sc_hd__or3b_1
X_27446_ _12149_ net2627 net84 VGND VGND VPWR VPWR _12150_ sky130_fd_sc_hd__mux2_1
X_24658_ _10412_ net1513 _10531_ _10534_ VGND VGND VPWR VPWR _02413_ sky130_fd_sc_hd__a31o_1
X_15391_ _13464_ _13922_ _13923_ VGND VGND VPWR VPWR _13924_ sky130_fd_sc_hd__and3_1
XFILLER_0_167_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27377_ _10724_ net2708 net86 VGND VGND VPWR VPWR _12108_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24589_ _10495_ VGND VGND VPWR VPWR _02383_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_189_5030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_22_clk clknet_5_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_22_clk sky130_fd_sc_hd__clkbuf_8
X_24050__578 clknet_1_0__leaf__10246_ VGND VGND VPWR VPWR net704 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_189_5041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17130_ _14185_ net3282 _04815_ VGND VGND VPWR VPWR _04822_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29116_ _13073_ VGND VGND VPWR VPWR _04332_ sky130_fd_sc_hd__clkbuf_1
X_26328_ _11081_ _11497_ VGND VGND VPWR VPWR _11499_ sky130_fd_sc_hd__and2_1
XFILLER_0_107_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_208_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29047_ _10069_ _13031_ VGND VGND VPWR VPWR _13037_ sky130_fd_sc_hd__and2_1
X_17061_ _04785_ VGND VGND VPWR VPWR _01506_ sky130_fd_sc_hd__clkbuf_1
X_26259_ _11461_ VGND VGND VPWR VPWR _03087_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16012_ net2135 _13275_ _14310_ VGND VGND VPWR VPWR _14344_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_1300 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_223_5845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_223_5856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17963_ rvcpu.dp.plem.ALUResultM\[14\] _05272_ _05270_ _13234_ _05306_ VGND VGND
+ VPWR VPWR _05334_ sky130_fd_sc_hd__a221o_2
X_29949_ net319 _01684_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[15\]\[8\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_89_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_89_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_18_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19702_ datamem.data_ram\[7\]\[0\] _06926_ _06955_ datamem.data_ram\[4\]\[0\] VGND
+ VGND VPWR VPWR _06998_ sky130_fd_sc_hd__a22o_1
X_16914_ _04707_ VGND VGND VPWR VPWR _01583_ sky130_fd_sc_hd__clkbuf_1
X_32960_ clknet_leaf_84_clk _04382_ VGND VGND VPWR VPWR datamem.data_ram\[6\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_17894_ _05266_ VGND VGND VPWR VPWR _05267_ sky130_fd_sc_hd__buf_4
XFILLER_0_217_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31911_ _04422_ net121 VGND VGND VPWR VPWR datamem.rd_data_mem\[16\] sky130_fd_sc_hd__dlxtn_1
X_19633_ _06666_ _06928_ VGND VGND VPWR VPWR _06929_ sky130_fd_sc_hd__nor2_1
X_23050__750 clknet_1_1__leaf__10090_ VGND VGND VPWR VPWR net876 sky130_fd_sc_hd__inv_2
XFILLER_0_217_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16845_ net3898 _14463_ _04670_ VGND VGND VPWR VPWR _04671_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_192_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32891_ clknet_leaf_165_clk _04313_ VGND VGND VPWR VPWR datamem.data_ram\[10\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19564_ _06585_ rvcpu.dp.plem.ALUResultM\[7\] VGND VGND VPWR VPWR _06860_ sky130_fd_sc_hd__nand2_8
X_31842_ clknet_leaf_163_clk _03296_ VGND VGND VPWR VPWR datamem.data_ram\[8\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_16776_ _04611_ VGND VGND VPWR VPWR _04634_ sky130_fd_sc_hd__buf_4
XFILLER_0_220_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18515_ _05860_ _05861_ _05874_ _05876_ VGND VGND VPWR VPWR _05877_ sky130_fd_sc_hd__a211o_1
X_15727_ _13268_ VGND VGND VPWR VPWR _14189_ sky130_fd_sc_hd__buf_4
XFILLER_0_34_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31773_ clknet_leaf_209_clk _03227_ VGND VGND VPWR VPWR datamem.data_ram\[1\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_19495_ datamem.data_ram\[24\]\[16\] _06647_ _06790_ datamem.data_ram\[25\]\[16\]
+ VGND VGND VPWR VPWR _06791_ sky130_fd_sc_hd__o22a_1
XFILLER_0_220_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18446_ _05652_ _00003_ VGND VGND VPWR VPWR _05809_ sky130_fd_sc_hd__nor2_4
X_30724_ clknet_leaf_191_clk _02459_ VGND VGND VPWR VPWR datamem.data_ram\[49\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_15658_ _14142_ VGND VGND VPWR VPWR _02182_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_174_4664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_4675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14609_ net1975 _13190_ _13181_ VGND VGND VPWR VPWR _13191_ sky130_fd_sc_hd__mux2_1
X_18377_ rvcpu.dp.plde.RD1E\[31\] _05266_ _05270_ _13172_ _05273_ VGND VGND VPWR VPWR
+ _05741_ sky130_fd_sc_hd__a221oi_4
X_30655_ clknet_leaf_197_clk _02390_ VGND VGND VPWR VPWR datamem.data_ram\[50\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15589_ net3427 _13210_ _14092_ VGND VGND VPWR VPWR _14102_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_13_clk clknet_5_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_13_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_141_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17328_ _04927_ VGND VGND VPWR VPWR _01381_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_209_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30586_ clknet_leaf_188_clk _02321_ VGND VGND VPWR VPWR datamem.data_ram\[53\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32325_ clknet_leaf_170_clk _03747_ VGND VGND VPWR VPWR datamem.data_ram\[31\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_17259_ _04890_ VGND VGND VPWR VPWR _01413_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_77_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_133_3682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20270_ datamem.data_ram\[38\]\[19\] _06764_ _07024_ datamem.data_ram\[36\]\[19\]
+ VGND VGND VPWR VPWR _07563_ sky130_fd_sc_hd__o22a_1
X_32256_ clknet_leaf_169_clk _03678_ VGND VGND VPWR VPWR datamem.data_ram\[34\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_133_3693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31207_ clknet_leaf_23_clk _02910_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCPlus4D\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_24027__558 clknet_1_1__leaf__10243_ VGND VGND VPWR VPWR net684 sky130_fd_sc_hd__inv_2
XFILLER_0_41_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32187_ clknet_leaf_241_clk _03609_ VGND VGND VPWR VPWR datamem.data_ram\[37\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3204 datamem.data_ram\[54\]\[16\] VGND VGND VPWR VPWR net4354 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3215 datamem.data_ram\[1\]\[9\] VGND VGND VPWR VPWR net4365 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3226 rvcpu.dp.rf.reg_file_arr\[7\]\[7\] VGND VGND VPWR VPWR net4376 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3237 datamem.data_ram\[60\]\[21\] VGND VGND VPWR VPWR net4387 sky130_fd_sc_hd__dlygate4sd3_1
X_31138_ clknet_leaf_214_clk _02873_ VGND VGND VPWR VPWR datamem.data_ram\[4\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2503 datamem.data_ram\[24\]\[19\] VGND VGND VPWR VPWR net3653 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3248 datamem.data_ram\[5\]\[10\] VGND VGND VPWR VPWR net4398 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3259 rvcpu.c.ad.opb5 VGND VGND VPWR VPWR net4409 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2514 datamem.data_ram\[37\]\[25\] VGND VGND VPWR VPWR net3664 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_36_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2525 rvcpu.dp.rf.reg_file_arr\[26\]\[4\] VGND VGND VPWR VPWR net3675 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_36_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2536 rvcpu.dp.rf.reg_file_arr\[28\]\[1\] VGND VGND VPWR VPWR net3686 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31069_ clknet_leaf_159_clk _02804_ VGND VGND VPWR VPWR datamem.data_ram\[9\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_23960_ _09248_ net3913 _10229_ VGND VGND VPWR VPWR _10234_ sky130_fd_sc_hd__mux2_1
Xhold1802 datamem.data_ram\[60\]\[9\] VGND VGND VPWR VPWR net2952 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2547 datamem.data_ram\[34\]\[8\] VGND VGND VPWR VPWR net3697 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_142_3907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1813 rvcpu.dp.rf.reg_file_arr\[12\]\[4\] VGND VGND VPWR VPWR net2963 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2558 datamem.data_ram\[37\]\[15\] VGND VGND VPWR VPWR net3708 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1824 datamem.data_ram\[13\]\[11\] VGND VGND VPWR VPWR net2974 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2569 datamem.data_ram\[6\]\[25\] VGND VGND VPWR VPWR net3719 sky130_fd_sc_hd__dlygate4sd3_1
X_22911_ _07019_ _10042_ _10044_ VGND VGND VPWR VPWR _10045_ sky130_fd_sc_hd__or3_1
XFILLER_0_166_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23483__130 clknet_1_0__leaf__10159_ VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_32_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1835 rvcpu.dp.rf.reg_file_arr\[0\]\[22\] VGND VGND VPWR VPWR net2985 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1846 datamem.data_ram\[26\]\[19\] VGND VGND VPWR VPWR net2996 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1857 rvcpu.dp.rf.reg_file_arr\[25\]\[9\] VGND VGND VPWR VPWR net3007 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1868 datamem.data_ram\[32\]\[26\] VGND VGND VPWR VPWR net3018 sky130_fd_sc_hd__dlygate4sd3_1
X_25630_ _11057_ net1543 _11077_ _11082_ VGND VGND VPWR VPWR _02837_ sky130_fd_sc_hd__a31o_1
Xhold1879 datamem.data_ram\[31\]\[16\] VGND VGND VPWR VPWR net3029 sky130_fd_sc_hd__dlygate4sd3_1
X_22842_ rvcpu.dp.rf.reg_file_arr\[0\]\[28\] rvcpu.dp.rf.reg_file_arr\[1\]\[28\] rvcpu.dp.rf.reg_file_arr\[2\]\[28\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[28\] _09463_ _09637_ VGND VGND VPWR VPWR _09980_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_223_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_190_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25561_ _09350_ _10051_ VGND VGND VPWR VPWR _11039_ sky130_fd_sc_hd__nand2_4
XFILLER_0_116_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22773_ rvcpu.dp.rf.reg_file_arr\[12\]\[24\] rvcpu.dp.rf.reg_file_arr\[13\]\[24\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[24\] rvcpu.dp.rf.reg_file_arr\[15\]\[24\] _09462_
+ _09721_ VGND VGND VPWR VPWR _09915_ sky130_fd_sc_hd__mux4_1
XFILLER_0_17_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27300_ _12061_ net1492 _12053_ _12063_ VGND VGND VPWR VPWR _03526_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_101_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24512_ _10449_ VGND VGND VPWR VPWR _02352_ sky130_fd_sc_hd__clkbuf_1
X_28280_ _12611_ VGND VGND VPWR VPWR _03958_ sky130_fd_sc_hd__clkbuf_1
X_21724_ _08960_ _08964_ _08968_ _08624_ VGND VGND VPWR VPWR _01045_ sky130_fd_sc_hd__o31a_1
XFILLER_0_91_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_900 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25492_ _10814_ net2101 _10999_ VGND VGND VPWR VPWR _11001_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27231_ _12022_ net1386 _12018_ _12027_ VGND VGND VPWR VPWR _03493_ sky130_fd_sc_hd__a31o_1
XFILLER_0_164_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24443_ _10057_ VGND VGND VPWR VPWR _10408_ sky130_fd_sc_hd__buf_2
X_21655_ _08531_ _08902_ _08512_ VGND VGND VPWR VPWR _08903_ sky130_fd_sc_hd__o21a_1
XFILLER_0_191_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27162_ _11970_ _11984_ VGND VGND VPWR VPWR _11987_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_62_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20606_ datamem.data_ram\[62\]\[13\] _06682_ _06671_ datamem.data_ram\[63\]\[13\]
+ _07896_ VGND VGND VPWR VPWR _07897_ sky130_fd_sc_hd__o221a_1
XFILLER_0_163_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24374_ _09330_ net3208 _10357_ VGND VGND VPWR VPWR _10365_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21586_ _08663_ _08834_ _08837_ _08575_ VGND VGND VPWR VPWR _08838_ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26113_ net1676 _11386_ VGND VGND VPWR VPWR _11392_ sky130_fd_sc_hd__and2_1
X_23325_ clknet_1_0__leaf__10130_ VGND VGND VPWR VPWR _10135_ sky130_fd_sc_hd__buf_1
X_27093_ _11825_ _11941_ VGND VGND VPWR VPWR _11943_ sky130_fd_sc_hd__and2_1
X_20537_ _07827_ VGND VGND VPWR VPWR _07828_ sky130_fd_sc_hd__buf_6
XFILLER_0_50_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26044_ _07203_ _10918_ _10897_ VGND VGND VPWR VPWR _11349_ sky130_fd_sc_hd__or3_1
XFILLER_0_160_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20468_ datamem.data_ram\[42\]\[20\] _06609_ _07242_ datamem.data_ram\[41\]\[20\]
+ VGND VGND VPWR VPWR _07760_ sky130_fd_sc_hd__o22a_1
XFILLER_0_63_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22207_ _09376_ VGND VGND VPWR VPWR _01120_ sky130_fd_sc_hd__clkbuf_1
X_23187_ _07132_ VGND VGND VPWR VPWR _10113_ sky130_fd_sc_hd__buf_8
X_20399_ _06595_ _07657_ _07690_ VGND VGND VPWR VPWR _07691_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_101_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23434__85 clknet_1_1__leaf__10155_ VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__inv_2
X_29803_ clknet_leaf_197_clk _01538_ VGND VGND VPWR VPWR datamem.data_ram\[59\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_22138_ _09338_ VGND VGND VPWR VPWR _01089_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_203_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27995_ _12457_ VGND VGND VPWR VPWR _03827_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14960_ _13415_ VGND VGND VPWR VPWR _13509_ sky130_fd_sc_hd__clkbuf_4
X_26946_ _11822_ _11854_ VGND VGND VPWR VPWR _11855_ sky130_fd_sc_hd__and2_1
X_29734_ net1080 _01469_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[21\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_22069_ _09285_ net3586 _09270_ VGND VGND VPWR VPWR _09286_ sky130_fd_sc_hd__mux2_1
Xhold9 rvcpu.dp.plem.ResultSrcM\[0\] VGND VGND VPWR VPWR net1159 sky130_fd_sc_hd__dlygate4sd3_1
X_26877_ _11725_ _11075_ VGND VGND VPWR VPWR _11810_ sky130_fd_sc_hd__nor2_2
X_14891_ _13441_ VGND VGND VPWR VPWR _13442_ sky130_fd_sc_hd__clkbuf_4
X_29665_ net1011 _01400_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[24\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_16630_ _14162_ net4208 _04551_ VGND VGND VPWR VPWR _04557_ sky130_fd_sc_hd__mux2_1
X_25828_ rvcpu.dp.pcreg.q\[22\] _11208_ VGND VGND VPWR VPWR _11214_ sky130_fd_sc_hd__nor2_1
X_28616_ _12702_ net2003 _12796_ VGND VGND VPWR VPWR _12804_ sky130_fd_sc_hd__mux2_1
XFILLER_0_226_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29596_ net950 _01331_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[26\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_16561_ _14162_ net2367 _04514_ VGND VGND VPWR VPWR _04520_ sky130_fd_sc_hd__mux2_1
X_25759_ _11159_ _11160_ _11152_ VGND VGND VPWR VPWR _11161_ sky130_fd_sc_hd__a21o_1
XFILLER_0_186_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28547_ _12766_ net3651 _12752_ VGND VGND VPWR VPWR _12767_ sky130_fd_sc_hd__mux2_1
X_15512_ _14009_ _14038_ _13357_ VGND VGND VPWR VPWR _14039_ sky130_fd_sc_hd__a21oi_1
X_18300_ _05664_ VGND VGND VPWR VPWR _05665_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19280_ rvcpu.dp.plfd.InstrD\[13\] _06577_ rvcpu.dp.plfd.InstrD\[14\] VGND VGND VPWR
+ VPWR _06578_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16492_ _04483_ VGND VGND VPWR VPWR _01797_ sky130_fd_sc_hd__clkbuf_1
X_28478_ _12721_ VGND VGND VPWR VPWR _04046_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_216_5671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_183_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18231_ rvcpu.dp.plde.RD1E\[7\] _05292_ _05341_ VGND VGND VPWR VPWR _05596_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_84_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_216_5682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15443_ _13328_ _13301_ _13858_ VGND VGND VPWR VPWR _13974_ sky130_fd_sc_hd__a21bo_1
X_27429_ _09255_ VGND VGND VPWR VPWR _12138_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_127_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23989__524 clknet_1_0__leaf__10239_ VGND VGND VPWR VPWR net650 sky130_fd_sc_hd__inv_2
X_18162_ rvcpu.dp.plde.RD1E\[25\] _05291_ _05526_ VGND VGND VPWR VPWR _05527_ sky130_fd_sc_hd__o21a_1
X_30440_ net778 _02175_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[29\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_15374_ _13785_ _13501_ _13905_ _13906_ _13907_ VGND VGND VPWR VPWR _13908_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_212_5579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17113_ _14168_ net4065 _04804_ VGND VGND VPWR VPWR _04813_ sky130_fd_sc_hd__mux2_1
X_18093_ _05460_ VGND VGND VPWR VPWR _05461_ sky130_fd_sc_hd__buf_2
X_30371_ net717 _02106_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[3\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32110_ clknet_leaf_120_clk _03532_ VGND VGND VPWR VPWR datamem.data_ram\[58\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap106 net111 VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__clkbuf_2
Xhold409 datamem.data_ram\[2\]\[5\] VGND VGND VPWR VPWR net1559 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap117 _08470_ VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__buf_1
X_17044_ _04776_ VGND VGND VPWR VPWR _01514_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_208_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_225_5907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32041_ clknet_leaf_130_clk _03463_ VGND VGND VPWR VPWR datamem.data_ram\[49\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_146_4007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_1278 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_221_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18995_ _06218_ _06329_ _05698_ VGND VGND VPWR VPWR _06330_ sky130_fd_sc_hd__mux2_1
XFILLER_0_178_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24100__608 clknet_1_1__leaf__10258_ VGND VGND VPWR VPWR net734 sky130_fd_sc_hd__inv_2
XFILLER_0_188_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17946_ _05317_ VGND VGND VPWR VPWR _05318_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_163_4398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1109 datamem.data_ram\[40\]\[22\] VGND VGND VPWR VPWR net2259 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_2_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_119_Right_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_206_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32943_ clknet_leaf_139_clk _04365_ VGND VGND VPWR VPWR datamem.data_ram\[6\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_105_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17877_ rvcpu.dp.plde.Rs1E\[1\] rvcpu.dp.plem.RdM\[1\] VGND VGND VPWR VPWR _05250_
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_105_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19616_ _05391_ _06911_ VGND VGND VPWR VPWR _06912_ sky130_fd_sc_hd__nand2_1
X_16828_ net4010 _14447_ _04659_ VGND VGND VPWR VPWR _04662_ sky130_fd_sc_hd__mux2_1
X_23660__259 clknet_1_1__leaf__10191_ VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__inv_2
X_32874_ clknet_leaf_56_clk _04296_ VGND VGND VPWR VPWR datamem.data_ram\[10\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_176_4715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_176_4726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31825_ clknet_leaf_104_clk _03279_ VGND VGND VPWR VPWR datamem.data_ram\[16\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19547_ datamem.data_ram\[21\]\[24\] _06724_ _06671_ datamem.data_ram\[23\]\[24\]
+ VGND VGND VPWR VPWR _06843_ sky130_fd_sc_hd__o22a_1
XFILLER_0_215_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16759_ _04625_ VGND VGND VPWR VPWR _01664_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_66_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31756_ clknet_leaf_72_clk _03210_ VGND VGND VPWR VPWR datamem.data_ram\[45\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_19478_ datamem.data_ram\[19\]\[16\] _06636_ VGND VGND VPWR VPWR _06774_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18429_ _05780_ _05782_ _05788_ _05792_ VGND VGND VPWR VPWR _05793_ sky130_fd_sc_hd__o211a_1
XFILLER_0_146_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30707_ clknet_leaf_195_clk _02442_ VGND VGND VPWR VPWR datamem.data_ram\[49\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31687_ clknet_leaf_37_clk _03145_ VGND VGND VPWR VPWR rvcpu.dp.pcreg.q\[5\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_150_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_3733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_568 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_3744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21440_ _08509_ _08512_ VGND VGND VPWR VPWR _08699_ sky130_fd_sc_hd__nand2_2
X_30638_ clknet_leaf_142_clk _02373_ VGND VGND VPWR VPWR datamem.data_ram\[51\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_487 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21371_ _08559_ VGND VGND VPWR VPWR _08632_ sky130_fd_sc_hd__buf_4
XFILLER_0_86_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22961__670 clknet_1_1__leaf__10081_ VGND VGND VPWR VPWR net796 sky130_fd_sc_hd__inv_2
X_30569_ clknet_leaf_195_clk _02304_ VGND VGND VPWR VPWR datamem.data_ram\[54\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_20322_ datamem.data_ram\[30\]\[4\] _07159_ _07612_ _07613_ VGND VGND VPWR VPWR _07614_
+ sky130_fd_sc_hd__a211o_1
X_32308_ clknet_leaf_256_clk _03730_ VGND VGND VPWR VPWR datamem.data_ram\[32\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_96_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24090_ _09291_ net2121 _10249_ VGND VGND VPWR VPWR _10257_ sky130_fd_sc_hd__mux2_1
Xhold910 datamem.data_ram\[19\]\[16\] VGND VGND VPWR VPWR net2060 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold921 rvcpu.dp.rf.reg_file_arr\[8\]\[4\] VGND VGND VPWR VPWR net2071 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold932 datamem.data_ram\[35\]\[15\] VGND VGND VPWR VPWR net2082 sky130_fd_sc_hd__dlygate4sd3_1
X_20253_ datamem.data_ram\[40\]\[3\] _06937_ _06958_ datamem.data_ram\[41\]\[3\] _07545_
+ VGND VGND VPWR VPWR _07546_ sky130_fd_sc_hd__a221o_1
Xhold943 rvcpu.dp.rf.reg_file_arr\[3\]\[6\] VGND VGND VPWR VPWR net2093 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold954 rvcpu.dp.rf.reg_file_arr\[29\]\[9\] VGND VGND VPWR VPWR net2104 sky130_fd_sc_hd__dlygate4sd3_1
X_32239_ clknet_leaf_277_clk _03661_ VGND VGND VPWR VPWR datamem.data_ram\[35\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_23057__756 clknet_1_0__leaf__10091_ VGND VGND VPWR VPWR net882 sky130_fd_sc_hd__inv_2
Xhold965 rvcpu.dp.plfd.PCD\[18\] VGND VGND VPWR VPWR net2115 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3001 datamem.data_ram\[58\]\[9\] VGND VGND VPWR VPWR net4151 sky130_fd_sc_hd__dlygate4sd3_1
Xhold976 datamem.data_ram\[13\]\[31\] VGND VGND VPWR VPWR net2126 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3012 datamem.data_ram\[28\]\[10\] VGND VGND VPWR VPWR net4162 sky130_fd_sc_hd__dlygate4sd3_1
Xhold987 rvcpu.dp.rf.reg_file_arr\[3\]\[12\] VGND VGND VPWR VPWR net2137 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3023 datamem.data_ram\[35\]\[20\] VGND VGND VPWR VPWR net4173 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_34_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20184_ datamem.data_ram\[0\]\[11\] _06779_ _06620_ datamem.data_ram\[4\]\[11\] VGND
+ VGND VPWR VPWR _07477_ sky130_fd_sc_hd__o22a_1
Xhold998 rvcpu.dp.rf.reg_file_arr\[19\]\[24\] VGND VGND VPWR VPWR net2148 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_34_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3034 datamem.data_ram\[14\]\[11\] VGND VGND VPWR VPWR net4184 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3045 rvcpu.dp.rf.reg_file_arr\[13\]\[9\] VGND VGND VPWR VPWR net4195 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2300 datamem.data_ram\[49\]\[11\] VGND VGND VPWR VPWR net3450 sky130_fd_sc_hd__dlygate4sd3_1
X_26800_ _11679_ _11762_ VGND VGND VPWR VPWR _11764_ sky130_fd_sc_hd__and2_1
Xhold3056 datamem.data_ram\[54\]\[21\] VGND VGND VPWR VPWR net4206 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2311 datamem.data_ram\[21\]\[23\] VGND VGND VPWR VPWR net3461 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2322 datamem.data_ram\[18\]\[20\] VGND VGND VPWR VPWR net3472 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3067 datamem.data_ram\[39\]\[16\] VGND VGND VPWR VPWR net4217 sky130_fd_sc_hd__dlygate4sd3_1
X_27780_ _12089_ net3645 _12326_ VGND VGND VPWR VPWR _12331_ sky130_fd_sc_hd__mux2_1
XFILLER_0_200_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24992_ _10442_ net3144 _10715_ VGND VGND VPWR VPWR _10717_ sky130_fd_sc_hd__mux2_1
Xhold3078 datamem.data_ram\[25\]\[12\] VGND VGND VPWR VPWR net4228 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2333 datamem.data_ram\[42\]\[11\] VGND VGND VPWR VPWR net3483 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3089 datamem.data_ram\[0\]\[13\] VGND VGND VPWR VPWR net4239 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2344 datamem.data_ram\[33\]\[15\] VGND VGND VPWR VPWR net3494 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1610 rvcpu.dp.rf.reg_file_arr\[12\]\[16\] VGND VGND VPWR VPWR net2760 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2355 datamem.data_ram\[30\]\[25\] VGND VGND VPWR VPWR net3505 sky130_fd_sc_hd__dlygate4sd3_1
X_26731_ _11721_ VGND VGND VPWR VPWR _03299_ sky130_fd_sc_hd__clkbuf_1
Xhold1621 datamem.data_ram\[32\]\[10\] VGND VGND VPWR VPWR net2771 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2366 datamem.data_ram\[3\]\[31\] VGND VGND VPWR VPWR net3516 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1632 rvcpu.dp.rf.reg_file_arr\[27\]\[17\] VGND VGND VPWR VPWR net2782 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2377 datamem.data_ram\[15\]\[9\] VGND VGND VPWR VPWR net3527 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2388 datamem.data_ram\[32\]\[19\] VGND VGND VPWR VPWR net3538 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1643 rvcpu.dp.rf.reg_file_arr\[22\]\[12\] VGND VGND VPWR VPWR net2793 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1654 rvcpu.dp.rf.reg_file_arr\[20\]\[30\] VGND VGND VPWR VPWR net2804 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2399 datamem.data_ram\[12\]\[26\] VGND VGND VPWR VPWR net3549 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1665 datamem.data_ram\[26\]\[9\] VGND VGND VPWR VPWR net2815 sky130_fd_sc_hd__dlygate4sd3_1
X_29450_ net812 _01185_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[30\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_26662_ _10060_ VGND VGND VPWR VPWR _11681_ sky130_fd_sc_hd__clkbuf_4
Xhold1676 datamem.data_ram\[1\]\[28\] VGND VGND VPWR VPWR net2826 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1687 datamem.data_ram\[42\]\[21\] VGND VGND VPWR VPWR net2837 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1698 datamem.data_ram\[51\]\[10\] VGND VGND VPWR VPWR net2848 sky130_fd_sc_hd__dlygate4sd3_1
X_28401_ _12445_ net3461 _12669_ VGND VGND VPWR VPWR _12677_ sky130_fd_sc_hd__mux2_1
X_25613_ _10733_ net3673 net53 VGND VGND VPWR VPWR _11071_ sky130_fd_sc_hd__mux2_1
Xclkbuf_0__10262_ _10262_ VGND VGND VPWR VPWR clknet_0__10262_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_223_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_211_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22825_ _09429_ _09961_ _09963_ VGND VGND VPWR VPWR _09964_ sky130_fd_sc_hd__a21o_1
X_29381_ clknet_leaf_267_clk _01116_ VGND VGND VPWR VPWR datamem.data_ram\[60\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_26593_ _11618_ net1817 _11639_ _11643_ VGND VGND VPWR VPWR _03239_ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28332_ _12371_ net3343 _12632_ VGND VGND VPWR VPWR _12640_ sky130_fd_sc_hd__mux2_1
X_25544_ _10570_ _10960_ _10998_ VGND VGND VPWR VPWR _11030_ sky130_fd_sc_hd__a21oi_4
Xclkbuf_0__10193_ _10193_ VGND VGND VPWR VPWR clknet_0__10193_ sky130_fd_sc_hd__clkbuf_16
X_22756_ _09481_ _09898_ VGND VGND VPWR VPWR _09899_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21707_ rvcpu.dp.rf.reg_file_arr\[16\]\[17\] rvcpu.dp.rf.reg_file_arr\[17\]\[17\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[17\] rvcpu.dp.rf.reg_file_arr\[19\]\[17\] _08703_
+ _08721_ VGND VGND VPWR VPWR _08952_ sky130_fd_sc_hd__mux4_1
X_28263_ _08133_ net106 VGND VGND VPWR VPWR _12602_ sky130_fd_sc_hd__nor2_8
X_25475_ _10076_ _10985_ VGND VGND VPWR VPWR _10994_ sky130_fd_sc_hd__and2_1
XFILLER_0_176_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22687_ _09511_ _09832_ VGND VGND VPWR VPWR _09833_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27214_ _07019_ _11109_ _11839_ VGND VGND VPWR VPWR _12017_ sky130_fd_sc_hd__or3_1
XFILLER_0_75_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_229_6007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24426_ _10395_ VGND VGND VPWR VPWR _02320_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28194_ _12447_ net3150 net46 VGND VGND VPWR VPWR _12565_ sky130_fd_sc_hd__mux2_1
X_21638_ rvcpu.dp.rf.reg_file_arr\[24\]\[13\] rvcpu.dp.rf.reg_file_arr\[25\]\[13\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[13\] rvcpu.dp.rf.reg_file_arr\[27\]\[13\] _08548_
+ _08526_ VGND VGND VPWR VPWR _08887_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_229_6018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27145_ _11974_ net1507 _11964_ _11975_ VGND VGND VPWR VPWR _03459_ sky130_fd_sc_hd__a31o_1
X_24357_ _09291_ net2397 _10348_ VGND VGND VPWR VPWR _10356_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21569_ _08817_ _08819_ _08821_ _08700_ VGND VGND VPWR VPWR _08822_ sky130_fd_sc_hd__a211o_1
XFILLER_0_23_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27076_ _11835_ _11924_ VGND VGND VPWR VPWR _11931_ sky130_fd_sc_hd__and2_1
X_15090_ _13478_ _13480_ _13527_ _13635_ _13438_ VGND VGND VPWR VPWR _13636_ sky130_fd_sc_hd__a41o_1
XFILLER_0_132_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24288_ _10317_ VGND VGND VPWR VPWR _02260_ sky130_fd_sc_hd__clkbuf_1
X_26027_ _11109_ _10980_ VGND VGND VPWR VPWR _11340_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_207_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17800_ _05193_ VGND VGND VPWR VPWR rvcpu.dp.SrcBFW_Mux.y\[4\] sky130_fd_sc_hd__clkbuf_2
X_23880__441 clknet_1_1__leaf__10221_ VGND VGND VPWR VPWR net567 sky130_fd_sc_hd__inv_2
X_18780_ _05805_ _06128_ _05695_ _05703_ VGND VGND VPWR VPWR _06129_ sky130_fd_sc_hd__a2bb2o_1
X_15992_ net2007 _13244_ _14333_ VGND VGND VPWR VPWR _14334_ sky130_fd_sc_hd__mux2_1
X_27978_ _12445_ net1937 _12431_ VGND VGND VPWR VPWR _12446_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_175_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14943_ _13295_ _13432_ VGND VGND VPWR VPWR _13492_ sky130_fd_sc_hd__or2_2
X_29717_ net1063 _01452_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[22\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_17731_ _13244_ net4310 _05140_ VGND VGND VPWR VPWR _05141_ sky130_fd_sc_hd__mux2_1
X_26929_ _11831_ net1598 _11841_ _11844_ VGND VGND VPWR VPWR _03374_ sky130_fd_sc_hd__a31o_1
X_14874_ _13425_ _13336_ VGND VGND VPWR VPWR _13426_ sky130_fd_sc_hd__nor2_1
X_29648_ net994 _01383_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[24\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17662_ _05081_ VGND VGND VPWR VPWR _05104_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_218_5722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19401_ _06696_ VGND VGND VPWR VPWR _06697_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_218_5733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16613_ _14145_ net3790 _04540_ VGND VGND VPWR VPWR _04548_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17593_ _05067_ VGND VGND VPWR VPWR _01240_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_187_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29579_ net933 _01314_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[26\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24056__584 clknet_1_0__leaf__10246_ VGND VGND VPWR VPWR net710 sky130_fd_sc_hd__inv_2
X_31610_ clknet_leaf_25_clk net1173 VGND VGND VPWR VPWR rvcpu.dp.plmw.PCPlus4W\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_16544_ _14145_ net4259 _04503_ VGND VGND VPWR VPWR _04511_ sky130_fd_sc_hd__mux2_1
X_19332_ _06627_ VGND VGND VPWR VPWR _06628_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_171_4601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32590_ clknet_leaf_73_clk _04012_ VGND VGND VPWR VPWR datamem.data_ram\[21\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19263_ _05275_ _05280_ VGND VGND VPWR VPWR _06564_ sky130_fd_sc_hd__and2_1
X_31541_ clknet_leaf_76_clk net1208 VGND VGND VPWR VPWR rvcpu.dp.plem.MemWriteM sky130_fd_sc_hd__dfxtp_1
X_16475_ _04474_ VGND VGND VPWR VPWR _01805_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15426_ _13292_ _13401_ _13628_ _13718_ VGND VGND VPWR VPWR _13957_ sky130_fd_sc_hd__or4_1
X_18214_ _05578_ VGND VGND VPWR VPWR _05579_ sky130_fd_sc_hd__clkbuf_4
X_19194_ _06503_ _06504_ VGND VGND VPWR VPWR _06505_ sky130_fd_sc_hd__xor2_1
XFILLER_0_182_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31472_ clknet_leaf_5_clk rvcpu.dp.SrcBFW_Mux.y\[30\] VGND VGND VPWR VPWR rvcpu.dp.plem.WriteDataM\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30423_ net761 _02158_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[29\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_15357_ _13888_ _13889_ _13891_ _13439_ VGND VGND VPWR VPWR _13892_ sky130_fd_sc_hd__a31o_1
X_18145_ _05506_ _05509_ VGND VGND VPWR VPWR _05510_ sky130_fd_sc_hd__and2_1
XFILLER_0_182_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_169_4541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18076_ _05441_ _05430_ VGND VGND VPWR VPWR _05444_ sky130_fd_sc_hd__and2_1
X_30354_ net700 _02089_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[3\]\[5\] sky130_fd_sc_hd__dfxtp_1
Xhold206 datamem.data_ram\[60\]\[6\] VGND VGND VPWR VPWR net1356 sky130_fd_sc_hd__dlygate4sd3_1
X_15288_ _13604_ _13505_ _13764_ VGND VGND VPWR VPWR _13826_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_169_4552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold217 datamem.data_ram\[47\]\[0\] VGND VGND VPWR VPWR net1367 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_169_4563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold228 datamem.data_ram\[13\]\[7\] VGND VGND VPWR VPWR net1378 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17027_ _04767_ VGND VGND VPWR VPWR _01522_ sky130_fd_sc_hd__clkbuf_1
Xhold239 datamem.data_ram\[39\]\[6\] VGND VGND VPWR VPWR net1389 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_145_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30285_ net631 _02020_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[5\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_165_4449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32024_ clknet_leaf_129_clk _03446_ VGND VGND VPWR VPWR datamem.data_ram\[51\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23413__66 clknet_1_1__leaf__10153_ VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__inv_2
X_18978_ _06313_ _06080_ VGND VGND VPWR VPWR _06314_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23130__806 clknet_1_0__leaf__10106_ VGND VGND VPWR VPWR net932 sky130_fd_sc_hd__inv_2
XFILLER_0_226_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_128_3570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17929_ _05300_ _05301_ VGND VGND VPWR VPWR _05302_ sky130_fd_sc_hd__and2_1
X_23379__1014 clknet_1_1__leaf__10139_ VGND VGND VPWR VPWR net1140 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_68_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20940_ _08227_ _08228_ _08229_ _07822_ _07868_ VGND VGND VPWR VPWR _08230_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_124_3467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32926_ clknet_leaf_3_clk _04348_ VGND VGND VPWR VPWR datamem.data_ram\[0\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_124_3478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_221_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32857_ clknet_leaf_55_clk _04279_ VGND VGND VPWR VPWR datamem.data_ram\[11\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_20871_ datamem.data_ram\[50\]\[14\] _07832_ VGND VGND VPWR VPWR _08161_ sky130_fd_sc_hd__and2_1
XFILLER_0_7_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22610_ rvcpu.dp.rf.reg_file_arr\[16\]\[16\] rvcpu.dp.rf.reg_file_arr\[17\]\[16\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[16\] rvcpu.dp.rf.reg_file_arr\[19\]\[16\] _09512_
+ _09513_ VGND VGND VPWR VPWR _09760_ sky130_fd_sc_hd__mux4_1
X_31808_ clknet_leaf_109_clk _03262_ VGND VGND VPWR VPWR datamem.data_ram\[17\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_221_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_193_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32788_ clknet_leaf_257_clk _04210_ VGND VGND VPWR VPWR datamem.data_ram\[14\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22541_ _09412_ _09690_ _09692_ _09694_ _09413_ VGND VGND VPWR VPWR _09695_ sky130_fd_sc_hd__a221o_1
X_31739_ net188 _03197_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[9\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25260_ _10538_ net1478 _10867_ _10871_ VGND VGND VPWR VPWR _02678_ sky130_fd_sc_hd__a31o_1
XFILLER_0_173_251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22472_ _09534_ _09629_ VGND VGND VPWR VPWR _09630_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_98_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24211_ _09322_ net2704 _10270_ VGND VGND VPWR VPWR _10276_ sky130_fd_sc_hd__mux2_1
X_21423_ _08523_ VGND VGND VPWR VPWR _08682_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_72_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25191_ _10833_ VGND VGND VPWR VPWR _02647_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_228_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21354_ rvcpu.dp.plde.funct3E\[0\] rvcpu.dp.Cout rvcpu.dp.plde.funct3E\[1\] rvcpu.dp.plde.funct3E\[2\]
+ VGND VGND VPWR VPWR _08616_ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20305_ _07227_ _07597_ VGND VGND VPWR VPWR _07598_ sky130_fd_sc_hd__nor2_1
X_28950_ _12741_ net4242 net67 VGND VGND VPWR VPWR _12982_ sky130_fd_sc_hd__mux2_1
Xhold740 rvcpu.dp.plfd.PCPlus4D\[9\] VGND VGND VPWR VPWR net1890 sky130_fd_sc_hd__dlygate4sd3_1
X_21285_ _08532_ VGND VGND VPWR VPWR _08547_ sky130_fd_sc_hd__clkbuf_4
Xhold751 rvcpu.dp.rf.reg_file_arr\[19\]\[13\] VGND VGND VPWR VPWR net1901 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_57_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold762 rvcpu.dp.rf.reg_file_arr\[11\]\[27\] VGND VGND VPWR VPWR net1912 sky130_fd_sc_hd__dlygate4sd3_1
X_27901_ _12391_ net1448 _12393_ _12401_ VGND VGND VPWR VPWR _03789_ sky130_fd_sc_hd__a31o_1
Xhold773 datamem.data_ram\[33\]\[23\] VGND VGND VPWR VPWR net1923 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20236_ _07071_ _07512_ _07517_ _07528_ VGND VGND VPWR VPWR _07529_ sky130_fd_sc_hd__a31o_1
XFILLER_0_124_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_229_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28881_ _12758_ net2877 _12941_ VGND VGND VPWR VPWR _12945_ sky130_fd_sc_hd__mux2_1
Xhold784 rvcpu.dp.rf.reg_file_arr\[6\]\[29\] VGND VGND VPWR VPWR net1934 sky130_fd_sc_hd__dlygate4sd3_1
Xhold795 rvcpu.dp.rf.reg_file_arr\[3\]\[8\] VGND VGND VPWR VPWR net1945 sky130_fd_sc_hd__dlygate4sd3_1
X_27832_ _09309_ VGND VGND VPWR VPWR _12361_ sky130_fd_sc_hd__clkbuf_2
X_20167_ _06712_ _07437_ _07448_ _07459_ _06797_ VGND VGND VPWR VPWR _07460_ sky130_fd_sc_hd__a32o_1
XFILLER_0_216_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2130 datamem.data_ram\[43\]\[25\] VGND VGND VPWR VPWR net3280 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2141 datamem.data_ram\[44\]\[16\] VGND VGND VPWR VPWR net3291 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2152 datamem.data_ram\[8\]\[19\] VGND VGND VPWR VPWR net3302 sky130_fd_sc_hd__dlygate4sd3_1
X_24975_ _10468_ net3260 net101 VGND VGND VPWR VPWR _10708_ sky130_fd_sc_hd__mux2_1
X_20098_ datamem.data_ram\[6\]\[10\] _06718_ _06656_ datamem.data_ram\[1\]\[10\] VGND
+ VGND VPWR VPWR _07392_ sky130_fd_sc_hd__o22a_1
Xhold2163 datamem.data_ram\[18\]\[28\] VGND VGND VPWR VPWR net3313 sky130_fd_sc_hd__dlygate4sd3_1
X_27763_ _12321_ VGND VGND VPWR VPWR _03731_ sky130_fd_sc_hd__clkbuf_1
Xhold2174 datamem.data_ram\[18\]\[18\] VGND VGND VPWR VPWR net3324 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2185 datamem.data_ram\[14\]\[24\] VGND VGND VPWR VPWR net3335 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1440 datamem.data_ram\[6\]\[24\] VGND VGND VPWR VPWR net2590 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1451 datamem.data_ram\[51\]\[15\] VGND VGND VPWR VPWR net2601 sky130_fd_sc_hd__dlygate4sd3_1
X_29502_ net864 _01237_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[28\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_26714_ _10826_ net3516 _11704_ VGND VGND VPWR VPWR _11712_ sky130_fd_sc_hd__mux2_1
Xhold2196 rvcpu.dp.rf.reg_file_arr\[30\]\[5\] VGND VGND VPWR VPWR net3346 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27694_ _12134_ net2570 _12280_ VGND VGND VPWR VPWR _12285_ sky130_fd_sc_hd__mux2_1
Xhold1462 rvcpu.dp.rf.reg_file_arr\[23\]\[7\] VGND VGND VPWR VPWR net2612 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1473 datamem.data_ram\[22\]\[16\] VGND VGND VPWR VPWR net2623 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1484 rvcpu.dp.rf.reg_file_arr\[30\]\[26\] VGND VGND VPWR VPWR net2634 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_200_5291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1495 rvcpu.dp.rf.reg_file_arr\[13\]\[20\] VGND VGND VPWR VPWR net2645 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26645_ _11665_ net1822 _11662_ _11669_ VGND VGND VPWR VPWR _03265_ sky130_fd_sc_hd__a31o_1
X_29433_ net795 _01168_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[30\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0__10245_ _10245_ VGND VGND VPWR VPWR clknet_0__10245_ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_0_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22808_ _09415_ _09945_ _09947_ _09473_ VGND VGND VPWR VPWR _09948_ sky130_fd_sc_hd__o211a_1
X_14590_ rvcpu.dp.plmw.RdW\[3\] VGND VGND VPWR VPWR _13175_ sky130_fd_sc_hd__inv_2
X_26576_ _11633_ VGND VGND VPWR VPWR _03232_ sky130_fd_sc_hd__clkbuf_1
X_29364_ clknet_leaf_180_clk _01099_ VGND VGND VPWR VPWR datamem.data_ram\[61\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_211_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22968__676 clknet_1_1__leaf__10082_ VGND VGND VPWR VPWR net802 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_192_5092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_1288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__10176_ _10176_ VGND VGND VPWR VPWR clknet_0__10176_ sky130_fd_sc_hd__clkbuf_16
X_28315_ _12462_ net3482 net72 VGND VGND VPWR VPWR _12631_ sky130_fd_sc_hd__mux2_1
X_25527_ _10838_ _11020_ _10998_ VGND VGND VPWR VPWR _11021_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_149_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29295_ clknet_leaf_1_clk _01030_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD1E\[2\] sky130_fd_sc_hd__dfxtp_1
X_22739_ _09476_ _09880_ _09882_ _09474_ VGND VGND VPWR VPWR _09883_ sky130_fd_sc_hd__o211a_1
XFILLER_0_165_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28246_ _12447_ net3438 net44 VGND VGND VPWR VPWR _12593_ sky130_fd_sc_hd__mux2_1
X_16260_ net2856 _14426_ _14489_ VGND VGND VPWR VPWR _14492_ sky130_fd_sc_hd__mux2_1
X_25458_ _10983_ VGND VGND VPWR VPWR _10984_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_109_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15211_ _13469_ _13745_ _13749_ _13752_ VGND VGND VPWR VPWR _13753_ sky130_fd_sc_hd__or4_1
X_24409_ _09291_ net3402 _10376_ VGND VGND VPWR VPWR _10384_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28177_ _12430_ net3022 _12555_ VGND VGND VPWR VPWR _12556_ sky130_fd_sc_hd__mux2_1
X_16191_ net1944 _14445_ _14443_ VGND VGND VPWR VPWR _14446_ sky130_fd_sc_hd__mux2_1
X_25389_ _09225_ _10051_ VGND VGND VPWR VPWR _10947_ sky130_fd_sc_hd__nand2_8
XTAP_TAPCELL_ROW_11_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15142_ _13488_ _13685_ _13581_ _13492_ _13527_ VGND VGND VPWR VPWR _13686_ sky130_fd_sc_hd__o41a_1
X_27128_ _07203_ _10326_ _11839_ VGND VGND VPWR VPWR _11963_ sky130_fd_sc_hd__or3_1
XFILLER_0_51_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15073_ _13289_ _13507_ _13511_ VGND VGND VPWR VPWR _13619_ sky130_fd_sc_hd__a21o_1
X_27059_ _11837_ _11911_ VGND VGND VPWR VPWR _11921_ sky130_fd_sc_hd__and2_1
X_19950_ datamem.data_ram\[51\]\[18\] _06633_ _07243_ datamem.data_ram\[49\]\[18\]
+ _06678_ VGND VGND VPWR VPWR _07244_ sky130_fd_sc_hd__o221a_1
X_18901_ _06240_ _06241_ VGND VGND VPWR VPWR _06242_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_691 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_207_5456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30070_ net432 _01805_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[12\]\[25\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_207_5467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19881_ rvcpu.dp.plem.ALUResultM\[7\] _06750_ VGND VGND VPWR VPWR _07176_ sky130_fd_sc_hd__or2_2
X_18832_ _05497_ _05727_ _05730_ _05495_ _06177_ VGND VGND VPWR VPWR _06178_ sky130_fd_sc_hd__a221o_1
X_23726__318 clknet_1_0__leaf__10198_ VGND VGND VPWR VPWR net444 sky130_fd_sc_hd__inv_2
XFILLER_0_101_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_208_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_184_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_160_4324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_4335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_199_5268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_4346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18763_ _06045_ _06112_ _05706_ VGND VGND VPWR VPWR _06113_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_199_5279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15975_ net2053 _13220_ _14322_ VGND VGND VPWR VPWR _14325_ sky130_fd_sc_hd__mux2_1
X_17714_ _13220_ net3851 _05129_ VGND VGND VPWR VPWR _05132_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14926_ _13314_ VGND VGND VPWR VPWR _13475_ sky130_fd_sc_hd__clkbuf_4
X_18694_ _05872_ _06047_ _05697_ VGND VGND VPWR VPWR _06048_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30972_ clknet_leaf_201_clk _02707_ VGND VGND VPWR VPWR datamem.data_ram\[39\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32711_ clknet_leaf_86_clk _04133_ VGND VGND VPWR VPWR datamem.data_ram\[17\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17645_ _05095_ VGND VGND VPWR VPWR _01216_ sky130_fd_sc_hd__clkbuf_1
X_14857_ _13408_ VGND VGND VPWR VPWR _13409_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_63_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_63_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32642_ clknet_leaf_156_clk _04064_ VGND VGND VPWR VPWR datamem.data_ram\[1\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14788_ _13340_ VGND VGND VPWR VPWR _13341_ sky130_fd_sc_hd__clkbuf_4
X_17576_ _13217_ net3770 _05057_ VGND VGND VPWR VPWR _05059_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_158_4286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_4297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19315_ _06610_ VGND VGND VPWR VPWR _06611_ sky130_fd_sc_hd__buf_8
X_16527_ _04501_ VGND VGND VPWR VPWR _01780_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32573_ clknet_leaf_287_clk _03995_ VGND VGND VPWR VPWR datamem.data_ram\[22\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31524_ clknet_leaf_45_clk net1210 VGND VGND VPWR VPWR rvcpu.dp.plem.PCPlus4M\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_19246_ _06548_ _06549_ VGND VGND VPWR VPWR _06550_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16458_ _14273_ VGND VGND VPWR VPWR _04464_ sky130_fd_sc_hd__inv_2
XFILLER_0_156_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15409_ _13665_ _13348_ _13940_ VGND VGND VPWR VPWR _13941_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_22_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19177_ _06488_ _06489_ VGND VGND VPWR VPWR _06490_ sky130_fd_sc_hd__nand2_1
X_31455_ clknet_leaf_5_clk rvcpu.dp.SrcBFW_Mux.y\[13\] VGND VGND VPWR VPWR rvcpu.dp.plem.WriteDataM\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16389_ _14559_ VGND VGND VPWR VPWR _01844_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18128_ _05490_ _05493_ VGND VGND VPWR VPWR _05494_ sky130_fd_sc_hd__nand2_1
X_30406_ net744 _02141_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[31\]\[17\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_93_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31386_ clknet_leaf_32_clk _03089_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCE\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23887__447 clknet_1_1__leaf__10222_ VGND VGND VPWR VPWR net573 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_93_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18059_ _05425_ _05426_ VGND VGND VPWR VPWR _05427_ sky130_fd_sc_hd__nor2_1
X_24106__614 clknet_1_0__leaf__10258_ VGND VGND VPWR VPWR net740 sky130_fd_sc_hd__inv_2
X_30337_ net683 _02072_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[4\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21070_ _07866_ _08357_ _08358_ VGND VGND VPWR VPWR _08359_ sky130_fd_sc_hd__and3_1
XFILLER_0_112_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30268_ net622 _02003_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[6\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20021_ datamem.data_ram\[46\]\[2\] _06950_ _06953_ datamem.data_ram\[44\]\[2\] VGND
+ VGND VPWR VPWR _07315_ sky130_fd_sc_hd__a22o_1
X_32007_ clknet_leaf_127_clk _03429_ VGND VGND VPWR VPWR datamem.data_ram\[27\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_171_Right_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_3518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30199_ net553 _01934_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[8\]\[18\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_126_3529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_193_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24760_ _10465_ net3227 _10589_ VGND VGND VPWR VPWR _10590_ sky130_fd_sc_hd__mux2_1
XFILLER_0_213_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21972_ rvcpu.dp.rf.reg_file_arr\[4\]\[31\] rvcpu.dp.rf.reg_file_arr\[5\]\[31\] rvcpu.dp.rf.reg_file_arr\[6\]\[31\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[31\] _08696_ _08825_ VGND VGND VPWR VPWR _09203_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_83_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_174_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23711_ clknet_1_0__leaf__10192_ VGND VGND VPWR VPWR _10197_ sky130_fd_sc_hd__buf_1
X_20923_ datamem.data_ram\[42\]\[22\] datamem.data_ram\[43\]\[22\] _07827_ VGND VGND
+ VPWR VPWR _08213_ sky130_fd_sc_hd__mux2_1
X_32909_ clknet_leaf_262_clk _04331_ VGND VGND VPWR VPWR datamem.data_ram\[7\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24691_ _10439_ net4147 _10552_ VGND VGND VPWR VPWR _10553_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26430_ _06461_ _11522_ VGND VGND VPWR VPWR _11564_ sky130_fd_sc_hd__and2_1
XFILLER_0_178_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23642_ _10187_ VGND VGND VPWR VPWR _01744_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20854_ _06680_ _06595_ VGND VGND VPWR VPWR _08144_ sky130_fd_sc_hd__nand2_8
XFILLER_0_193_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26361_ _11501_ net1445 _11510_ _11514_ VGND VGND VPWR VPWR _03136_ sky130_fd_sc_hd__a31o_1
XFILLER_0_3_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20785_ datamem.data_ram\[17\]\[30\] _07832_ VGND VGND VPWR VPWR _08075_ sky130_fd_sc_hd__or2_1
X_28100_ _12456_ net3307 net75 VGND VGND VPWR VPWR _12515_ sky130_fd_sc_hd__mux2_1
X_25312_ _10814_ net2803 _10899_ VGND VGND VPWR VPWR _10901_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29080_ _13054_ VGND VGND VPWR VPWR _04315_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22524_ _09441_ _09678_ VGND VGND VPWR VPWR _09679_ sky130_fd_sc_hd__nor2_1
X_26292_ net1291 _11478_ VGND VGND VPWR VPWR _11479_ sky130_fd_sc_hd__and2_1
XFILLER_0_91_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_487 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28031_ _12439_ net4436 _12473_ VGND VGND VPWR VPWR _12478_ sky130_fd_sc_hd__mux2_1
X_25243_ _10861_ VGND VGND VPWR VPWR _02671_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22455_ _09613_ VGND VGND VPWR VPWR _01131_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_59_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21406_ _08542_ _08665_ VGND VGND VPWR VPWR _08666_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_59_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25174_ _10822_ net3919 net58 VGND VGND VPWR VPWR _10823_ sky130_fd_sc_hd__mux2_1
XFILLER_0_228_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22386_ rvcpu.dp.rf.reg_file_arr\[4\]\[4\] rvcpu.dp.rf.reg_file_arr\[5\]\[4\] rvcpu.dp.rf.reg_file_arr\[6\]\[4\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[4\] _09423_ _09424_ VGND VGND VPWR VPWR _09548_ sky130_fd_sc_hd__mux4_1
X_23946__500 clknet_1_1__leaf__10228_ VGND VGND VPWR VPWR net626 sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_284_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_284_clk
+ sky130_fd_sc_hd__clkbuf_8
X_21337_ rvcpu.ALUResultE\[23\] _06294_ _06305_ rvcpu.ALUResultE\[29\] VGND VGND VPWR
+ VPWR _08599_ sky130_fd_sc_hd__or4_1
XFILLER_0_20_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29982_ net352 _01717_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[14\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_202_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28933_ _12972_ VGND VGND VPWR VPWR _04250_ sky130_fd_sc_hd__clkbuf_1
Xhold570 rvcpu.dp.plfd.PCD\[19\] VGND VGND VPWR VPWR net1720 sky130_fd_sc_hd__dlygate4sd3_1
X_21268_ _08523_ _08529_ VGND VGND VPWR VPWR _08530_ sky130_fd_sc_hd__nor2_1
Xhold581 datamem.data_ram\[15\]\[1\] VGND VGND VPWR VPWR net1731 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_229_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold592 rvcpu.dp.plem.ALUResultM\[2\] VGND VGND VPWR VPWR net1742 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20219_ datamem.data_ram\[26\]\[3\] _07136_ _07508_ _07511_ VGND VGND VPWR VPWR _07512_
+ sky130_fd_sc_hd__a211o_1
X_28864_ _12694_ net3716 _12932_ VGND VGND VPWR VPWR _12936_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21199_ _08481_ VGND VGND VPWR VPWR _04418_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_202_5342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27815_ _12350_ VGND VGND VPWR VPWR _03754_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_202_5353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28795_ _12899_ VGND VGND VPWR VPWR _04185_ sky130_fd_sc_hd__clkbuf_1
X_15760_ _14149_ net2767 _14199_ VGND VGND VPWR VPWR _14209_ sky130_fd_sc_hd__mux2_1
X_27746_ _12312_ VGND VGND VPWR VPWR _03723_ sky130_fd_sc_hd__clkbuf_1
X_24958_ _10698_ VGND VGND VPWR VPWR _02549_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_216_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1270 datamem.data_ram\[38\]\[25\] VGND VGND VPWR VPWR net2420 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_194_5143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_194_5154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14711_ rvcpu.dp.plmw.ALUResultW\[3\] rvcpu.dp.plmw.ReadDataW\[3\] rvcpu.dp.plmw.PCPlus4W\[3\]
+ rvcpu.dp.plmw.lAuiPCW\[3\] rvcpu.dp.plmw.ResultSrcW\[0\] rvcpu.dp.plmw.ResultSrcW\[1\]
+ VGND VGND VPWR VPWR _13268_ sky130_fd_sc_hd__mux4_2
Xhold1281 rvcpu.dp.rf.reg_file_arr\[27\]\[3\] VGND VGND VPWR VPWR net2431 sky130_fd_sc_hd__dlygate4sd3_1
X_15691_ _14164_ net2833 _14152_ VGND VGND VPWR VPWR _14165_ sky130_fd_sc_hd__mux2_1
Xhold1292 datamem.data_ram\[58\]\[30\] VGND VGND VPWR VPWR net2442 sky130_fd_sc_hd__dlygate4sd3_1
X_24889_ _10661_ VGND VGND VPWR VPWR _02517_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_410 _06647_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27677_ _12275_ VGND VGND VPWR VPWR _03691_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_212_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_421 _06776_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_213_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14642_ rvcpu.dp.plmw.ALUResultW\[20\] rvcpu.dp.plmw.ReadDataW\[20\] rvcpu.dp.plmw.PCPlus4W\[20\]
+ rvcpu.dp.plmw.lAuiPCW\[20\] _13169_ _13171_ VGND VGND VPWR VPWR _13216_ sky130_fd_sc_hd__mux4_2
XFILLER_0_157_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29416_ clknet_leaf_12_clk _01151_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD2E\[27\] sky130_fd_sc_hd__dfxtp_1
X_17430_ _04981_ VGND VGND VPWR VPWR _01325_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_432 _06815_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26628_ _10782_ _11659_ _11660_ net1349 VGND VGND VPWR VPWR _03257_ sky130_fd_sc_hd__a22o_1
XFILLER_0_185_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_443 _07023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_454 _08125_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_465 _08744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_476 _09317_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_0__10228_ _10228_ VGND VGND VPWR VPWR clknet_0__10228_ sky130_fd_sc_hd__clkbuf_16
XANTENNA_487 _09478_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17361_ _14143_ net4219 _04938_ VGND VGND VPWR VPWR _04945_ sky130_fd_sc_hd__mux2_1
X_29347_ clknet_leaf_196_clk _01082_ VGND VGND VPWR VPWR datamem.data_ram\[61\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__10128_ clknet_0__10128_ VGND VGND VPWR VPWR clknet_1_1__leaf__10128_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_498 _11078_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26559_ _11624_ VGND VGND VPWR VPWR _03224_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19100_ rvcpu.dp.plde.ImmExtE\[11\] rvcpu.dp.plde.PCE\[11\] VGND VGND VPWR VPWR _06422_
+ sky130_fd_sc_hd__nand2_1
X_16312_ net4028 _14478_ _14511_ VGND VGND VPWR VPWR _14519_ sky130_fd_sc_hd__mux2_1
X_17292_ _04908_ VGND VGND VPWR VPWR _01398_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__10159_ _10159_ VGND VGND VPWR VPWR clknet_0__10159_ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_153_4161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29278_ _13160_ VGND VGND VPWR VPWR _04407_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_193_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_153_4172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19031_ _06360_ _06361_ VGND VGND VPWR VPWR _06362_ sky130_fd_sc_hd__nand2_1
X_16243_ net1967 _14480_ _14464_ VGND VGND VPWR VPWR _14481_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28229_ _12430_ net3084 _12583_ VGND VGND VPWR VPWR _12584_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_563 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23378__1013 clknet_1_1__leaf__10139_ VGND VGND VPWR VPWR net1139 sky130_fd_sc_hd__inv_2
X_31240_ clknet_leaf_35_clk _02943_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCD\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_207_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16174_ _13200_ VGND VGND VPWR VPWR _14434_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_209_5507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_209_5518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15125_ _13664_ _13667_ _13669_ VGND VGND VPWR VPWR _13670_ sky130_fd_sc_hd__or3b_1
Xclkbuf_leaf_275_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_275_clk
+ sky130_fd_sc_hd__clkbuf_8
X_31171_ clknet_leaf_13_clk rvcpu.ALUResultE\[30\] VGND VGND VPWR VPWR rvcpu.dp.plem.ALUResultM\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30122_ net484 _01857_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[10\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_15056_ _13291_ _13578_ VGND VGND VPWR VPWR _13603_ sky130_fd_sc_hd__nand2_1
X_19933_ _07153_ _07179_ _07226_ _07227_ VGND VGND VPWR VPWR _07228_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_112_3190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_183_4880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30053_ net415 _01788_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[12\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19864_ _06978_ VGND VGND VPWR VPWR _07159_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_183_4891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18815_ _05504_ _05727_ _06161_ VGND VGND VPWR VPWR _06162_ sky130_fd_sc_hd__a21oi_1
X_19795_ datamem.data_ram\[62\]\[9\] _06629_ _06620_ datamem.data_ram\[60\]\[9\] VGND
+ VGND VPWR VPWR _07090_ sky130_fd_sc_hd__o22a_1
X_18746_ _05693_ _05805_ _05935_ VGND VGND VPWR VPWR _06097_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_121_3404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15958_ net2836 _13195_ _14311_ VGND VGND VPWR VPWR _14316_ sky130_fd_sc_hd__mux2_1
X_14909_ _13291_ _13304_ VGND VGND VPWR VPWR _13459_ sky130_fd_sc_hd__nor2_1
XFILLER_0_204_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18677_ _06031_ _05865_ _05820_ VGND VGND VPWR VPWR _06032_ sky130_fd_sc_hd__o21a_1
X_30955_ clknet_leaf_277_clk _02690_ VGND VGND VPWR VPWR datamem.data_ram\[3\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15889_ _14279_ VGND VGND VPWR VPWR _02080_ sky130_fd_sc_hd__clkbuf_1
X_17628_ _05086_ VGND VGND VPWR VPWR _01224_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_176_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_82_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30886_ clknet_leaf_222_clk _02621_ VGND VGND VPWR VPWR datamem.data_ram\[42\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_82_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32625_ clknet_leaf_93_clk _04047_ VGND VGND VPWR VPWR datamem.data_ram\[1\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_176_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_175_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17559_ _13190_ net4241 _05046_ VGND VGND VPWR VPWR _05050_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_1278 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_3355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32556_ clknet_leaf_233_clk _03978_ VGND VGND VPWR VPWR datamem.data_ram\[22\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20570_ datamem.data_ram\[38\]\[13\] datamem.data_ram\[39\]\[13\] _07829_ VGND VGND
+ VPWR VPWR _07861_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31507_ clknet_leaf_66_clk net1288 VGND VGND VPWR VPWR rvcpu.dp.plem.PCPlus4M\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_19229_ rvcpu.dp.plde.ImmExtE\[27\] rvcpu.dp.plde.PCE\[27\] VGND VGND VPWR VPWR _06535_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_144_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32487_ clknet_leaf_186_clk _03909_ VGND VGND VPWR VPWR datamem.data_ram\[25\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_574 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22240_ _08592_ VGND VGND VPWR VPWR _09406_ sky130_fd_sc_hd__buf_6
XFILLER_0_5_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31438_ clknet_leaf_102_clk _03141_ VGND VGND VPWR VPWR datamem.data_ram\[14\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_266_clk clknet_5_19__leaf_clk VGND VGND VPWR VPWR clknet_leaf_266_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_147_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22171_ _09318_ net2732 _09352_ VGND VGND VPWR VPWR _09357_ sky130_fd_sc_hd__mux2_1
X_31369_ clknet_leaf_13_clk _03072_ VGND VGND VPWR VPWR rvcpu.dp.plde.ImmExtE\[18\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_2_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23136__812 clknet_1_0__leaf__10106_ VGND VGND VPWR VPWR net938 sky130_fd_sc_hd__inv_2
X_21122_ datamem.data_ram\[46\]\[23\] _07831_ _08410_ _07838_ VGND VGND VPWR VPWR
+ _08411_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_54_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25930_ net1326 _11279_ VGND VGND VPWR VPWR _11285_ sky130_fd_sc_hd__or2_1
X_21053_ _08340_ _08341_ _07819_ VGND VGND VPWR VPWR _08342_ sky130_fd_sc_hd__mux2_1
XFILLER_0_226_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__10079_ clknet_0__10079_ VGND VGND VPWR VPWR clknet_1_0__leaf__10079_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_185_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20004_ _06714_ _07292_ _07297_ _06594_ VGND VGND VPWR VPWR _07298_ sky130_fd_sc_hd__a31o_1
X_25861_ _11239_ _11240_ VGND VGND VPWR VPWR _11241_ sky130_fd_sc_hd__nor2_1
XFILLER_0_199_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24812_ _10619_ VGND VGND VPWR VPWR _02482_ sky130_fd_sc_hd__clkbuf_1
X_27600_ _12234_ VGND VGND VPWR VPWR _03655_ sky130_fd_sc_hd__clkbuf_1
X_25792_ rvcpu.dp.pcreg.q\[14\] _11182_ VGND VGND VPWR VPWR _11186_ sky130_fd_sc_hd__or2_1
X_28580_ _12784_ VGND VGND VPWR VPWR _04085_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_213_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27531_ _12125_ net2821 _12197_ VGND VGND VPWR VPWR _12198_ sky130_fd_sc_hd__mux2_1
X_24743_ _10385_ net2960 _10580_ VGND VGND VPWR VPWR _10581_ sky130_fd_sc_hd__mux2_1
X_21955_ rvcpu.dp.rf.reg_file_arr\[4\]\[30\] rvcpu.dp.rf.reg_file_arr\[5\]\[30\] rvcpu.dp.rf.reg_file_arr\[6\]\[30\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[30\] _08628_ _08856_ VGND VGND VPWR VPWR _09187_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_68_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_210_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20906_ datamem.data_ram\[8\]\[22\] _07191_ _08191_ _08195_ VGND VGND VPWR VPWR _08196_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_139_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27462_ _12160_ VGND VGND VPWR VPWR _03591_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_48_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24674_ _10385_ net2813 _10543_ VGND VGND VPWR VPWR _10544_ sky130_fd_sc_hd__mux2_1
X_21886_ rvcpu.dp.rf.reg_file_arr\[4\]\[26\] rvcpu.dp.rf.reg_file_arr\[5\]\[26\] rvcpu.dp.rf.reg_file_arr\[6\]\[26\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[26\] _08839_ _08840_ VGND VGND VPWR VPWR _09122_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_49_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29201_ _13118_ VGND VGND VPWR VPWR _04372_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_104_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26413_ _11524_ rvcpu.ALUResultE\[10\] _11173_ _11526_ VGND VGND VPWR VPWR _11553_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_178_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20837_ _07635_ datamem.data_ram\[30\]\[14\] VGND VGND VPWR VPWR _08127_ sky130_fd_sc_hd__or2_1
X_27393_ _10668_ _10898_ _11713_ VGND VGND VPWR VPWR _12116_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_166_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26344_ _10780_ _11507_ VGND VGND VPWR VPWR _11508_ sky130_fd_sc_hd__nor2_2
X_29132_ _09251_ net2017 _13076_ VGND VGND VPWR VPWR _13082_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20768_ _08054_ _08055_ _08056_ _08057_ VGND VGND VPWR VPWR _08058_ sky130_fd_sc_hd__or4_1
XFILLER_0_181_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23223__873 clknet_1_0__leaf__10124_ VGND VGND VPWR VPWR net999 sky130_fd_sc_hd__inv_2
XFILLER_0_181_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22507_ rvcpu.dp.rf.reg_file_arr\[12\]\[10\] rvcpu.dp.rf.reg_file_arr\[13\]\[10\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[10\] rvcpu.dp.rf.reg_file_arr\[15\]\[10\] _09386_
+ _09467_ VGND VGND VPWR VPWR _09663_ sky130_fd_sc_hd__mux4_2
X_29063_ _13045_ VGND VGND VPWR VPWR _04307_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26275_ net1627 _11467_ VGND VGND VPWR VPWR _11470_ sky130_fd_sc_hd__and2_1
XFILLER_0_107_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20699_ datamem.data_ram\[0\]\[5\] _06937_ _06961_ datamem.data_ram\[3\]\[5\] _06742_
+ VGND VGND VPWR VPWR _07990_ sky130_fd_sc_hd__a221o_1
XFILLER_0_107_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25226_ _10852_ VGND VGND VPWR VPWR _02663_ sky130_fd_sc_hd__clkbuf_1
X_28014_ _12365_ net4264 net97 VGND VGND VPWR VPWR _12469_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22438_ rvcpu.dp.rf.reg_file_arr\[28\]\[7\] rvcpu.dp.rf.reg_file_arr\[30\]\[7\] rvcpu.dp.rf.reg_file_arr\[29\]\[7\]
+ rvcpu.dp.rf.reg_file_arr\[31\]\[7\] _09446_ _09402_ VGND VGND VPWR VPWR _09597_
+ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_257_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_257_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_165_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25157_ _09297_ VGND VGND VPWR VPWR _10811_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_0_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22369_ _09385_ VGND VGND VPWR VPWR _09532_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_206_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25088_ _10775_ VGND VGND VPWR VPWR _02602_ sky130_fd_sc_hd__clkbuf_1
X_29965_ net335 _01700_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[15\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28916_ _12963_ VGND VGND VPWR VPWR _04242_ sky130_fd_sc_hd__clkbuf_1
X_16930_ _04715_ VGND VGND VPWR VPWR _01575_ sky130_fd_sc_hd__clkbuf_1
X_29896_ net274 _01631_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[17\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_196_5205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16861_ net2499 _14480_ _04670_ VGND VGND VPWR VPWR _04679_ sky130_fd_sc_hd__mux2_1
X_28847_ _12741_ net4184 net69 VGND VGND VPWR VPWR _12927_ sky130_fd_sc_hd__mux2_1
X_18600_ _05957_ _05592_ _05933_ VGND VGND VPWR VPWR _05958_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_221_5795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15812_ _14237_ VGND VGND VPWR VPWR _02115_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_217_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19580_ datamem.data_ram\[32\]\[8\] _06821_ _06618_ datamem.data_ram\[36\]\[8\] VGND
+ VGND VPWR VPWR _06876_ sky130_fd_sc_hd__o22a_1
X_28778_ _12890_ VGND VGND VPWR VPWR _04177_ sky130_fd_sc_hd__clkbuf_1
X_16792_ _04642_ VGND VGND VPWR VPWR _01648_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_176_1294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18531_ _05603_ _05565_ _05566_ _05570_ _05668_ _05663_ VGND VGND VPWR VPWR _05892_
+ sky130_fd_sc_hd__mux4_1
X_15743_ _14200_ VGND VGND VPWR VPWR _02155_ sky130_fd_sc_hd__clkbuf_1
X_27729_ _12303_ VGND VGND VPWR VPWR _03715_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_198_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24135__640 clknet_1_1__leaf__10261_ VGND VGND VPWR VPWR net766 sky130_fd_sc_hd__inv_2
XFILLER_0_169_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18462_ _05643_ _05636_ _05637_ _05632_ _05682_ _05579_ VGND VGND VPWR VPWR _05825_
+ sky130_fd_sc_hd__mux4_1
X_30740_ clknet_leaf_200_clk _02475_ VGND VGND VPWR VPWR datamem.data_ram\[47\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_240 _11047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23541__166 clknet_1_1__leaf__10173_ VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__inv_2
X_15674_ _14153_ VGND VGND VPWR VPWR _02177_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_155_4212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_4223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_251 _13195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_201_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17413_ _14195_ net2699 _04937_ VGND VGND VPWR VPWR _04972_ sky130_fd_sc_hd__mux2_1
XANTENNA_262 _13216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14625_ rvcpu.dp.plmw.ALUResultW\[24\] rvcpu.dp.plmw.ReadDataW\[24\] rvcpu.dp.plmw.PCPlus4W\[24\]
+ rvcpu.dp.plmw.lAuiPCW\[24\] _13192_ _13193_ VGND VGND VPWR VPWR _13203_ sky130_fd_sc_hd__mux4_2
XFILLER_0_158_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_273 _13235_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18393_ _05286_ _05662_ VGND VGND VPWR VPWR _05757_ sky130_fd_sc_hd__nor2_1
XANTENNA_284 _13266_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30671_ clknet_leaf_178_clk _02406_ VGND VGND VPWR VPWR datamem.data_ram\[50\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_295 _13588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_4109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32410_ clknet_leaf_238_clk _03832_ VGND VGND VPWR VPWR datamem.data_ram\[28\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_17344_ _04935_ VGND VGND VPWR VPWR _01373_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_184_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32341_ clknet_leaf_246_clk _03763_ VGND VGND VPWR VPWR datamem.data_ram\[30\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17275_ _04898_ VGND VGND VPWR VPWR _01405_ sky130_fd_sc_hd__clkbuf_1
X_19014_ _05707_ _06282_ _06347_ VGND VGND VPWR VPWR _06348_ sky130_fd_sc_hd__o21a_1
XFILLER_0_10_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload204 clknet_leaf_198_clk VGND VGND VPWR VPWR clkload204/Y sky130_fd_sc_hd__bufinv_16
Xclkload215 clknet_leaf_166_clk VGND VGND VPWR VPWR clkload215/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_114_3230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16226_ _14469_ VGND VGND VPWR VPWR _01925_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_183_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_114_3241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32272_ clknet_leaf_201_clk _03694_ VGND VGND VPWR VPWR datamem.data_ram\[33\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload226 clknet_leaf_165_clk VGND VGND VPWR VPWR clkload226/Y sky130_fd_sc_hd__bufinv_16
Xclkload237 clknet_leaf_117_clk VGND VGND VPWR VPWR clkload237/Y sky130_fd_sc_hd__clkinv_1
Xclkload248 clknet_leaf_151_clk VGND VGND VPWR VPWR clkload248/Y sky130_fd_sc_hd__inv_8
XFILLER_0_113_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_248_clk clknet_5_17__leaf_clk VGND VGND VPWR VPWR clknet_leaf_248_clk
+ sky130_fd_sc_hd__clkbuf_8
X_31223_ clknet_leaf_39_clk _02926_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCD\[12\] sky130_fd_sc_hd__dfxtp_1
Xclkload259 clknet_leaf_146_clk VGND VGND VPWR VPWR clkload259/Y sky130_fd_sc_hd__inv_6
X_16157_ net3331 _14420_ _14422_ VGND VGND VPWR VPWR _14423_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_185_4931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_185_4942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_110_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15108_ _13392_ _13523_ _13536_ VGND VGND VPWR VPWR _13653_ sky130_fd_sc_hd__a21o_1
X_31154_ clknet_leaf_69_clk rvcpu.ALUResultE\[13\] VGND VGND VPWR VPWR rvcpu.dp.plem.ALUResultM\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16088_ net3489 _13173_ _14385_ VGND VGND VPWR VPWR _14386_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_181_4828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15039_ _13282_ _13415_ VGND VGND VPWR VPWR _13586_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_181_4839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19916_ datamem.data_ram\[34\]\[17\] _06612_ _06863_ datamem.data_ram\[35\]\[17\]
+ _06776_ VGND VGND VPWR VPWR _07211_ sky130_fd_sc_hd__o221a_1
XFILLER_0_139_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30105_ net467 _01840_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[11\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_31085_ clknet_leaf_101_clk _02820_ VGND VGND VPWR VPWR datamem.data_ram\[21\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2707 rvcpu.dp.rf.reg_file_arr\[28\]\[29\] VGND VGND VPWR VPWR net3857 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2718 rvcpu.dp.rf.reg_file_arr\[17\]\[22\] VGND VGND VPWR VPWR net3868 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_71_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2729 rvcpu.dp.rf.reg_file_arr\[27\]\[16\] VGND VGND VPWR VPWR net3879 sky130_fd_sc_hd__dlygate4sd3_1
X_30036_ net398 _01771_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[13\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_19847_ datamem.data_ram\[54\]\[1\] _06952_ _06969_ datamem.data_ram\[53\]\[1\] VGND
+ VGND VPWR VPWR _07142_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_144_3960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19778_ datamem.data_ram\[39\]\[9\] _06761_ _06700_ datamem.data_ram\[33\]\[9\] VGND
+ VGND VPWR VPWR _07073_ sky130_fd_sc_hd__o22a_1
XFILLER_0_74_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18729_ _05436_ VGND VGND VPWR VPWR _06081_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_140_3846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31987_ clknet_leaf_117_clk _03409_ VGND VGND VPWR VPWR datamem.data_ram\[37\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23166__838 clknet_1_1__leaf__10110_ VGND VGND VPWR VPWR net964 sky130_fd_sc_hd__inv_2
X_23704__298 clknet_1_0__leaf__10196_ VGND VGND VPWR VPWR net424 sky130_fd_sc_hd__inv_2
X_21740_ _08842_ _08983_ VGND VGND VPWR VPWR _08984_ sky130_fd_sc_hd__or2_1
XFILLER_0_149_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30938_ clknet_leaf_181_clk _02673_ VGND VGND VPWR VPWR datamem.data_ram\[40\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
Xwire78 _12346_ VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__buf_4
XFILLER_0_171_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21671_ _08514_ _08917_ VGND VGND VPWR VPWR _08918_ sky130_fd_sc_hd__or2_1
X_30869_ clknet_leaf_64_clk _02604_ VGND VGND VPWR VPWR datamem.data_ram\[42\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23410_ clknet_1_0__leaf__10078_ VGND VGND VPWR VPWR _10152_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_43_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32608_ clknet_leaf_183_clk _04030_ VGND VGND VPWR VPWR datamem.data_ram\[20\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_20622_ datamem.data_ram\[14\]\[13\] _07912_ VGND VGND VPWR VPWR _07913_ sky130_fd_sc_hd__or2_1
X_24390_ _09256_ net4379 _10367_ VGND VGND VPWR VPWR _10374_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32539_ clknet_leaf_78_clk _03961_ VGND VGND VPWR VPWR datamem.data_ram\[23\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20553_ _06614_ VGND VGND VPWR VPWR _07844_ sky130_fd_sc_hd__buf_6
XFILLER_0_85_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_580 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26060_ _11091_ _11351_ VGND VGND VPWR VPWR _11359_ sky130_fd_sc_hd__and2_1
XFILLER_0_144_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_229_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20484_ datamem.data_ram\[56\]\[20\] _06820_ _06617_ datamem.data_ram\[60\]\[20\]
+ _07775_ VGND VGND VPWR VPWR _07776_ sky130_fd_sc_hd__o221a_1
XFILLER_0_15_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25011_ _10727_ net2239 _10725_ VGND VGND VPWR VPWR _10728_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_239_clk clknet_5_17__leaf_clk VGND VGND VPWR VPWR clknet_leaf_239_clk
+ sky130_fd_sc_hd__clkbuf_8
X_22223_ _09388_ VGND VGND VPWR VPWR _09389_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_120_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22154_ _09285_ net2983 net62 VGND VGND VPWR VPWR _09347_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21105_ _08382_ _08386_ _06860_ _08393_ VGND VGND VPWR VPWR _08394_ sky130_fd_sc_hd__o211a_1
X_29750_ net1096 _01485_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[21\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_26962_ _11752_ VGND VGND VPWR VPWR _11863_ sky130_fd_sc_hd__clkbuf_4
X_22085_ _07132_ VGND VGND VPWR VPWR _09299_ sky130_fd_sc_hd__buf_6
Xfanout121 _00000_ VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__buf_1
X_24004__537 clknet_1_0__leaf__10241_ VGND VGND VPWR VPWR net663 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_7_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28701_ _12749_ net4102 net42 VGND VGND VPWR VPWR _12849_ sky130_fd_sc_hd__mux2_1
X_25913_ net1821 _11263_ VGND VGND VPWR VPWR _11276_ sky130_fd_sc_hd__or2_1
X_21036_ _06851_ _08317_ _08324_ _07176_ VGND VGND VPWR VPWR _08325_ sky130_fd_sc_hd__a211o_1
X_29681_ net1027 _01416_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[23\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26893_ _11672_ _11810_ VGND VGND VPWR VPWR _11819_ sky130_fd_sc_hd__and2_1
XFILLER_0_227_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28632_ _12812_ VGND VGND VPWR VPWR _04109_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25844_ rvcpu.dp.pcreg.q\[25\] _11221_ VGND VGND VPWR VPWR _11227_ sky130_fd_sc_hd__nor2_1
X_23377__1012 clknet_1_1__leaf__10139_ VGND VGND VPWR VPWR net1138 sky130_fd_sc_hd__inv_2
XFILLER_0_214_567 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28563_ _12775_ VGND VGND VPWR VPWR _04077_ sky130_fd_sc_hd__clkbuf_1
X_25775_ _11171_ _11172_ _11149_ VGND VGND VPWR VPWR _11173_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_214_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27514_ _12080_ net3476 net99 VGND VGND VPWR VPWR _12189_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24726_ _10439_ net3611 _10571_ VGND VGND VPWR VPWR _10572_ sky130_fd_sc_hd__mux2_1
X_21938_ rvcpu.dp.rf.reg_file_arr\[0\]\[29\] rvcpu.dp.rf.reg_file_arr\[1\]\[29\] rvcpu.dp.rf.reg_file_arr\[2\]\[29\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[29\] _08525_ _08528_ VGND VGND VPWR VPWR _09171_
+ sky130_fd_sc_hd__mux4_1
X_28494_ _12727_ net1498 _12723_ _12731_ VGND VGND VPWR VPWR _04052_ sky130_fd_sc_hd__a31o_1
XFILLER_0_195_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23679__275 clknet_1_0__leaf__10194_ VGND VGND VPWR VPWR net401 sky130_fd_sc_hd__inv_2
X_24657_ _10408_ _10532_ VGND VGND VPWR VPWR _10534_ sky130_fd_sc_hd__and2_1
X_27445_ _09278_ VGND VGND VPWR VPWR _12149_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_78_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21869_ rvcpu.dp.rf.reg_file_arr\[0\]\[25\] rvcpu.dp.rf.reg_file_arr\[1\]\[25\] rvcpu.dp.rf.reg_file_arr\[2\]\[25\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[25\] _08550_ _08554_ VGND VGND VPWR VPWR _09106_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_194_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15390_ _13298_ _13374_ _13604_ _13635_ _13438_ VGND VGND VPWR VPWR _13923_ sky130_fd_sc_hd__o311a_1
XFILLER_0_182_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27376_ _10598_ _12106_ _11713_ VGND VGND VPWR VPWR _12107_ sky130_fd_sc_hd__a21oi_1
X_24588_ _10392_ net2940 _10491_ VGND VGND VPWR VPWR _10495_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_189_5020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_189_5031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29115_ _09284_ net3648 _13067_ VGND VGND VPWR VPWR _13073_ sky130_fd_sc_hd__mux2_1
X_26327_ _11353_ net1806 _11496_ _11498_ VGND VGND VPWR VPWR _03118_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_189_5042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23539_ clknet_1_0__leaf__10172_ VGND VGND VPWR VPWR _10173_ sky130_fd_sc_hd__buf_1
XFILLER_0_52_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_1308 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17060_ net2814 _14474_ _04779_ VGND VGND VPWR VPWR _04785_ sky130_fd_sc_hd__mux2_1
X_29046_ _13018_ net1636 _13030_ _13036_ VGND VGND VPWR VPWR _04299_ sky130_fd_sc_hd__a31o_1
XFILLER_0_208_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26258_ net1377 _11432_ VGND VGND VPWR VPWR _11461_ sky130_fd_sc_hd__and2_1
XFILLER_0_122_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16011_ _14343_ VGND VGND VPWR VPWR _02022_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_208_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25209_ _10843_ VGND VGND VPWR VPWR _02655_ sky130_fd_sc_hd__clkbuf_1
X_26189_ _11431_ VGND VGND VPWR VPWR _03047_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_223_5846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17962_ _05325_ _05331_ _05332_ VGND VGND VPWR VPWR _05333_ sky130_fd_sc_hd__a21o_1
X_29948_ net318 _01683_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[15\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_223_5857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19701_ _06949_ VGND VGND VPWR VPWR _06997_ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_29_Left_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16913_ net2889 _14463_ _04706_ VGND VGND VPWR VPWR _04707_ sky130_fd_sc_hd__mux2_1
XFILLER_0_224_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17893_ _05265_ VGND VGND VPWR VPWR _05266_ sky130_fd_sc_hd__buf_4
X_29879_ net257 _01614_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[17\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23924__480 clknet_1_1__leaf__10226_ VGND VGND VPWR VPWR net606 sky130_fd_sc_hd__inv_2
X_19632_ _06622_ _06640_ VGND VGND VPWR VPWR _06928_ sky130_fd_sc_hd__nand2_4
X_31910_ _04421_ net118 VGND VGND VPWR VPWR datamem.rd_data_mem\[15\] sky130_fd_sc_hd__dlxtn_1
XFILLER_0_217_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16844_ _04647_ VGND VGND VPWR VPWR _04670_ sky130_fd_sc_hd__buf_4
X_32890_ clknet_leaf_158_clk _04312_ VGND VGND VPWR VPWR datamem.data_ram\[10\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31841_ clknet_leaf_165_clk _03295_ VGND VGND VPWR VPWR datamem.data_ram\[8\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_19563_ _06714_ _06853_ _06858_ VGND VGND VPWR VPWR _06859_ sky130_fd_sc_hd__or3_1
X_23623__241 clknet_1_1__leaf__10180_ VGND VGND VPWR VPWR net367 sky130_fd_sc_hd__inv_2
X_16775_ _04633_ VGND VGND VPWR VPWR _01656_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_189_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18514_ _05582_ _05654_ _05875_ VGND VGND VPWR VPWR _05876_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_17_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15726_ _14188_ VGND VGND VPWR VPWR _02160_ sky130_fd_sc_hd__clkbuf_1
X_19494_ _06789_ VGND VGND VPWR VPWR _06790_ sky130_fd_sc_hd__buf_8
XFILLER_0_125_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31772_ clknet_leaf_213_clk _03226_ VGND VGND VPWR VPWR datamem.data_ram\[1\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_24180__21 clknet_1_0__leaf__10265_ VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__inv_2
XFILLER_0_73_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18445_ _05236_ _05652_ rvcpu.dp.plde.ALUControlE\[1\] VGND VGND VPWR VPWR _05808_
+ sky130_fd_sc_hd__and3b_2
X_30723_ clknet_leaf_177_clk _02458_ VGND VGND VPWR VPWR datamem.data_ram\[49\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_15657_ _14141_ net3233 _14131_ VGND VGND VPWR VPWR _14142_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_174_4665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_1_Left_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_200_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_174_4676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_38_Left_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14608_ _13189_ VGND VGND VPWR VPWR _13190_ sky130_fd_sc_hd__buf_4
X_18376_ _05740_ VGND VGND VPWR VPWR rvcpu.ALUResultE\[31\] sky130_fd_sc_hd__buf_1
X_30654_ clknet_leaf_217_clk _02389_ VGND VGND VPWR VPWR datamem.data_ram\[50\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_15588_ _14101_ VGND VGND VPWR VPWR _02211_ sky130_fd_sc_hd__clkbuf_1
X_17327_ net4437 _13250_ _04924_ VGND VGND VPWR VPWR _04927_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30585_ clknet_leaf_178_clk _02320_ VGND VGND VPWR VPWR datamem.data_ram\[53\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_32324_ clknet_leaf_88_clk _03746_ VGND VGND VPWR VPWR datamem.data_ram\[31\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17258_ _14177_ net4047 _04887_ VGND VGND VPWR VPWR _04890_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_77_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_3683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16209_ net4257 _14457_ _14443_ VGND VGND VPWR VPWR _14458_ sky130_fd_sc_hd__mux2_1
X_32255_ clknet_leaf_86_clk _03677_ VGND VGND VPWR VPWR datamem.data_ram\[34\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_133_3694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17189_ _04853_ VGND VGND VPWR VPWR _01446_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31206_ clknet_leaf_27_clk _02909_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCPlus4D\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32186_ clknet_leaf_259_clk _03608_ VGND VGND VPWR VPWR datamem.data_ram\[37\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3205 datamem.data_ram\[62\]\[18\] VGND VGND VPWR VPWR net4355 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold3216 rvcpu.dp.rf.reg_file_arr\[25\]\[27\] VGND VGND VPWR VPWR net4366 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_47_Left_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_228_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold3227 rvcpu.dp.rf.reg_file_arr\[22\]\[4\] VGND VGND VPWR VPWR net4377 sky130_fd_sc_hd__dlygate4sd3_1
X_31137_ clknet_leaf_235_clk _02872_ VGND VGND VPWR VPWR datamem.data_ram\[4\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3238 datamem.data_ram\[53\]\[13\] VGND VGND VPWR VPWR net4388 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3249 datamem.data_ram\[60\]\[18\] VGND VGND VPWR VPWR net4399 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_36_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2504 datamem.data_ram\[21\]\[28\] VGND VGND VPWR VPWR net3654 sky130_fd_sc_hd__dlygate4sd3_1
X_23784__370 clknet_1_0__leaf__10204_ VGND VGND VPWR VPWR net496 sky130_fd_sc_hd__inv_2
Xhold2515 datamem.data_ram\[28\]\[26\] VGND VGND VPWR VPWR net3665 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_36_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2526 rvcpu.dp.rf.reg_file_arr\[26\]\[17\] VGND VGND VPWR VPWR net3676 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31068_ clknet_leaf_281_clk _02803_ VGND VGND VPWR VPWR datamem.data_ram\[8\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2537 rvcpu.dp.rf.reg_file_arr\[13\]\[30\] VGND VGND VPWR VPWR net3687 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1803 rvcpu.dp.rf.reg_file_arr\[25\]\[30\] VGND VGND VPWR VPWR net2953 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2548 datamem.data_ram\[23\]\[12\] VGND VGND VPWR VPWR net3698 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2559 datamem.data_ram\[26\]\[11\] VGND VGND VPWR VPWR net3709 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1814 datamem.data_ram\[13\]\[25\] VGND VGND VPWR VPWR net2964 sky130_fd_sc_hd__dlygate4sd3_1
X_22910_ _10043_ VGND VGND VPWR VPWR _10044_ sky130_fd_sc_hd__clkbuf_4
Xhold1825 datamem.data_ram\[11\]\[27\] VGND VGND VPWR VPWR net2975 sky130_fd_sc_hd__dlygate4sd3_1
X_30019_ net381 _01754_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[13\]\[6\] sky130_fd_sc_hd__dfxtp_1
Xhold1836 datamem.data_ram\[37\]\[27\] VGND VGND VPWR VPWR net2986 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1847 datamem.data_ram\[30\]\[10\] VGND VGND VPWR VPWR net2997 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1858 datamem.data_ram\[37\]\[18\] VGND VGND VPWR VPWR net3008 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1869 datamem.data_ram\[50\]\[9\] VGND VGND VPWR VPWR net3019 sky130_fd_sc_hd__dlygate4sd3_1
X_22841_ rvcpu.dp.rf.reg_file_arr\[4\]\[28\] rvcpu.dp.rf.reg_file_arr\[5\]\[28\] rvcpu.dp.rf.reg_file_arr\[6\]\[28\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[28\] _09386_ _09419_ VGND VGND VPWR VPWR _09979_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_190_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25560_ _11038_ VGND VGND VPWR VPWR _02811_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22772_ rvcpu.dp.rf.reg_file_arr\[8\]\[24\] rvcpu.dp.rf.reg_file_arr\[10\]\[24\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[24\] rvcpu.dp.rf.reg_file_arr\[11\]\[24\] _09483_
+ _09656_ VGND VGND VPWR VPWR _09914_ sky130_fd_sc_hd__mux4_1
XFILLER_0_151_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24511_ _10448_ datamem.data_ram\[52\]\[20\] _10440_ VGND VGND VPWR VPWR _10449_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21723_ _08547_ _08965_ _08967_ _08652_ VGND VGND VPWR VPWR _08968_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_56_Left_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25491_ _11000_ VGND VGND VPWR VPWR _02780_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_192_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27230_ _11978_ _12019_ VGND VGND VPWR VPWR _12027_ sky130_fd_sc_hd__and2_1
X_24442_ _10056_ net2036 _10404_ _10407_ VGND VGND VPWR VPWR _02324_ sky130_fd_sc_hd__a31o_1
XFILLER_0_137_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21654_ rvcpu.dp.rf.reg_file_arr\[28\]\[14\] rvcpu.dp.rf.reg_file_arr\[30\]\[14\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[14\] rvcpu.dp.rf.reg_file_arr\[31\]\[14\] _08533_
+ _08636_ VGND VGND VPWR VPWR _08902_ sky130_fd_sc_hd__mux4_1
XFILLER_0_163_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_191_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27161_ _11974_ net1520 _11983_ _11986_ VGND VGND VPWR VPWR _03464_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_62_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20605_ datamem.data_ram\[58\]\[13\] _06728_ _06686_ datamem.data_ram\[60\]\[13\]
+ VGND VGND VPWR VPWR _07896_ sky130_fd_sc_hd__o22a_1
X_24373_ _10364_ VGND VGND VPWR VPWR _02298_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_62_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21585_ _08835_ _08836_ VGND VGND VPWR VPWR _08837_ sky130_fd_sc_hd__or2_1
XFILLER_0_151_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26112_ _11391_ VGND VGND VPWR VPWR _03009_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_201_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27092_ _11938_ net2172 _11940_ _11942_ VGND VGND VPWR VPWR _03439_ sky130_fd_sc_hd__a31o_1
X_20536_ _07826_ VGND VGND VPWR VPWR _07827_ sky130_fd_sc_hd__buf_6
XFILLER_0_7_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26043_ _11121_ net1828 _11339_ _11348_ VGND VGND VPWR VPWR _02984_ sky130_fd_sc_hd__a31o_1
XFILLER_0_127_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23419__72 clknet_1_0__leaf__10153_ VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__inv_2
X_20467_ datamem.data_ram\[45\]\[20\] _06702_ _06619_ datamem.data_ram\[44\]\[20\]
+ VGND VGND VPWR VPWR _07759_ sky130_fd_sc_hd__o22a_1
XFILLER_0_28_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22206_ _09282_ net3606 _09371_ VGND VGND VPWR VPWR _09376_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_65_Left_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23335__974 clknet_1_0__leaf__10135_ VGND VGND VPWR VPWR net1100 sky130_fd_sc_hd__inv_2
X_20398_ _06712_ _07668_ _07679_ _07689_ _06796_ VGND VGND VPWR VPWR _07690_ sky130_fd_sc_hd__a32o_1
X_29802_ clknet_leaf_205_clk _01537_ VGND VGND VPWR VPWR datamem.data_ram\[59\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_22137_ _09252_ net4064 _09332_ VGND VGND VPWR VPWR _09338_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27994_ _12456_ net3803 net76 VGND VGND VPWR VPWR _12457_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29733_ net1079 _01468_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[21\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_23034__735 clknet_1_1__leaf__10089_ VGND VGND VPWR VPWR net861 sky130_fd_sc_hd__inv_2
X_26945_ _09351_ _11112_ _11609_ VGND VGND VPWR VPWR _11854_ sky130_fd_sc_hd__and3_1
X_22068_ _09284_ VGND VGND VPWR VPWR _09285_ sky130_fd_sc_hd__buf_2
X_21019_ datamem.data_ram\[55\]\[31\] _06667_ _08307_ _06676_ VGND VGND VPWR VPWR
+ _08308_ sky130_fd_sc_hd__o211a_1
X_29664_ net1010 _01399_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[24\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_26876_ _11808_ VGND VGND VPWR VPWR _11809_ sky130_fd_sc_hd__buf_2
X_14890_ _13312_ _13313_ VGND VGND VPWR VPWR _13441_ sky130_fd_sc_hd__or2_2
XFILLER_0_214_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23114__792 clknet_1_1__leaf__10104_ VGND VGND VPWR VPWR net918 sky130_fd_sc_hd__inv_2
X_28615_ _12803_ VGND VGND VPWR VPWR _04101_ sky130_fd_sc_hd__clkbuf_1
X_25827_ rvcpu.dp.pcreg.q\[22\] _11208_ VGND VGND VPWR VPWR _11213_ sky130_fd_sc_hd__and2_1
X_29595_ net949 _01330_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[26\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_28546_ _09259_ VGND VGND VPWR VPWR _12766_ sky130_fd_sc_hd__buf_2
X_16560_ _04519_ VGND VGND VPWR VPWR _01765_ sky130_fd_sc_hd__clkbuf_1
X_25758_ _13823_ _13876_ VGND VGND VPWR VPWR _11160_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15511_ _13297_ _13546_ _13294_ _13292_ VGND VGND VPWR VPWR _14038_ sky130_fd_sc_hd__a211o_1
XFILLER_0_35_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24709_ _10562_ VGND VGND VPWR VPWR _02436_ sky130_fd_sc_hd__clkbuf_1
X_16491_ net2697 _14451_ _04478_ VGND VGND VPWR VPWR _04483_ sky130_fd_sc_hd__mux2_1
X_28477_ _12462_ net3493 _12713_ VGND VGND VPWR VPWR _12721_ sky130_fd_sc_hd__mux2_1
X_25689_ _11105_ net1768 _11111_ _11116_ VGND VGND VPWR VPWR _02862_ sky130_fd_sc_hd__a31o_1
XFILLER_0_128_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_216_5672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18230_ _05356_ _05593_ _05594_ VGND VGND VPWR VPWR _05595_ sky130_fd_sc_hd__o21a_1
XFILLER_0_155_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_216_5683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15442_ _13431_ _13628_ _13642_ VGND VGND VPWR VPWR _13973_ sky130_fd_sc_hd__o21a_1
X_27428_ _12137_ VGND VGND VPWR VPWR _03580_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_210_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_182_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18161_ rvcpu.dp.plem.ALUResultM\[25\] _05293_ _05340_ _13200_ VGND VGND VPWR VPWR
+ _05526_ sky130_fd_sc_hd__o22a_1
XFILLER_0_5_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15373_ _13407_ _13448_ _13366_ VGND VGND VPWR VPWR _13907_ sky130_fd_sc_hd__a21o_1
X_27359_ _12080_ net3561 _12097_ VGND VGND VPWR VPWR _12098_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17112_ _04812_ VGND VGND VPWR VPWR _01482_ sky130_fd_sc_hd__clkbuf_1
X_18092_ _05458_ _05459_ VGND VGND VPWR VPWR _05460_ sky130_fd_sc_hd__and2_1
XFILLER_0_145_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30370_ net716 _02105_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[3\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap107 net108 VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_2
X_17043_ net2043 _14457_ _04768_ VGND VGND VPWR VPWR _04776_ sky130_fd_sc_hd__mux2_1
X_29029_ _13026_ VGND VGND VPWR VPWR _04292_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32040_ clknet_leaf_132_clk _03462_ VGND VGND VPWR VPWR datamem.data_ram\[50\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_146_4008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18994_ _06271_ _06328_ _05707_ VGND VGND VPWR VPWR _06329_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23467__115 clknet_1_0__leaf__10158_ VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__inv_2
X_17945_ _05315_ _05316_ VGND VGND VPWR VPWR _05317_ sky130_fd_sc_hd__and2_1
XFILLER_0_209_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_225_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_4399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_218_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32942_ clknet_leaf_134_clk _04364_ VGND VGND VPWR VPWR datamem.data_ram\[6\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_105_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17876_ rvcpu.dp.plde.Rs1E\[1\] rvcpu.dp.plem.RdM\[1\] VGND VGND VPWR VPWR _05249_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_105_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23547__172 clknet_1_0__leaf__10173_ VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__inv_2
XFILLER_0_75_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_105_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19615_ _06591_ _05386_ VGND VGND VPWR VPWR _06911_ sky130_fd_sc_hd__nor2_2
XFILLER_0_221_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16827_ _04661_ VGND VGND VPWR VPWR _01624_ sky130_fd_sc_hd__clkbuf_1
X_32873_ clknet_leaf_56_clk _04295_ VGND VGND VPWR VPWR datamem.data_ram\[10\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_176_4716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_176_4727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31824_ clknet_leaf_105_clk _03278_ VGND VGND VPWR VPWR datamem.data_ram\[16\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_19546_ datamem.data_ram\[26\]\[24\] _06612_ _06838_ _06841_ VGND VGND VPWR VPWR
+ _06842_ sky130_fd_sc_hd__o211a_1
X_16758_ net2824 _14445_ _04623_ VGND VGND VPWR VPWR _04625_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_220_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_66_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15709_ _13250_ VGND VGND VPWR VPWR _14177_ sky130_fd_sc_hd__buf_4
X_31755_ clknet_leaf_58_clk _03209_ VGND VGND VPWR VPWR datamem.data_ram\[45\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_19477_ _06753_ _06759_ _06772_ VGND VGND VPWR VPWR _06773_ sky130_fd_sc_hd__or3_2
XFILLER_0_220_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16689_ _04588_ VGND VGND VPWR VPWR _01697_ sky130_fd_sc_hd__clkbuf_1
X_18428_ _05394_ _05719_ _05790_ _05732_ _05791_ VGND VGND VPWR VPWR _05792_ sky130_fd_sc_hd__o32a_1
XFILLER_0_57_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30706_ clknet_leaf_216_clk _02441_ VGND VGND VPWR VPWR datamem.data_ram\[49\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31686_ clknet_leaf_37_clk _03144_ VGND VGND VPWR VPWR rvcpu.dp.pcreg.q\[4\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_158_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18359_ _05659_ _05722_ _05723_ VGND VGND VPWR VPWR _05724_ sky130_fd_sc_hd__o21ai_2
X_30637_ clknet_leaf_143_clk _02372_ VGND VGND VPWR VPWR datamem.data_ram\[51\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_135_3734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_3745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23816__399 clknet_1_0__leaf__10207_ VGND VGND VPWR VPWR net525 sky130_fd_sc_hd__inv_2
XFILLER_0_16_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21370_ _08535_ VGND VGND VPWR VPWR _08631_ sky130_fd_sc_hd__buf_4
X_30568_ clknet_leaf_142_clk _02303_ VGND VGND VPWR VPWR datamem.data_ram\[54\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_831 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20321_ datamem.data_ram\[27\]\[4\] _06943_ _06926_ datamem.data_ram\[31\]\[4\] _06776_
+ VGND VGND VPWR VPWR _07613_ sky130_fd_sc_hd__a221o_1
XFILLER_0_25_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32307_ clknet_leaf_241_clk _03729_ VGND VGND VPWR VPWR datamem.data_ram\[32\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_23376__1011 clknet_1_1__leaf__10139_ VGND VGND VPWR VPWR net1137 sky130_fd_sc_hd__inv_2
XFILLER_0_141_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold900 rvcpu.dp.rf.reg_file_arr\[6\]\[6\] VGND VGND VPWR VPWR net2050 sky130_fd_sc_hd__dlygate4sd3_1
X_30499_ clknet_leaf_140_clk _02234_ VGND VGND VPWR VPWR datamem.data_ram\[57\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold911 rvcpu.dp.rf.reg_file_arr\[2\]\[16\] VGND VGND VPWR VPWR net2061 sky130_fd_sc_hd__dlygate4sd3_1
Xhold922 datamem.data_ram\[35\]\[3\] VGND VGND VPWR VPWR net2072 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_222_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20252_ datamem.data_ram\[46\]\[3\] _06951_ _06954_ datamem.data_ram\[44\]\[3\] VGND
+ VGND VPWR VPWR _07545_ sky130_fd_sc_hd__a22o_1
Xhold933 datamem.data_ram\[4\]\[23\] VGND VGND VPWR VPWR net2083 sky130_fd_sc_hd__dlygate4sd3_1
X_32238_ clknet_leaf_272_clk _03660_ VGND VGND VPWR VPWR datamem.data_ram\[35\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold944 rvcpu.dp.rf.reg_file_arr\[11\]\[25\] VGND VGND VPWR VPWR net2094 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold955 rvcpu.dp.rf.reg_file_arr\[7\]\[13\] VGND VGND VPWR VPWR net2105 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold966 rvcpu.dp.rf.reg_file_arr\[3\]\[19\] VGND VGND VPWR VPWR net2116 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3002 datamem.data_ram\[16\]\[23\] VGND VGND VPWR VPWR net4152 sky130_fd_sc_hd__dlygate4sd3_1
Xhold977 rvcpu.dp.rf.reg_file_arr\[8\]\[19\] VGND VGND VPWR VPWR net2127 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3013 rvcpu.dp.rf.reg_file_arr\[31\]\[31\] VGND VGND VPWR VPWR net4163 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3024 datamem.data_ram\[21\]\[17\] VGND VGND VPWR VPWR net4174 sky130_fd_sc_hd__dlygate4sd3_1
X_32169_ clknet_leaf_226_clk _03591_ VGND VGND VPWR VPWR datamem.data_ram\[37\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_34_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20183_ datamem.data_ram\[9\]\[11\] _06701_ _07472_ _07475_ VGND VGND VPWR VPWR _07476_
+ sky130_fd_sc_hd__o211a_1
Xhold988 rvcpu.dp.rf.reg_file_arr\[1\]\[1\] VGND VGND VPWR VPWR net2138 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold999 rvcpu.dp.rf.reg_file_arr\[8\]\[18\] VGND VGND VPWR VPWR net2149 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3035 rvcpu.dp.rf.reg_file_arr\[29\]\[8\] VGND VGND VPWR VPWR net4185 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3046 datamem.data_ram\[12\]\[29\] VGND VGND VPWR VPWR net4196 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2301 rvcpu.dp.rf.reg_file_arr\[30\]\[0\] VGND VGND VPWR VPWR net3451 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2312 datamem.data_ram\[34\]\[7\] VGND VGND VPWR VPWR net3462 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold3057 datamem.data_ram\[27\]\[16\] VGND VGND VPWR VPWR net4207 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3068 rvcpu.dp.rf.reg_file_arr\[25\]\[17\] VGND VGND VPWR VPWR net4218 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2323 rvcpu.dp.rf.reg_file_arr\[0\]\[6\] VGND VGND VPWR VPWR net3473 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24991_ _10716_ VGND VGND VPWR VPWR _02564_ sky130_fd_sc_hd__clkbuf_1
Xhold3079 rvcpu.dp.rf.reg_file_arr\[16\]\[25\] VGND VGND VPWR VPWR net4229 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2334 rvcpu.dp.rf.reg_file_arr\[0\]\[9\] VGND VGND VPWR VPWR net3484 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1600 rvcpu.dp.rf.reg_file_arr\[17\]\[17\] VGND VGND VPWR VPWR net2750 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2345 datamem.data_ram\[20\]\[17\] VGND VGND VPWR VPWR net3495 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26730_ _10764_ net3684 _11714_ VGND VGND VPWR VPWR _11721_ sky130_fd_sc_hd__mux2_1
Xhold2356 rvcpu.dp.rf.reg_file_arr\[23\]\[22\] VGND VGND VPWR VPWR net3506 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1611 datamem.data_ram\[34\]\[28\] VGND VGND VPWR VPWR net2761 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2367 datamem.data_ram\[45\]\[16\] VGND VGND VPWR VPWR net3517 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1622 datamem.data_ram\[21\]\[11\] VGND VGND VPWR VPWR net2772 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1633 rvcpu.dp.rf.reg_file_arr\[24\]\[30\] VGND VGND VPWR VPWR net2783 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2378 datamem.data_ram\[54\]\[24\] VGND VGND VPWR VPWR net3528 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1644 datamem.data_ram\[13\]\[26\] VGND VGND VPWR VPWR net2794 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2389 datamem.data_ram\[14\]\[30\] VGND VGND VPWR VPWR net3539 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1655 rvcpu.dp.rf.reg_file_arr\[29\]\[6\] VGND VGND VPWR VPWR net2805 sky130_fd_sc_hd__dlygate4sd3_1
X_26661_ _11665_ net1688 _11675_ _11680_ VGND VGND VPWR VPWR _03270_ sky130_fd_sc_hd__a31o_1
XFILLER_0_212_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1666 rvcpu.dp.rf.reg_file_arr\[10\]\[25\] VGND VGND VPWR VPWR net2816 sky130_fd_sc_hd__dlygate4sd3_1
X_23873_ clknet_1_1__leaf__10203_ VGND VGND VPWR VPWR _10221_ sky130_fd_sc_hd__buf_1
Xhold1677 rvcpu.dp.rf.reg_file_arr\[20\]\[13\] VGND VGND VPWR VPWR net2827 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1688 rvcpu.dp.rf.reg_file_arr\[16\]\[18\] VGND VGND VPWR VPWR net2838 sky130_fd_sc_hd__dlygate4sd3_1
X_28400_ _12676_ VGND VGND VPWR VPWR _04013_ sky130_fd_sc_hd__clkbuf_1
Xhold1699 datamem.data_ram\[48\]\[8\] VGND VGND VPWR VPWR net2849 sky130_fd_sc_hd__dlygate4sd3_1
X_25612_ _11070_ VGND VGND VPWR VPWR _02831_ sky130_fd_sc_hd__clkbuf_1
X_22824_ _09433_ _09962_ _09789_ VGND VGND VPWR VPWR _09963_ sky130_fd_sc_hd__a21o_1
Xclkbuf_0__10261_ _10261_ VGND VGND VPWR VPWR clknet_0__10261_ sky130_fd_sc_hd__clkbuf_16
X_29380_ clknet_leaf_145_clk _01115_ VGND VGND VPWR VPWR datamem.data_ram\[60\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__10161_ clknet_0__10161_ VGND VGND VPWR VPWR clknet_1_1__leaf__10161_
+ sky130_fd_sc_hd__clkbuf_16
X_26592_ _11083_ _11640_ VGND VGND VPWR VPWR _11643_ sky130_fd_sc_hd__and2_1
XFILLER_0_168_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_184_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28331_ _12639_ VGND VGND VPWR VPWR _03981_ sky130_fd_sc_hd__clkbuf_1
X_25543_ _11029_ VGND VGND VPWR VPWR _02803_ sky130_fd_sc_hd__clkbuf_1
X_22755_ rvcpu.dp.rf.reg_file_arr\[12\]\[23\] rvcpu.dp.rf.reg_file_arr\[13\]\[23\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[23\] rvcpu.dp.rf.reg_file_arr\[15\]\[23\] _09462_
+ _09721_ VGND VGND VPWR VPWR _09898_ sky130_fd_sc_hd__mux4_1
Xclkbuf_0__10192_ _10192_ VGND VGND VPWR VPWR clknet_0__10192_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_56_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21706_ _08943_ _08947_ _08951_ _08625_ VGND VGND VPWR VPWR _01044_ sky130_fd_sc_hd__o31a_1
X_25474_ _10991_ net1449 _10984_ _10993_ VGND VGND VPWR VPWR _02770_ sky130_fd_sc_hd__a31o_1
XFILLER_0_164_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28262_ _07125_ VGND VGND VPWR VPWR _12601_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_82_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22686_ rvcpu.dp.rf.reg_file_arr\[16\]\[20\] rvcpu.dp.rf.reg_file_arr\[17\]\[20\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[20\] rvcpu.dp.rf.reg_file_arr\[19\]\[20\] _09512_
+ _09513_ VGND VGND VPWR VPWR _09832_ sky130_fd_sc_hd__mux4_1
XFILLER_0_66_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27213_ _12005_ net1639 _12007_ _12016_ VGND VGND VPWR VPWR _03486_ sky130_fd_sc_hd__a31o_1
X_24425_ _10394_ datamem.data_ram\[53\]\[12\] _10386_ VGND VGND VPWR VPWR _10395_
+ sky130_fd_sc_hd__mux2_1
X_21637_ rvcpu.dp.rf.reg_file_arr\[28\]\[13\] rvcpu.dp.rf.reg_file_arr\[30\]\[13\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[13\] rvcpu.dp.rf.reg_file_arr\[31\]\[13\] _08559_
+ _08636_ VGND VGND VPWR VPWR _08886_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_229_6008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28193_ _12279_ _12345_ _12482_ VGND VGND VPWR VPWR _12564_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_229_6019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27144_ _11946_ _11966_ VGND VGND VPWR VPWR _11975_ sky130_fd_sc_hd__and2_1
X_24356_ _10355_ VGND VGND VPWR VPWR _02290_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21568_ _08695_ _08820_ VGND VGND VPWR VPWR _08821_ sky130_fd_sc_hd__and2_1
XFILLER_0_90_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_185_Right_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_5_16__f_clk clknet_2_2_0_clk VGND VGND VPWR VPWR clknet_5_16__leaf_clk sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_73_Left_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27075_ _11919_ net1733 _11923_ _11930_ VGND VGND VPWR VPWR _03434_ sky130_fd_sc_hd__a31o_1
X_20519_ datamem.data_ram\[29\]\[21\] _06865_ _06672_ datamem.data_ram\[31\]\[21\]
+ VGND VGND VPWR VPWR _07810_ sky130_fd_sc_hd__o22a_1
XFILLER_0_16_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24287_ _09267_ net2858 _10316_ VGND VGND VPWR VPWR _10317_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21499_ _08663_ _08752_ _08754_ _08652_ VGND VGND VPWR VPWR _08755_ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26026_ _11338_ VGND VGND VPWR VPWR _11339_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_127_1074 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_207_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27977_ _09259_ VGND VGND VPWR VPWR _12445_ sky130_fd_sc_hd__clkbuf_2
X_15991_ _14310_ VGND VGND VPWR VPWR _14333_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_206_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29716_ net1062 _01451_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[22\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_17730_ _05117_ VGND VGND VPWR VPWR _05140_ sky130_fd_sc_hd__buf_4
XFILLER_0_206_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14942_ _13449_ _13490_ _13429_ VGND VGND VPWR VPWR _13491_ sky130_fd_sc_hd__o21ai_1
X_26928_ _11825_ _11842_ VGND VGND VPWR VPWR _11844_ sky130_fd_sc_hd__and2_1
XFILLER_0_175_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_82_Left_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29647_ net993 _01382_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[24\]\[10\] sky130_fd_sc_hd__dfxtp_1
Xhold2890 rvcpu.dp.rf.reg_file_arr\[21\]\[10\] VGND VGND VPWR VPWR net4040 sky130_fd_sc_hd__dlygate4sd3_1
X_17661_ _05103_ VGND VGND VPWR VPWR _01208_ sky130_fd_sc_hd__clkbuf_1
X_14873_ _13380_ VGND VGND VPWR VPWR _13425_ sky130_fd_sc_hd__buf_4
XFILLER_0_215_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26859_ _11795_ net1490 _11797_ _11799_ VGND VGND VPWR VPWR _03349_ sky130_fd_sc_hd__a31o_1
XFILLER_0_203_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19400_ _06695_ VGND VGND VPWR VPWR _06696_ sky130_fd_sc_hd__clkbuf_8
X_16612_ _04547_ VGND VGND VPWR VPWR _01733_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_218_5723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_218_5734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29578_ net932 _01313_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[26\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_17592_ _13241_ net3035 _05057_ VGND VGND VPWR VPWR _05067_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19331_ _06626_ VGND VGND VPWR VPWR _06627_ sky130_fd_sc_hd__clkbuf_8
X_28529_ _12754_ net3955 _12752_ VGND VGND VPWR VPWR _12755_ sky130_fd_sc_hd__mux2_1
X_16543_ _04510_ VGND VGND VPWR VPWR _01773_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_171_4602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19262_ _06563_ VGND VGND VPWR VPWR rvcpu.dp.lAuiPCE\[31\] sky130_fd_sc_hd__clkbuf_1
X_31540_ clknet_leaf_75_clk net1261 VGND VGND VPWR VPWR rvcpu.dp.plem.funct3M\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16474_ net2618 _14434_ _04467_ VGND VGND VPWR VPWR _04474_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18213_ _05384_ _05385_ VGND VGND VPWR VPWR _05578_ sky130_fd_sc_hd__and2_1
X_15425_ _13572_ _13939_ _13944_ _13956_ VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__o31a_1
XFILLER_0_155_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19193_ _06487_ _06491_ _06496_ _06495_ VGND VGND VPWR VPWR _06504_ sky130_fd_sc_hd__a31o_1
X_31471_ clknet_leaf_5_clk rvcpu.dp.SrcBFW_Mux.y\[29\] VGND VGND VPWR VPWR rvcpu.dp.plem.WriteDataM\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18144_ rvcpu.dp.plde.ImmExtE\[16\] rvcpu.dp.SrcBFW_Mux.y\[16\] _05278_ VGND VGND
+ VPWR VPWR _05509_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_91_Left_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30422_ net760 _02157_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[29\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_15356_ _13533_ _13890_ _13478_ VGND VGND VPWR VPWR _13891_ sky130_fd_sc_hd__o21a_1
XFILLER_0_124_831 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_152_Right_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18075_ _05425_ VGND VGND VPWR VPWR _05443_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_130_3620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30353_ net699 _02088_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[3\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_15287_ _13823_ _13350_ _13824_ VGND VGND VPWR VPWR _13825_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_169_4542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold207 datamem.data_ram\[43\]\[6\] VGND VGND VPWR VPWR net1357 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_169_4553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__10181_ clknet_0__10181_ VGND VGND VPWR VPWR clknet_1_0__leaf__10181_
+ sky130_fd_sc_hd__clkbuf_16
Xhold218 datamem.data_ram\[7\]\[6\] VGND VGND VPWR VPWR net1368 sky130_fd_sc_hd__dlygate4sd3_1
Xhold229 datamem.data_ram\[16\]\[7\] VGND VGND VPWR VPWR net1379 sky130_fd_sc_hd__dlygate4sd3_1
X_17026_ net2451 _14440_ _04757_ VGND VGND VPWR VPWR _04767_ sky130_fd_sc_hd__mux2_1
XFILLER_0_229_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30284_ clknet_leaf_196_clk _02019_ VGND VGND VPWR VPWR datamem.data_ram\[58\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32023_ clknet_leaf_129_clk _03445_ VGND VGND VPWR VPWR datamem.data_ram\[51\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_91_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18977_ _05866_ _06004_ VGND VGND VPWR VPWR _06313_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_128_3560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17928_ rvcpu.dp.plde.ImmExtE\[28\] rvcpu.dp.SrcBFW_Mux.y\[28\] _05279_ VGND VGND
+ VPWR VPWR _05301_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_3571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22991__697 clknet_1_0__leaf__10084_ VGND VGND VPWR VPWR net823 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_68_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32925_ clknet_leaf_255_clk _04347_ VGND VGND VPWR VPWR datamem.data_ram\[0\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_68_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17859_ _05179_ _05180_ rvcpu.dp.plde.RD2E\[5\] VGND VGND VPWR VPWR _05234_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_124_3468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_3479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20870_ datamem.data_ram\[53\]\[14\] _07037_ _06806_ datamem.data_ram\[52\]\[14\]
+ VGND VGND VPWR VPWR _08160_ sky130_fd_sc_hd__o22a_1
X_32856_ clknet_leaf_185_clk _04278_ VGND VGND VPWR VPWR datamem.data_ram\[11\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_221_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31807_ clknet_leaf_108_clk _03261_ VGND VGND VPWR VPWR datamem.data_ram\[17\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19529_ datamem.data_ram\[46\]\[24\] _06626_ _06812_ datamem.data_ram\[43\]\[24\]
+ _06599_ VGND VGND VPWR VPWR _06825_ sky130_fd_sc_hd__o221a_1
X_32787_ clknet_leaf_250_clk _04209_ VGND VGND VPWR VPWR datamem.data_ram\[14\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22540_ _09399_ _09693_ _09472_ VGND VGND VPWR VPWR _09694_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_27_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31738_ net187 _03196_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[9\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22471_ rvcpu.dp.rf.reg_file_arr\[12\]\[8\] rvcpu.dp.rf.reg_file_arr\[13\]\[8\] rvcpu.dp.rf.reg_file_arr\[14\]\[8\]
+ rvcpu.dp.rf.reg_file_arr\[15\]\[8\] _09552_ _09382_ VGND VGND VPWR VPWR _09629_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_228_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31669_ clknet_leaf_68_clk net1253 VGND VGND VPWR VPWR rvcpu.dp.plmw.ALUResultW\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24210_ _10275_ VGND VGND VPWR VPWR _02224_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_98_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21422_ _08675_ _08677_ _08680_ _08626_ _08510_ VGND VGND VPWR VPWR _08681_ sky130_fd_sc_hd__a221o_1
X_25190_ _10731_ net3638 net57 VGND VGND VPWR VPWR _10833_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21353_ rvcpu.dp.plde.funct3E\[0\] rvcpu.dp.Cout VGND VGND VPWR VPWR _08615_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20304_ _07574_ _07596_ VGND VGND VPWR VPWR _07597_ sky130_fd_sc_hd__nor2_2
Xhold730 rvcpu.dp.rf.reg_file_arr\[1\]\[28\] VGND VGND VPWR VPWR net1880 sky130_fd_sc_hd__dlygate4sd3_1
X_21284_ _08511_ _08545_ VGND VGND VPWR VPWR _08546_ sky130_fd_sc_hd__nor2_1
XFILLER_0_163_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold741 rvcpu.dp.rf.reg_file_arr\[1\]\[29\] VGND VGND VPWR VPWR net1891 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27900_ _11978_ _12394_ VGND VGND VPWR VPWR _12401_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23864__426 clknet_1_1__leaf__10220_ VGND VGND VPWR VPWR net552 sky130_fd_sc_hd__inv_2
Xhold752 rvcpu.dp.rf.reg_file_arr\[4\]\[6\] VGND VGND VPWR VPWR net1902 sky130_fd_sc_hd__dlygate4sd3_1
X_20235_ _06753_ _07522_ _07527_ _06713_ VGND VGND VPWR VPWR _07528_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_57_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold763 rvcpu.dp.rf.reg_file_arr\[6\]\[23\] VGND VGND VPWR VPWR net1913 sky130_fd_sc_hd__dlygate4sd3_1
X_28880_ _12944_ VGND VGND VPWR VPWR _04225_ sky130_fd_sc_hd__clkbuf_1
Xhold774 rvcpu.dp.rf.reg_file_arr\[17\]\[18\] VGND VGND VPWR VPWR net1924 sky130_fd_sc_hd__dlygate4sd3_1
Xhold785 datamem.data_ram\[62\]\[31\] VGND VGND VPWR VPWR net1935 sky130_fd_sc_hd__dlygate4sd3_1
Xhold796 rvcpu.dp.rf.reg_file_arr\[30\]\[14\] VGND VGND VPWR VPWR net1946 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_228_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27831_ _12360_ VGND VGND VPWR VPWR _03760_ sky130_fd_sc_hd__clkbuf_1
X_20166_ _07449_ _07450_ _07453_ _07458_ VGND VGND VPWR VPWR _07459_ sky130_fd_sc_hd__a31o_1
Xhold2120 rvcpu.dp.rf.reg_file_arr\[21\]\[31\] VGND VGND VPWR VPWR net3270 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2131 datamem.data_ram\[45\]\[25\] VGND VGND VPWR VPWR net3281 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2142 datamem.data_ram\[5\]\[29\] VGND VGND VPWR VPWR net3292 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2153 rvcpu.dp.rf.reg_file_arr\[14\]\[27\] VGND VGND VPWR VPWR net3303 sky130_fd_sc_hd__dlygate4sd3_1
X_27762_ _12151_ net2506 net48 VGND VGND VPWR VPWR _12321_ sky130_fd_sc_hd__mux2_1
X_24974_ _10707_ VGND VGND VPWR VPWR _02556_ sky130_fd_sc_hd__clkbuf_1
X_20097_ datamem.data_ram\[2\]\[10\] _06804_ _06687_ datamem.data_ram\[4\]\[10\] VGND
+ VGND VPWR VPWR _07391_ sky130_fd_sc_hd__o22a_1
Xhold2164 rvcpu.dp.rf.reg_file_arr\[31\]\[1\] VGND VGND VPWR VPWR net3314 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2175 rvcpu.dp.rf.reg_file_arr\[27\]\[25\] VGND VGND VPWR VPWR net3325 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1430 rvcpu.dp.rf.reg_file_arr\[31\]\[12\] VGND VGND VPWR VPWR net2580 sky130_fd_sc_hd__dlygate4sd3_1
X_29501_ net863 _01236_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[28\]\[8\] sky130_fd_sc_hd__dfxtp_1
Xhold1441 datamem.data_ram\[39\]\[28\] VGND VGND VPWR VPWR net2591 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2186 datamem.data_ram\[42\]\[25\] VGND VGND VPWR VPWR net3336 sky130_fd_sc_hd__dlygate4sd3_1
X_26713_ _11711_ VGND VGND VPWR VPWR _03291_ sky130_fd_sc_hd__clkbuf_1
Xhold2197 datamem.data_ram\[37\]\[24\] VGND VGND VPWR VPWR net3347 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1452 rvcpu.dp.rf.reg_file_arr\[29\]\[20\] VGND VGND VPWR VPWR net2602 sky130_fd_sc_hd__dlygate4sd3_1
X_27693_ _12284_ VGND VGND VPWR VPWR _03698_ sky130_fd_sc_hd__clkbuf_1
Xhold1463 datamem.data_ram\[61\]\[31\] VGND VGND VPWR VPWR net2613 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1474 rvcpu.dp.rf.reg_file_arr\[16\]\[23\] VGND VGND VPWR VPWR net2624 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1485 datamem.data_ram\[35\]\[31\] VGND VGND VPWR VPWR net2635 sky130_fd_sc_hd__dlygate4sd3_1
X_29432_ net794 _01167_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[30\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_26644_ _11645_ _11663_ VGND VGND VPWR VPWR _11669_ sky130_fd_sc_hd__and2_1
XFILLER_0_212_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_200_5292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1496 rvcpu.dp.rf.reg_file_arr\[23\]\[25\] VGND VGND VPWR VPWR net2646 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_211_131 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0__10244_ _10244_ VGND VGND VPWR VPWR clknet_0__10244_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_131_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22807_ _09636_ _09946_ VGND VGND VPWR VPWR _09947_ sky130_fd_sc_hd__or2_1
X_29363_ clknet_leaf_174_clk _01098_ VGND VGND VPWR VPWR datamem.data_ram\[61\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26511__63 clknet_1_0__leaf__11602_ VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__inv_2
X_26575_ _10731_ net2736 _11629_ VGND VGND VPWR VPWR _11633_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20999_ datamem.data_ram\[26\]\[15\] _06608_ _06631_ datamem.data_ram\[27\]\[15\]
+ VGND VGND VPWR VPWR _08288_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_0_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_192_5093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28314_ _12630_ VGND VGND VPWR VPWR _03973_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_196_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0__10175_ _10175_ VGND VGND VPWR VPWR clknet_0__10175_ sky130_fd_sc_hd__clkbuf_16
X_25526_ _08151_ _09268_ VGND VGND VPWR VPWR _11020_ sky130_fd_sc_hd__nor2_4
XFILLER_0_223_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29294_ clknet_leaf_1_clk _01029_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD1E\[1\] sky130_fd_sc_hd__dfxtp_1
X_22738_ _09469_ _09881_ VGND VGND VPWR VPWR _09882_ sky130_fd_sc_hd__or2_1
XFILLER_0_109_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28245_ _10979_ _12345_ _12573_ VGND VGND VPWR VPWR _12592_ sky130_fd_sc_hd__a21oi_1
X_25457_ _07182_ _10932_ _10044_ VGND VGND VPWR VPWR _10983_ sky130_fd_sc_hd__or3_1
XFILLER_0_165_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22669_ rvcpu.dp.rf.reg_file_arr\[20\]\[19\] rvcpu.dp.rf.reg_file_arr\[21\]\[19\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[19\] rvcpu.dp.rf.reg_file_arr\[23\]\[19\] _09401_
+ _09430_ VGND VGND VPWR VPWR _09816_ sky130_fd_sc_hd__mux4_1
X_15210_ _13750_ _13751_ _13573_ VGND VGND VPWR VPWR _13752_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_129_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24408_ _10383_ VGND VGND VPWR VPWR _02314_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28176_ _12279_ _12335_ _12482_ VGND VGND VPWR VPWR _12555_ sky130_fd_sc_hd__a21oi_4
X_16190_ _13216_ VGND VGND VPWR VPWR _14445_ sky130_fd_sc_hd__buf_4
X_25388_ _08133_ VGND VGND VPWR VPWR _10946_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_11_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15141_ _13328_ _13289_ VGND VGND VPWR VPWR _13685_ sky130_fd_sc_hd__nor2_1
X_27127_ _11956_ net1796 _11952_ _11962_ VGND VGND VPWR VPWR _03454_ sky130_fd_sc_hd__a31o_1
XFILLER_0_106_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24339_ _09260_ net4386 _10338_ VGND VGND VPWR VPWR _10346_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15072_ _13338_ _13617_ _13501_ VGND VGND VPWR VPWR _13618_ sky130_fd_sc_hd__a21oi_1
X_27058_ _11919_ net1870 _11910_ _11920_ VGND VGND VPWR VPWR _03427_ sky130_fd_sc_hd__a31o_1
X_18900_ _05461_ _05627_ _06228_ _05655_ VGND VGND VPWR VPWR _06241_ sky130_fd_sc_hd__a31o_1
XFILLER_0_120_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26009_ net18 _11317_ VGND VGND VPWR VPWR _11330_ sky130_fd_sc_hd__or2_1
X_19880_ datamem.data_ram\[17\]\[1\] _06997_ _07171_ _07174_ VGND VGND VPWR VPWR _07175_
+ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_207_5457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_207_5468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18831_ _05494_ _05732_ VGND VGND VPWR VPWR _06177_ sky130_fd_sc_hd__nor2_1
XFILLER_0_207_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_160_4325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_4336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_4347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18762_ _05307_ _05437_ _05610_ _05408_ _05665_ _05670_ VGND VGND VPWR VPWR _06112_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_199_5269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15974_ _14324_ VGND VGND VPWR VPWR _02040_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_172_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17713_ _05131_ VGND VGND VPWR VPWR _01184_ sky130_fd_sc_hd__clkbuf_1
X_14925_ _13333_ _13364_ VGND VGND VPWR VPWR _13474_ sky130_fd_sc_hd__nand2_2
XFILLER_0_136_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18693_ _06046_ VGND VGND VPWR VPWR _06047_ sky130_fd_sc_hd__inv_2
X_30971_ clknet_leaf_208_clk _02706_ VGND VGND VPWR VPWR datamem.data_ram\[39\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold90 rvcpu.dp.plde.PCPlus4E\[15\] VGND VGND VPWR VPWR net1240 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_136_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32710_ clknet_leaf_83_clk _04132_ VGND VGND VPWR VPWR datamem.data_ram\[17\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_17644_ net2358 _13216_ _05093_ VGND VGND VPWR VPWR _05095_ sky130_fd_sc_hd__mux2_1
X_14856_ _13312_ _13313_ VGND VGND VPWR VPWR _13408_ sky130_fd_sc_hd__and2_1
XFILLER_0_76_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23375__1010 clknet_1_0__leaf__10139_ VGND VGND VPWR VPWR net1136 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_63_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32641_ clknet_leaf_159_clk _04063_ VGND VGND VPWR VPWR datamem.data_ram\[1\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_17575_ _05058_ VGND VGND VPWR VPWR _01249_ sky130_fd_sc_hd__clkbuf_1
X_14787_ _13288_ _13286_ VGND VGND VPWR VPWR _13340_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_221_Right_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_175_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_158_4276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_158_4287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19314_ _06609_ VGND VGND VPWR VPWR _06610_ sky130_fd_sc_hd__buf_8
XFILLER_0_202_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_4298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16526_ net4146 _14486_ _04466_ VGND VGND VPWR VPWR _04501_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32572_ clknet_leaf_253_clk _03994_ VGND VGND VPWR VPWR datamem.data_ram\[22\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_31523_ clknet_leaf_47_clk net1180 VGND VGND VPWR VPWR rvcpu.dp.plem.PCPlus4M\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_19245_ rvcpu.dp.plde.ImmExtE\[29\] rvcpu.dp.plde.PCE\[29\] VGND VGND VPWR VPWR _06549_
+ sky130_fd_sc_hd__nand2_1
X_16457_ _04463_ VGND VGND VPWR VPWR _01812_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15408_ _13649_ VGND VGND VPWR VPWR _13940_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_22_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19176_ _06473_ _06476_ _06481_ _06480_ VGND VGND VPWR VPWR _06489_ sky130_fd_sc_hd__a31o_1
XFILLER_0_143_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31454_ clknet_leaf_7_clk rvcpu.dp.SrcBFW_Mux.y\[12\] VGND VGND VPWR VPWR rvcpu.dp.plem.WriteDataM\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_22_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16388_ net2018 _14486_ _14524_ VGND VGND VPWR VPWR _14559_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18127_ rvcpu.dp.plde.ImmExtE\[18\] rvcpu.dp.SrcBFW_Mux.y\[18\] _05278_ VGND VGND
+ VPWR VPWR _05493_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_3294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30405_ net743 _02140_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[31\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_15339_ _13409_ _13459_ _13488_ _13521_ VGND VGND VPWR VPWR _13875_ sky130_fd_sc_hd__a31o_1
XFILLER_0_14_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31385_ clknet_leaf_32_clk _03088_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCE\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_93_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18058_ _05421_ _05424_ VGND VGND VPWR VPWR _05426_ sky130_fd_sc_hd__nor2_1
X_30336_ net682 _02071_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[4\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17009_ _04758_ VGND VGND VPWR VPWR _01531_ sky130_fd_sc_hd__clkbuf_1
X_30267_ net621 _02002_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[6\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20020_ datamem.data_ram\[38\]\[2\] _06951_ _07310_ _07313_ VGND VGND VPWR VPWR _07314_
+ sky130_fd_sc_hd__a211o_1
X_32006_ clknet_leaf_133_clk _03428_ VGND VGND VPWR VPWR datamem.data_ram\[52\]\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_158_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_226_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_3508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_3519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30198_ net552 _01933_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[8\]\[17\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_52_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21971_ _09196_ _09198_ _09201_ _08557_ VGND VGND VPWR VPWR _09202_ sky130_fd_sc_hd__a22o_1
XFILLER_0_213_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_193_1267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20922_ datamem.data_ram\[40\]\[22\] datamem.data_ram\[41\]\[22\] _07827_ VGND VGND
+ VPWR VPWR _08212_ sky130_fd_sc_hd__mux2_1
X_24690_ _10542_ _10114_ _10501_ VGND VGND VPWR VPWR _10552_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_55_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32908_ clknet_leaf_258_clk _04330_ VGND VGND VPWR VPWR datamem.data_ram\[7\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23641_ _09282_ net3085 _10182_ VGND VGND VPWR VPWR _10187_ sky130_fd_sc_hd__mux2_1
X_20853_ datamem.data_ram\[1\]\[14\] _06658_ _08140_ _08142_ VGND VGND VPWR VPWR _08143_
+ sky130_fd_sc_hd__o211a_1
X_32839_ clknet_leaf_282_clk _04261_ VGND VGND VPWR VPWR datamem.data_ram\[12\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26360_ _11083_ _11511_ VGND VGND VPWR VPWR _11514_ sky130_fd_sc_hd__and2_1
XFILLER_0_194_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23572_ clknet_1_0__leaf__10172_ VGND VGND VPWR VPWR _10176_ sky130_fd_sc_hd__buf_1
XFILLER_0_159_591 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20784_ datamem.data_ram\[2\]\[30\] _07023_ _06739_ datamem.data_ram\[3\]\[30\] _08073_
+ VGND VGND VPWR VPWR _08074_ sky130_fd_sc_hd__o221a_1
XFILLER_0_187_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25311_ _10900_ VGND VGND VPWR VPWR _02700_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_46_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22523_ _09442_ _09673_ _09675_ _09677_ VGND VGND VPWR VPWR _09678_ sky130_fd_sc_hd__o2bb2a_1
X_26291_ _11413_ VGND VGND VPWR VPWR _11478_ sky130_fd_sc_hd__buf_2
XFILLER_0_76_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_228_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28030_ _12477_ VGND VGND VPWR VPWR _03842_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25242_ _10731_ net2668 net55 VGND VGND VPWR VPWR _10861_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22454_ _09389_ _09602_ _09607_ _09612_ VGND VGND VPWR VPWR _09613_ sky130_fd_sc_hd__and4_1
XFILLER_0_134_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_924 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21405_ rvcpu.dp.rf.reg_file_arr\[8\]\[2\] rvcpu.dp.rf.reg_file_arr\[10\]\[2\] rvcpu.dp.rf.reg_file_arr\[9\]\[2\]
+ rvcpu.dp.rf.reg_file_arr\[11\]\[2\] _08560_ _08561_ VGND VGND VPWR VPWR _08665_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_59_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25173_ _09321_ VGND VGND VPWR VPWR _10822_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_59_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22385_ rvcpu.dp.rf.reg_file_arr\[0\]\[4\] rvcpu.dp.rf.reg_file_arr\[1\]\[4\] rvcpu.dp.rf.reg_file_arr\[2\]\[4\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[4\] _09417_ _09419_ VGND VGND VPWR VPWR _09547_ sky130_fd_sc_hd__mux4_1
XFILLER_0_161_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21336_ _08588_ _08597_ rvcpu.dp.hu.ResultSrcE0 VGND VGND VPWR VPWR _08598_ sky130_fd_sc_hd__o21ai_4
X_29981_ net351 _01716_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[14\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28932_ _12758_ net2655 _12968_ VGND VGND VPWR VPWR _12972_ sky130_fd_sc_hd__mux2_1
Xhold560 datamem.data_ram\[14\]\[3\] VGND VGND VPWR VPWR net1710 sky130_fd_sc_hd__dlygate4sd3_1
X_21267_ rvcpu.dp.rf.reg_file_arr\[20\]\[0\] rvcpu.dp.rf.reg_file_arr\[21\]\[0\] rvcpu.dp.rf.reg_file_arr\[22\]\[0\]
+ rvcpu.dp.rf.reg_file_arr\[23\]\[0\] _08525_ _08528_ VGND VGND VPWR VPWR _08529_
+ sky130_fd_sc_hd__mux4_1
Xhold571 datamem.data_ram\[19\]\[4\] VGND VGND VPWR VPWR net1721 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold582 datamem.data_ram\[5\]\[1\] VGND VGND VPWR VPWR net1732 sky130_fd_sc_hd__dlygate4sd3_1
Xhold593 datamem.data_ram\[17\]\[5\] VGND VGND VPWR VPWR net1743 sky130_fd_sc_hd__dlygate4sd3_1
X_20218_ datamem.data_ram\[25\]\[3\] _06949_ _07510_ _06680_ VGND VGND VPWR VPWR _07511_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_229_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28863_ _12935_ VGND VGND VPWR VPWR _04217_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_204_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21198_ _08471_ _08480_ VGND VGND VPWR VPWR _08481_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27814_ _12149_ net2991 net78 VGND VGND VPWR VPWR _12350_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_217_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_202_5332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20149_ datamem.data_ram\[58\]\[27\] _06611_ _07438_ _07441_ VGND VGND VPWR VPWR
+ _07442_ sky130_fd_sc_hd__o211a_1
XFILLER_0_218_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_205_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_202_5343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28794_ _12739_ net4186 net70 VGND VGND VPWR VPWR _12899_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_202_5354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27745_ _12134_ net2578 _12307_ VGND VGND VPWR VPWR _12312_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24957_ _10388_ net2992 _10696_ VGND VGND VPWR VPWR _10698_ sky130_fd_sc_hd__mux2_1
XFILLER_0_188_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1260 datamem.data_ram\[11\]\[29\] VGND VGND VPWR VPWR net2410 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_213_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14710_ _13267_ VGND VGND VPWR VPWR _03176_ sky130_fd_sc_hd__clkbuf_1
Xhold1271 rvcpu.dp.rf.reg_file_arr\[3\]\[24\] VGND VGND VPWR VPWR net2421 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_194_5144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1282 datamem.data_ram\[42\]\[24\] VGND VGND VPWR VPWR net2432 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_194_5155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1293 datamem.data_ram\[15\]\[16\] VGND VGND VPWR VPWR net2443 sky130_fd_sc_hd__dlygate4sd3_1
X_27676_ _12089_ net3141 net51 VGND VGND VPWR VPWR _12275_ sky130_fd_sc_hd__mux2_1
X_15690_ _13231_ VGND VGND VPWR VPWR _14164_ sky130_fd_sc_hd__buf_4
X_24888_ _10442_ net3647 _10659_ VGND VGND VPWR VPWR _10661_ sky130_fd_sc_hd__mux2_1
XANTENNA_400 _06617_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_411 _06647_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29415_ clknet_leaf_11_clk _01150_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD2E\[26\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_422 _06776_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_200_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26627_ _10064_ _11659_ _11660_ net1348 VGND VGND VPWR VPWR _03256_ sky130_fd_sc_hd__a22o_1
XANTENNA_433 _06821_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14641_ _13215_ VGND VGND VPWR VPWR _03193_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_213_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_444 _07070_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23839_ _09322_ net2687 _10210_ VGND VGND VPWR VPWR _10216_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_455 _08144_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_0__10227_ _10227_ VGND VGND VPWR VPWR clknet_0__10227_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_71_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_466 _08744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_1_1__f__10127_ clknet_0__10127_ VGND VGND VPWR VPWR clknet_1_1__leaf__10127_
+ sky130_fd_sc_hd__clkbuf_16
X_29346_ clknet_leaf_205_clk _01081_ VGND VGND VPWR VPWR datamem.data_ram\[61\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_477 _09317_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17360_ _04944_ VGND VGND VPWR VPWR _01358_ sky130_fd_sc_hd__clkbuf_1
X_26558_ _10818_ net2966 _11620_ VGND VGND VPWR VPWR _11624_ sky130_fd_sc_hd__mux2_1
XANTENNA_488 _09490_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_499 _11089_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_1194 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16311_ _14518_ VGND VGND VPWR VPWR _01881_ sky130_fd_sc_hd__clkbuf_1
X_25509_ _10405_ _11010_ VGND VGND VPWR VPWR _11011_ sky130_fd_sc_hd__and2_1
Xclkbuf_0__10158_ _10158_ VGND VGND VPWR VPWR clknet_0__10158_ sky130_fd_sc_hd__clkbuf_16
X_17291_ net4439 _13197_ _04902_ VGND VGND VPWR VPWR _04908_ sky130_fd_sc_hd__mux2_1
X_29277_ _09297_ net2342 _13159_ VGND VGND VPWR VPWR _13160_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_153_4162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19030_ rvcpu.dp.plde.ImmExtE\[2\] rvcpu.dp.plde.PCE\[2\] VGND VGND VPWR VPWR _06361_
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_153_4173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28228_ _10979_ _12335_ _12573_ VGND VGND VPWR VPWR _12583_ sky130_fd_sc_hd__a21oi_4
X_16242_ _13268_ VGND VGND VPWR VPWR _14480_ sky130_fd_sc_hd__buf_4
XFILLER_0_153_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__10089_ _10089_ VGND VGND VPWR VPWR clknet_0__10089_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_36_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16173_ _14433_ VGND VGND VPWR VPWR _01942_ sky130_fd_sc_hd__clkbuf_1
X_28159_ _12279_ _12325_ _12482_ VGND VGND VPWR VPWR _12546_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_209_5508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_209_5519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_328 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15124_ _13668_ _13451_ _13423_ _13324_ VGND VGND VPWR VPWR _13669_ sky130_fd_sc_hd__a211o_1
XFILLER_0_140_439 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31170_ clknet_leaf_13_clk rvcpu.ALUResultE\[29\] VGND VGND VPWR VPWR rvcpu.dp.plem.ALUResultM\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_3180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30121_ net483 _01856_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[10\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15055_ _13449_ _13490_ _13597_ _13601_ _13327_ VGND VGND VPWR VPWR _13602_ sky130_fd_sc_hd__o311a_1
X_19932_ rvcpu.dp.plem.ALUResultM\[0\] _06586_ _06987_ _06915_ VGND VGND VPWR VPWR
+ _07227_ sky130_fd_sc_hd__o31a_1
XFILLER_0_120_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_3191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19863_ datamem.data_ram\[2\]\[1\] _07136_ _07133_ datamem.data_ram\[1\]\[1\] _07157_
+ VGND VGND VPWR VPWR _07158_ sky130_fd_sc_hd__a221o_1
X_30052_ net414 _01787_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[12\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_183_4881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_4892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24187__27 clknet_1_1__leaf__10266_ VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__inv_2
XFILLER_0_208_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18814_ _05503_ _05785_ _05974_ _05502_ VGND VGND VPWR VPWR _06161_ sky130_fd_sc_hd__a2bb2o_1
X_19794_ datamem.data_ram\[50\]\[9\] _07023_ _07084_ _07088_ VGND VGND VPWR VPWR _07089_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_223_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18745_ _05941_ _06095_ _05697_ VGND VGND VPWR VPWR _06096_ sky130_fd_sc_hd__mux2_1
X_15957_ _14315_ VGND VGND VPWR VPWR _02048_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_121_3405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14908_ rvcpu.dp.pcreg.q\[8\] _13313_ VGND VGND VPWR VPWR _13458_ sky130_fd_sc_hd__nand2_4
XFILLER_0_163_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18676_ _06029_ _06030_ VGND VGND VPWR VPWR _06031_ sky130_fd_sc_hd__nand2_1
X_30954_ clknet_leaf_279_clk _02689_ VGND VGND VPWR VPWR datamem.data_ram\[3\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_86_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15888_ net3310 _13190_ _14275_ VGND VGND VPWR VPWR _14279_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17627_ net4360 _13189_ _05082_ VGND VGND VPWR VPWR _05086_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14839_ _13387_ _13391_ VGND VGND VPWR VPWR _13392_ sky130_fd_sc_hd__nand2_2
X_30885_ clknet_leaf_224_clk _02620_ VGND VGND VPWR VPWR datamem.data_ram\[42\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_82_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_82_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32624_ clknet_leaf_274_clk _04046_ VGND VGND VPWR VPWR datamem.data_ram\[20\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_17558_ _05049_ VGND VGND VPWR VPWR _01257_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16509_ _04492_ VGND VGND VPWR VPWR _01789_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_119_3345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23592__213 clknet_1_1__leaf__10177_ VGND VGND VPWR VPWR net339 sky130_fd_sc_hd__inv_2
X_32555_ clknet_leaf_240_clk _03977_ VGND VGND VPWR VPWR datamem.data_ram\[22\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_3356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17489_ _13187_ net4005 _05010_ VGND VGND VPWR VPWR _05013_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31506_ clknet_leaf_67_clk net1277 VGND VGND VPWR VPWR rvcpu.dp.plem.PCPlus4M\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_19228_ _06533_ _06530_ _06527_ VGND VGND VPWR VPWR _06534_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_160_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32486_ clknet_leaf_246_clk _03908_ VGND VGND VPWR VPWR datamem.data_ram\[25\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31437_ clknet_leaf_103_clk _03140_ VGND VGND VPWR VPWR datamem.data_ram\[14\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_19159_ rvcpu.dp.plde.ImmExtE\[18\] rvcpu.dp.plde.PCE\[18\] VGND VGND VPWR VPWR _06474_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_147_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_586 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24069__595 clknet_1_1__leaf__10248_ VGND VGND VPWR VPWR net721 sky130_fd_sc_hd__inv_2
XFILLER_0_169_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22170_ _09356_ VGND VGND VPWR VPWR _01103_ sky130_fd_sc_hd__clkbuf_1
X_31368_ clknet_leaf_17_clk _03071_ VGND VGND VPWR VPWR rvcpu.dp.plde.ImmExtE\[17\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_83_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21121_ _06666_ datamem.data_ram\[47\]\[23\] VGND VGND VPWR VPWR _08410_ sky130_fd_sc_hd__and2_1
X_30319_ net665 _02054_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[4\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_54_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31299_ clknet_leaf_40_clk _03002_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCPlus4E\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23709__303 clknet_1_1__leaf__10196_ VGND VGND VPWR VPWR net429 sky130_fd_sc_hd__inv_2
X_21052_ datamem.data_ram\[34\]\[31\] datamem.data_ram\[35\]\[31\] _07911_ VGND VGND
+ VPWR VPWR _08341_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__10078_ clknet_0__10078_ VGND VGND VPWR VPWR clknet_1_0__leaf__10078_
+ sky130_fd_sc_hd__clkbuf_16
X_20003_ datamem.data_ram\[27\]\[2\] _06942_ _07293_ _07296_ VGND VGND VPWR VPWR _07297_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_201_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25860_ rvcpu.dp.pcreg.q\[28\] _11234_ VGND VGND VPWR VPWR _11240_ sky130_fd_sc_hd__nor2_1
XFILLER_0_214_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24811_ _10452_ net3628 _10612_ VGND VGND VPWR VPWR _10619_ sky130_fd_sc_hd__mux2_1
XFILLER_0_226_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25791_ rvcpu.dp.pcreg.q\[14\] _11182_ VGND VGND VPWR VPWR _11185_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27530_ _10542_ _10908_ _12168_ VGND VGND VPWR VPWR _12197_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_2_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24742_ _10570_ _10347_ _10501_ VGND VGND VPWR VPWR _10580_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_2_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21954_ rvcpu.dp.rf.reg_file_arr\[0\]\[30\] rvcpu.dp.rf.reg_file_arr\[1\]\[30\] rvcpu.dp.rf.reg_file_arr\[2\]\[30\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[30\] _08566_ _08569_ VGND VGND VPWR VPWR _09186_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_96_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20905_ datamem.data_ram\[9\]\[22\] _06701_ _08194_ _07081_ VGND VGND VPWR VPWR _08195_
+ sky130_fd_sc_hd__o211a_1
X_27461_ _12080_ net3347 net83 VGND VGND VPWR VPWR _12160_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24673_ _10542_ _10092_ _10501_ VGND VGND VPWR VPWR _10543_ sky130_fd_sc_hd__a21oi_4
X_21885_ _08682_ _09118_ _09120_ _08558_ VGND VGND VPWR VPWR _09121_ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29200_ _09321_ net3239 _13112_ VGND VGND VPWR VPWR _13118_ sky130_fd_sc_hd__mux2_1
X_26412_ _06418_ _11522_ VGND VGND VPWR VPWR _11552_ sky130_fd_sc_hd__and2_1
XFILLER_0_193_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20836_ datamem.data_ram\[28\]\[14\] datamem.data_ram\[29\]\[14\] _07828_ VGND VGND
+ VPWR VPWR _08126_ sky130_fd_sc_hd__mux2_1
X_27392_ _12115_ VGND VGND VPWR VPWR _03566_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_13_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29131_ _13081_ VGND VGND VPWR VPWR _04339_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26343_ _11039_ _10600_ VGND VGND VPWR VPWR _11507_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_13_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20767_ datamem.data_ram\[53\]\[6\] _06970_ _07125_ datamem.data_ram\[55\]\[6\] VGND
+ VGND VPWR VPWR _08057_ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_572 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29062_ _09281_ net2778 net65 VGND VGND VPWR VPWR _13045_ sky130_fd_sc_hd__mux2_1
X_22506_ _09441_ _09661_ VGND VGND VPWR VPWR _09662_ sky130_fd_sc_hd__nor2_1
X_26274_ _11469_ VGND VGND VPWR VPWR _03094_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20698_ datamem.data_ram\[5\]\[5\] _06969_ _06955_ datamem.data_ram\[4\]\[5\] VGND
+ VGND VPWR VPWR _07989_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_767 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28013_ _12468_ VGND VGND VPWR VPWR _03834_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25225_ _10758_ net3969 _10848_ VGND VGND VPWR VPWR _10852_ sky130_fd_sc_hd__mux2_1
X_22437_ _09511_ _09595_ VGND VGND VPWR VPWR _09596_ sky130_fd_sc_hd__or2_1
XFILLER_0_162_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25156_ _10810_ VGND VGND VPWR VPWR _02635_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22368_ _09415_ _09527_ _09530_ VGND VGND VPWR VPWR _09531_ sky130_fd_sc_hd__a21o_1
X_21319_ rvcpu.dp.plfd.InstrD\[16\] VGND VGND VPWR VPWR _08581_ sky130_fd_sc_hd__inv_2
X_24107_ clknet_1_0__leaf__10244_ VGND VGND VPWR VPWR _10259_ sky130_fd_sc_hd__buf_1
X_25087_ _10737_ net2117 _10768_ VGND VGND VPWR VPWR _10775_ sky130_fd_sc_hd__mux2_1
X_29964_ net334 _01699_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[15\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22299_ _09463_ VGND VGND VPWR VPWR _09464_ sky130_fd_sc_hd__buf_6
XFILLER_0_130_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28915_ _12694_ net4126 _12959_ VGND VGND VPWR VPWR _12963_ sky130_fd_sc_hd__mux2_1
Xhold390 datamem.data_ram\[60\]\[4\] VGND VGND VPWR VPWR net1540 sky130_fd_sc_hd__dlygate4sd3_1
X_29895_ net273 _01630_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[17\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_16860_ _04678_ VGND VGND VPWR VPWR _01608_ sky130_fd_sc_hd__clkbuf_1
X_28846_ _12926_ VGND VGND VPWR VPWR _04209_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_217_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_196_5206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15811_ net1930 _13173_ _14236_ VGND VGND VPWR VPWR _14237_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_221_5796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28777_ _12756_ net4123 _12887_ VGND VGND VPWR VPWR _12890_ sky130_fd_sc_hd__mux2_1
X_16791_ net2220 _14478_ _04634_ VGND VGND VPWR VPWR _04642_ sky130_fd_sc_hd__mux2_1
X_25989_ net8 _11317_ VGND VGND VPWR VPWR _11319_ sky130_fd_sc_hd__or2_1
X_18530_ _05890_ VGND VGND VPWR VPWR _05891_ sky130_fd_sc_hd__inv_2
XFILLER_0_204_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15742_ _14127_ net4163 _14199_ VGND VGND VPWR VPWR _14200_ sky130_fd_sc_hd__mux2_1
X_27728_ _12089_ net3094 net49 VGND VGND VPWR VPWR _12303_ sky130_fd_sc_hd__mux2_1
XFILLER_0_204_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1090 rvcpu.dp.rf.reg_file_arr\[28\]\[16\] VGND VGND VPWR VPWR net2240 sky130_fd_sc_hd__dlygate4sd3_1
X_18461_ _05822_ _05823_ _05674_ VGND VGND VPWR VPWR _05824_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_217_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27659_ _12151_ net3881 net79 VGND VGND VPWR VPWR _12266_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15673_ _14151_ net3884 _14152_ VGND VGND VPWR VPWR _14153_ sky130_fd_sc_hd__mux2_1
XANTENNA_230 _10072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_193_clk clknet_5_22__leaf_clk VGND VGND VPWR VPWR clknet_leaf_193_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_241 _11083_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_4213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17412_ _04971_ VGND VGND VPWR VPWR _01333_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_252 _13195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_4224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14624_ _13202_ VGND VGND VPWR VPWR _03197_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_263 _13216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_185_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18392_ _05300_ _05663_ _05755_ VGND VGND VPWR VPWR _05756_ sky130_fd_sc_hd__o21ai_1
X_30670_ clknet_leaf_177_clk _02405_ VGND VGND VPWR VPWR datamem.data_ram\[50\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_274 _13235_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23083__764 clknet_1_1__leaf__10091_ VGND VGND VPWR VPWR net890 sky130_fd_sc_hd__inv_2
XANTENNA_285 _13272_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_201_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_296 _13638_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29329_ clknet_leaf_145_clk _01064_ VGND VGND VPWR VPWR datamem.data_ram\[62\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_17343_ rvcpu.dp.rf.reg_file_arr\[24\]\[1\] _13274_ _04901_ VGND VGND VPWR VPWR _04935_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_184_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32340_ clknet_leaf_232_clk _03762_ VGND VGND VPWR VPWR datamem.data_ram\[30\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_17274_ _14193_ net3021 _04864_ VGND VGND VPWR VPWR _04898_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_183_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19013_ _05755_ _06345_ _06346_ _05671_ _05677_ VGND VGND VPWR VPWR _06347_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_114_3220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16225_ net2279 _14468_ _14464_ VGND VGND VPWR VPWR _14469_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_114_3231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload205 clknet_leaf_199_clk VGND VGND VPWR VPWR clkload205/Y sky130_fd_sc_hd__clkinv_1
XFILLER_0_107_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32271_ clknet_leaf_187_clk _03693_ VGND VGND VPWR VPWR datamem.data_ram\[33\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload216 clknet_leaf_167_clk VGND VGND VPWR VPWR clkload216/Y sky130_fd_sc_hd__clkinv_1
XTAP_TAPCELL_ROW_114_3242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload227 clknet_leaf_91_clk VGND VGND VPWR VPWR clkload227/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_141_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload238 clknet_leaf_118_clk VGND VGND VPWR VPWR clkload238/Y sky130_fd_sc_hd__inv_6
XFILLER_0_12_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31222_ clknet_leaf_38_clk _02925_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCD\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload249 clknet_leaf_152_clk VGND VGND VPWR VPWR clkload249/Y sky130_fd_sc_hd__bufinv_16
X_16156_ _14421_ VGND VGND VPWR VPWR _14422_ sky130_fd_sc_hd__buf_4
XFILLER_0_80_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_185_4932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_185_4943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15107_ _13463_ _13641_ _13647_ _13651_ VGND VGND VPWR VPWR _13652_ sky130_fd_sc_hd__a211o_1
XFILLER_0_140_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31153_ clknet_leaf_69_clk rvcpu.ALUResultE\[12\] VGND VGND VPWR VPWR rvcpu.dp.plem.ALUResultM\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16087_ _14384_ VGND VGND VPWR VPWR _14385_ sky130_fd_sc_hd__buf_4
XFILLER_0_224_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_181_4829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30104_ net466 _01839_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[11\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_15038_ _13332_ _13562_ _13427_ VGND VGND VPWR VPWR _13585_ sky130_fd_sc_hd__or3_1
X_19915_ datamem.data_ram\[37\]\[17\] _06664_ _06658_ datamem.data_ram\[33\]\[17\]
+ VGND VGND VPWR VPWR _07210_ sky130_fd_sc_hd__o22a_1
XFILLER_0_227_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31084_ clknet_leaf_114_clk _02819_ VGND VGND VPWR VPWR datamem.data_ram\[20\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2708 datamem.data_ram\[20\]\[13\] VGND VGND VPWR VPWR net3858 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2719 datamem.data_ram\[51\]\[12\] VGND VGND VPWR VPWR net3869 sky130_fd_sc_hd__dlygate4sd3_1
X_30035_ net397 _01770_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[13\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_19846_ _07131_ _07135_ _07140_ VGND VGND VPWR VPWR _07141_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_88_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19777_ datamem.data_ram\[38\]\[9\] _06683_ _06688_ datamem.data_ram\[36\]\[9\] VGND
+ VGND VPWR VPWR _07072_ sky130_fd_sc_hd__o22a_1
X_16989_ net1943 _14472_ _04742_ VGND VGND VPWR VPWR _04747_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_108_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18728_ _05917_ _06079_ _05697_ VGND VGND VPWR VPWR _06080_ sky130_fd_sc_hd__mux2_1
X_31986_ clknet_leaf_116_clk _03408_ VGND VGND VPWR VPWR datamem.data_ram\[37\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_140_3847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_140_3858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18659_ _05998_ _05999_ _06014_ VGND VGND VPWR VPWR rvcpu.ALUResultE\[8\] sky130_fd_sc_hd__a21o_1
X_30937_ clknet_leaf_264_clk _02672_ VGND VGND VPWR VPWR datamem.data_ram\[40\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_204_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_203_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_184_clk clknet_5_22__leaf_clk VGND VGND VPWR VPWR clknet_leaf_184_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_188_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xwire68 _12950_ VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__buf_4
XFILLER_0_203_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_176_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23600__220 clknet_1_1__leaf__10178_ VGND VGND VPWR VPWR net346 sky130_fd_sc_hd__inv_2
XFILLER_0_176_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21670_ rvcpu.dp.rf.reg_file_arr\[16\]\[15\] rvcpu.dp.rf.reg_file_arr\[17\]\[15\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[15\] rvcpu.dp.rf.reg_file_arr\[19\]\[15\] _08799_
+ _08800_ VGND VGND VPWR VPWR _08917_ sky130_fd_sc_hd__mux4_2
XFILLER_0_4_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30868_ clknet_leaf_3_clk _02603_ VGND VGND VPWR VPWR datamem.data_ram\[43\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23207__858 clknet_1_1__leaf__10112_ VGND VGND VPWR VPWR net984 sky130_fd_sc_hd__inv_2
XFILLER_0_8_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_191_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20621_ _07911_ VGND VGND VPWR VPWR _07912_ sky130_fd_sc_hd__buf_6
XFILLER_0_175_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32607_ clknet_leaf_183_clk _04029_ VGND VGND VPWR VPWR datamem.data_ram\[20\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_1106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30799_ clknet_leaf_202_clk _02534_ VGND VGND VPWR VPWR datamem.data_ram\[45\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20552_ datamem.data_ram\[0\]\[21\] datamem.data_ram\[1\]\[21\] datamem.data_ram\[2\]\[21\]
+ datamem.data_ram\[3\]\[21\] _07837_ _07822_ VGND VGND VPWR VPWR _07843_ sky130_fd_sc_hd__mux4_1
X_32538_ clknet_leaf_81_clk _03960_ VGND VGND VPWR VPWR datamem.data_ram\[23\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_138_3798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32469_ clknet_leaf_78_clk _03891_ VGND VGND VPWR VPWR datamem.data_ram\[26\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_20483_ datamem.data_ram\[63\]\[20\] _06668_ _06654_ datamem.data_ram\[57\]\[20\]
+ VGND VGND VPWR VPWR _07775_ sky130_fd_sc_hd__o22a_1
XFILLER_0_162_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25010_ _09272_ VGND VGND VPWR VPWR _10727_ sky130_fd_sc_hd__buf_2
X_22222_ _09380_ _09383_ _09386_ _09387_ _08622_ VGND VGND VPWR VPWR _09388_ sky130_fd_sc_hd__o41a_1
XFILLER_0_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22153_ _09346_ VGND VGND VPWR VPWR _01096_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_203_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21104_ _06615_ _08387_ _08392_ _06677_ VGND VGND VPWR VPWR _08393_ sky130_fd_sc_hd__a211o_1
X_26961_ _11849_ net1421 _11853_ _11862_ VGND VGND VPWR VPWR _03388_ sky130_fd_sc_hd__a31o_1
X_22084_ _09297_ VGND VGND VPWR VPWR _09298_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_160_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28700_ _12848_ VGND VGND VPWR VPWR _04141_ sky130_fd_sc_hd__clkbuf_1
X_25912_ _11153_ VGND VGND VPWR VPWR _11275_ sky130_fd_sc_hd__buf_2
X_21035_ _08321_ _08322_ _08323_ VGND VGND VPWR VPWR _08324_ sky130_fd_sc_hd__and3_1
X_29680_ net1026 _01415_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[23\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_7_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26892_ _11813_ net1575 _11809_ _11818_ VGND VGND VPWR VPWR _03363_ sky130_fd_sc_hd__a31o_1
X_28631_ _12764_ net2035 _12805_ VGND VGND VPWR VPWR _12812_ sky130_fd_sc_hd__mux2_1
X_25843_ rvcpu.dp.pcreg.q\[25\] _11221_ VGND VGND VPWR VPWR _11226_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_198_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28562_ _12700_ net2203 _12768_ VGND VGND VPWR VPWR _12775_ sky130_fd_sc_hd__mux2_1
X_24119__625 clknet_1_1__leaf__10260_ VGND VGND VPWR VPWR net751 sky130_fd_sc_hd__inv_2
X_25774_ rvcpu.dp.pcreg.q\[10\] _11168_ VGND VGND VPWR VPWR _11172_ sky130_fd_sc_hd__nor2_1
XFILLER_0_214_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23599__219 clknet_1_1__leaf__10178_ VGND VGND VPWR VPWR net345 sky130_fd_sc_hd__inv_2
XFILLER_0_97_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27513_ _10542_ _10898_ _12168_ VGND VGND VPWR VPWR _12188_ sky130_fd_sc_hd__a21oi_2
X_24725_ _10570_ _10337_ _10501_ VGND VGND VPWR VPWR _10571_ sky130_fd_sc_hd__a21oi_4
X_28493_ _11976_ _12724_ VGND VGND VPWR VPWR _12731_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_175_clk clknet_5_24__leaf_clk VGND VGND VPWR VPWR clknet_leaf_175_clk
+ sky130_fd_sc_hd__clkbuf_8
X_21937_ rvcpu.dp.rf.reg_file_arr\[4\]\[29\] rvcpu.dp.rf.reg_file_arr\[5\]\[29\] rvcpu.dp.rf.reg_file_arr\[6\]\[29\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[29\] _08578_ _08684_ VGND VGND VPWR VPWR _09170_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_210_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27444_ _12148_ VGND VGND VPWR VPWR _03585_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24656_ _10412_ net1446 _10531_ _10533_ VGND VGND VPWR VPWR _02412_ sky130_fd_sc_hd__a31o_1
XFILLER_0_38_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21868_ rvcpu.dp.rf.reg_file_arr\[4\]\[25\] rvcpu.dp.rf.reg_file_arr\[5\]\[25\] rvcpu.dp.rf.reg_file_arr\[6\]\[25\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[25\] _08839_ _08840_ VGND VGND VPWR VPWR _09105_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_210_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_194_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20819_ datamem.data_ram\[31\]\[30\] _07860_ _06934_ datamem.data_ram\[25\]\[30\]
+ VGND VGND VPWR VPWR _08109_ sky130_fd_sc_hd__o22a_1
X_27375_ net112 _10896_ VGND VGND VPWR VPWR _12106_ sky130_fd_sc_hd__nor2_8
X_21799_ rvcpu.dp.rf.reg_file_arr\[16\]\[22\] rvcpu.dp.rf.reg_file_arr\[17\]\[22\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[22\] rvcpu.dp.rf.reg_file_arr\[19\]\[22\] _08799_
+ _08800_ VGND VGND VPWR VPWR _09039_ sky130_fd_sc_hd__mux4_1
X_24587_ _10494_ VGND VGND VPWR VPWR _02382_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_182_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_189_5021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29114_ _13072_ VGND VGND VPWR VPWR _04331_ sky130_fd_sc_hd__clkbuf_1
X_26326_ _11078_ _11497_ VGND VGND VPWR VPWR _11498_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_189_5032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23538_ clknet_1_0__leaf__10078_ VGND VGND VPWR VPWR _10172_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_189_5043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29045_ _10066_ _13031_ VGND VGND VPWR VPWR _13036_ sky130_fd_sc_hd__and2_1
XFILLER_0_135_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26257_ _11460_ VGND VGND VPWR VPWR _03086_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16010_ net2674 _13272_ _14333_ VGND VGND VPWR VPWR _14343_ sky130_fd_sc_hd__mux2_1
X_25208_ _10818_ net3086 net56 VGND VGND VPWR VPWR _10843_ sky130_fd_sc_hd__mux2_1
X_26188_ rvcpu.ALUControl\[0\] _11408_ VGND VGND VPWR VPWR _11431_ sky130_fd_sc_hd__and2_1
XFILLER_0_104_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_227_5950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25139_ _10801_ VGND VGND VPWR VPWR _02627_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_148_4050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17961_ _05320_ _05323_ VGND VGND VPWR VPWR _05332_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_223_5836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29947_ net317 _01682_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[15\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_223_5847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_223_5858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19700_ _06777_ _06992_ _06995_ VGND VGND VPWR VPWR _06996_ sky130_fd_sc_hd__or3_1
X_16912_ _04683_ VGND VGND VPWR VPWR _04706_ sky130_fd_sc_hd__buf_4
X_23312__953 clknet_1_1__leaf__10133_ VGND VGND VPWR VPWR net1079 sky130_fd_sc_hd__inv_2
X_17892_ _05264_ VGND VGND VPWR VPWR _05265_ sky130_fd_sc_hd__clkbuf_4
X_29878_ net256 _01613_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[17\]\[9\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_205_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19631_ _06926_ VGND VGND VPWR VPWR _06927_ sky130_fd_sc_hd__clkbuf_4
X_16843_ _04669_ VGND VGND VPWR VPWR _01616_ sky130_fd_sc_hd__clkbuf_1
X_28829_ _12917_ VGND VGND VPWR VPWR _04201_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_219_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31840_ clknet_leaf_158_clk _03294_ VGND VGND VPWR VPWR datamem.data_ram\[8\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_19562_ datamem.data_ram\[3\]\[24\] _06829_ _06854_ _06857_ VGND VGND VPWR VPWR _06858_
+ sky130_fd_sc_hd__o211a_1
X_16774_ net1955 _14461_ _04623_ VGND VGND VPWR VPWR _04633_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_215_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_189_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18513_ _05383_ _05577_ _05581_ VGND VGND VPWR VPWR _05875_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_17_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15725_ _14187_ net3195 _14173_ VGND VGND VPWR VPWR _14188_ sky130_fd_sc_hd__mux2_1
X_19493_ _06655_ VGND VGND VPWR VPWR _06789_ sky130_fd_sc_hd__clkbuf_8
X_31771_ clknet_leaf_235_clk _03225_ VGND VGND VPWR VPWR datamem.data_ram\[1\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_166_clk clknet_5_24__leaf_clk VGND VGND VPWR VPWR clknet_leaf_166_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_17_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18444_ _05799_ _05800_ _05804_ _05806_ VGND VGND VPWR VPWR _05807_ sky130_fd_sc_hd__o211a_1
X_30722_ clknet_leaf_189_clk _02457_ VGND VGND VPWR VPWR datamem.data_ram\[49\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15656_ _13197_ VGND VGND VPWR VPWR _14141_ sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_199_Right_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_174_4666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_4677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14607_ rvcpu.dp.plmw.ALUResultW\[28\] rvcpu.dp.plmw.ReadDataW\[28\] rvcpu.dp.plmw.PCPlus4W\[28\]
+ rvcpu.dp.plmw.lAuiPCW\[28\] _13168_ _13170_ VGND VGND VPWR VPWR _13189_ sky130_fd_sc_hd__mux4_2
XFILLER_0_146_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18375_ _05240_ _05560_ _05739_ VGND VGND VPWR VPWR _05740_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30653_ clknet_leaf_207_clk _02388_ VGND VGND VPWR VPWR datamem.data_ram\[50\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_15587_ net3542 _13207_ _14092_ VGND VGND VPWR VPWR _14101_ sky130_fd_sc_hd__mux2_1
XFILLER_0_200_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_185_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17326_ _04926_ VGND VGND VPWR VPWR _01382_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_172_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30584_ clknet_leaf_188_clk _02319_ VGND VGND VPWR VPWR datamem.data_ram\[53\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_32323_ clknet_leaf_170_clk _03745_ VGND VGND VPWR VPWR datamem.data_ram\[31\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17257_ _04889_ VGND VGND VPWR VPWR _01414_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_77_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16208_ _13234_ VGND VGND VPWR VPWR _14457_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_77_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32254_ clknet_leaf_89_clk _03676_ VGND VGND VPWR VPWR datamem.data_ram\[34\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_133_3684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17188_ _14175_ net4037 _04851_ VGND VGND VPWR VPWR _04853_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_3695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31205_ clknet_leaf_31_clk _02908_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCPlus4D\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16139_ _14412_ VGND VGND VPWR VPWR _01955_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32185_ clknet_leaf_241_clk _03607_ VGND VGND VPWR VPWR datamem.data_ram\[37\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold3206 datamem.data_ram\[55\]\[13\] VGND VGND VPWR VPWR net4356 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold3217 rvcpu.dp.rf.reg_file_arr\[22\]\[14\] VGND VGND VPWR VPWR net4367 sky130_fd_sc_hd__dlygate4sd3_1
X_31136_ clknet_leaf_214_clk _02871_ VGND VGND VPWR VPWR datamem.data_ram\[4\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3228 datamem.data_ram\[53\]\[11\] VGND VGND VPWR VPWR net4378 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold3239 datamem.data_ram\[52\]\[15\] VGND VGND VPWR VPWR net4389 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_102_Left_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2505 rvcpu.dp.rf.reg_file_arr\[9\]\[1\] VGND VGND VPWR VPWR net3655 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2516 datamem.data_ram\[50\]\[20\] VGND VGND VPWR VPWR net3666 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_36_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2527 rvcpu.dp.rf.reg_file_arr\[25\]\[14\] VGND VGND VPWR VPWR net3677 sky130_fd_sc_hd__dlygate4sd3_1
X_31067_ clknet_leaf_279_clk _02802_ VGND VGND VPWR VPWR datamem.data_ram\[8\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2538 rvcpu.dp.rf.reg_file_arr\[12\]\[14\] VGND VGND VPWR VPWR net3688 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1804 datamem.data_ram\[17\]\[22\] VGND VGND VPWR VPWR net2954 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_166_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_3909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2549 rvcpu.dp.rf.reg_file_arr\[26\]\[1\] VGND VGND VPWR VPWR net3699 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1815 rvcpu.dp.rf.reg_file_arr\[15\]\[5\] VGND VGND VPWR VPWR net2965 sky130_fd_sc_hd__dlygate4sd3_1
X_30018_ net380 _01753_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[13\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_23287__930 clknet_1_0__leaf__10131_ VGND VGND VPWR VPWR net1056 sky130_fd_sc_hd__inv_2
XFILLER_0_208_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19829_ datamem.data_ram\[32\]\[1\] _07122_ _07123_ datamem.data_ram\[36\]\[1\] VGND
+ VGND VPWR VPWR _07124_ sky130_fd_sc_hd__a22o_1
Xhold1826 datamem.data_ram\[2\]\[12\] VGND VGND VPWR VPWR net2976 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1837 rvcpu.dp.rf.reg_file_arr\[12\]\[12\] VGND VGND VPWR VPWR net2987 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1848 datamem.data_ram\[25\]\[24\] VGND VGND VPWR VPWR net2998 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1859 rvcpu.dp.rf.reg_file_arr\[30\]\[28\] VGND VGND VPWR VPWR net3009 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22840_ _09413_ _09977_ VGND VGND VPWR VPWR _09978_ sky130_fd_sc_hd__nor2_1
XFILLER_0_194_1192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_157_clk clknet_5_27__leaf_clk VGND VGND VPWR VPWR clknet_leaf_157_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_17_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22771_ _09429_ _09910_ _09912_ VGND VGND VPWR VPWR _09913_ sky130_fd_sc_hd__a21o_1
XFILLER_0_91_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31969_ clknet_leaf_130_clk _03391_ VGND VGND VPWR VPWR datamem.data_ram\[54\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24510_ _09247_ VGND VGND VPWR VPWR _10448_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_101_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21722_ _08842_ _08966_ VGND VGND VPWR VPWR _08967_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25490_ _10811_ net3828 _10999_ VGND VGND VPWR VPWR _11000_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_101_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_166_Right_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_74_Right_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_111_Left_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24441_ _10405_ _10406_ VGND VGND VPWR VPWR _10407_ sky130_fd_sc_hd__and2_1
XFILLER_0_176_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21653_ _08673_ _08900_ VGND VGND VPWR VPWR _08901_ sky130_fd_sc_hd__or2_1
XFILLER_0_136_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27160_ _11968_ _11984_ VGND VGND VPWR VPWR _11986_ sky130_fd_sc_hd__and2_1
X_20604_ datamem.data_ram\[56\]\[13\] _06837_ _06657_ datamem.data_ram\[57\]\[13\]
+ _07894_ VGND VGND VPWR VPWR _07895_ sky130_fd_sc_hd__o221a_1
X_24372_ _09326_ net4285 net61 VGND VGND VPWR VPWR _10364_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21584_ rvcpu.dp.rf.reg_file_arr\[0\]\[10\] rvcpu.dp.rf.reg_file_arr\[1\]\[10\] rvcpu.dp.rf.reg_file_arr\[2\]\[10\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[10\] _08550_ _08528_ VGND VGND VPWR VPWR _08836_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_90_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26111_ net1736 _11386_ VGND VGND VPWR VPWR _11391_ sky130_fd_sc_hd__and2_1
X_20535_ _07825_ VGND VGND VPWR VPWR _07826_ sky130_fd_sc_hd__buf_6
X_27091_ _11822_ _11941_ VGND VGND VPWR VPWR _11942_ sky130_fd_sc_hd__and2_1
XFILLER_0_144_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23490__136 clknet_1_0__leaf__10160_ VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__inv_2
XFILLER_0_127_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26042_ _11064_ _11340_ VGND VGND VPWR VPWR _11348_ sky130_fd_sc_hd__and2_1
X_20466_ _07752_ _07757_ _06796_ VGND VGND VPWR VPWR _07758_ sky130_fd_sc_hd__o21a_1
XFILLER_0_132_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22205_ _09375_ VGND VGND VPWR VPWR _01119_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23570__193 clknet_1_0__leaf__10175_ VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__inv_2
X_20397_ _07031_ _07681_ _07683_ _07688_ VGND VGND VPWR VPWR _07689_ sky130_fd_sc_hd__a31o_1
XFILLER_0_101_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_120_Left_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_83_Right_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22136_ _09337_ VGND VGND VPWR VPWR _01088_ sky130_fd_sc_hd__clkbuf_1
X_29801_ clknet_leaf_218_clk _01536_ VGND VGND VPWR VPWR datamem.data_ram\[59\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_27993_ _09281_ VGND VGND VPWR VPWR _12456_ sky130_fd_sc_hd__buf_2
XFILLER_0_218_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23908__465 clknet_1_1__leaf__10225_ VGND VGND VPWR VPWR net591 sky130_fd_sc_hd__inv_2
X_26944_ _11852_ VGND VGND VPWR VPWR _11853_ sky130_fd_sc_hd__buf_2
X_22067_ rvcpu.dp.plem.WriteDataM\[5\] _09264_ _09265_ rvcpu.dp.plem.WriteDataM\[13\]
+ VGND VGND VPWR VPWR _09284_ sky130_fd_sc_hd__a22o_4
X_29732_ net1078 _01467_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[22\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21018_ datamem.data_ram\[48\]\[31\] _06643_ _08306_ _06940_ VGND VGND VPWR VPWR
+ _08307_ sky130_fd_sc_hd__o22a_1
X_29663_ net1009 _01398_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[24\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_26875_ _11725_ _11075_ VGND VGND VPWR VPWR _11808_ sky130_fd_sc_hd__or2_1
XFILLER_0_215_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23607__226 clknet_1_1__leaf__10179_ VGND VGND VPWR VPWR net352 sky130_fd_sc_hd__inv_2
XFILLER_0_215_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28614_ _12700_ net3263 _12796_ VGND VGND VPWR VPWR _12803_ sky130_fd_sc_hd__mux2_1
X_25826_ _11212_ VGND VGND VPWR VPWR _02903_ sky130_fd_sc_hd__clkbuf_1
X_29594_ net948 _01329_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[26\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28545_ _12765_ VGND VGND VPWR VPWR _04069_ sky130_fd_sc_hd__clkbuf_1
X_25757_ _13823_ _13876_ VGND VGND VPWR VPWR _11159_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_148_clk clknet_5_29__leaf_clk VGND VGND VPWR VPWR clknet_leaf_148_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_35_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15510_ _13542_ _13622_ VGND VGND VPWR VPWR _14037_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_92_Right_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24708_ _10465_ net4031 net59 VGND VGND VPWR VPWR _10562_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_179_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16490_ _04482_ VGND VGND VPWR VPWR _01798_ sky130_fd_sc_hd__clkbuf_1
X_28476_ _12720_ VGND VGND VPWR VPWR _04045_ sky130_fd_sc_hd__clkbuf_1
X_25688_ _11083_ _11113_ VGND VGND VPWR VPWR _11116_ sky130_fd_sc_hd__and2_1
XFILLER_0_35_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15441_ _13573_ _13970_ _13971_ _13475_ _13368_ VGND VGND VPWR VPWR _13972_ sky130_fd_sc_hd__o221a_1
X_27427_ _12136_ net3903 _12126_ VGND VGND VPWR VPWR _12137_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_133_Right_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_216_5673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24639_ _10523_ VGND VGND VPWR VPWR _02405_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_216_5684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18160_ _05454_ _05482_ _05514_ _05524_ VGND VGND VPWR VPWR _05525_ sky130_fd_sc_hd__a31o_2
X_15372_ _13694_ _13656_ _13865_ VGND VGND VPWR VPWR _13906_ sky130_fd_sc_hd__or3_1
X_27358_ _10520_ _10997_ _11713_ VGND VGND VPWR VPWR _12097_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_142_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17111_ _14166_ net2712 _04804_ VGND VGND VPWR VPWR _04812_ sky130_fd_sc_hd__mux2_1
X_26309_ _11487_ VGND VGND VPWR VPWR _03111_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18091_ _05456_ _05457_ VGND VGND VPWR VPWR _05459_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27289_ _12036_ net1600 _12053_ _12057_ VGND VGND VPWR VPWR _03521_ sky130_fd_sc_hd__a31o_1
XFILLER_0_151_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17042_ _04775_ VGND VGND VPWR VPWR _01515_ sky130_fd_sc_hd__clkbuf_1
X_29028_ _12745_ net4240 _13020_ VGND VGND VPWR VPWR _13026_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_146_4009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_1211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_4492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18993_ _05713_ _05708_ _05768_ VGND VGND VPWR VPWR _06328_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17944_ _05313_ _05314_ VGND VGND VPWR VPWR _05316_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_218_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17875_ rvcpu.dp.plde.Rs1E\[3\] VGND VGND VPWR VPWR _05248_ sky130_fd_sc_hd__inv_2
X_32941_ clknet_leaf_152_clk _04363_ VGND VGND VPWR VPWR datamem.data_ram\[6\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_105_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_105_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19614_ _06862_ _06909_ _06586_ VGND VGND VPWR VPWR _06910_ sky130_fd_sc_hd__mux2_1
XFILLER_0_219_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16826_ net2077 _14445_ _04659_ VGND VGND VPWR VPWR _04661_ sky130_fd_sc_hd__mux2_1
X_32872_ clknet_leaf_281_clk _04294_ VGND VGND VPWR VPWR datamem.data_ram\[11\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_191_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_205_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_176_4717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31823_ clknet_leaf_105_clk _03277_ VGND VGND VPWR VPWR datamem.data_ram\[16\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_176_4728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16757_ _04624_ VGND VGND VPWR VPWR _01665_ sky130_fd_sc_hd__clkbuf_1
X_19545_ datamem.data_ram\[25\]\[24\] _06790_ _06840_ _06810_ VGND VGND VPWR VPWR
+ _06841_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_139_clk clknet_5_31__leaf_clk VGND VGND VPWR VPWR clknet_leaf_139_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_66_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15708_ _14176_ VGND VGND VPWR VPWR _02166_ sky130_fd_sc_hd__clkbuf_1
X_31754_ clknet_leaf_58_clk _03208_ VGND VGND VPWR VPWR datamem.data_ram\[45\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_66_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19476_ datamem.data_ram\[51\]\[16\] _06739_ _06762_ _06771_ VGND VGND VPWR VPWR
+ _06772_ sky130_fd_sc_hd__o211a_1
X_16688_ _14151_ net2471 _04587_ VGND VGND VPWR VPWR _04588_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30705_ clknet_leaf_219_clk _02440_ VGND VGND VPWR VPWR datamem.data_ram\[49\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18427_ _05576_ _05771_ VGND VGND VPWR VPWR _05791_ sky130_fd_sc_hd__nand2_1
X_15639_ _13174_ rvcpu.dp.plmw.RdW\[3\] _13176_ VGND VGND VPWR VPWR _14129_ sky130_fd_sc_hd__and3_2
XPHY_EDGE_ROW_100_Right_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31685_ clknet_leaf_38_clk _03143_ VGND VGND VPWR VPWR rvcpu.dp.pcreg.q\[3\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_158_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_963 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24033__564 clknet_1_0__leaf__10243_ VGND VGND VPWR VPWR net690 sky130_fd_sc_hd__inv_2
XFILLER_0_185_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18358_ rvcpu.dp.plde.ALUControlE\[0\] rvcpu.dp.plde.ALUControlE\[2\] rvcpu.dp.plde.ALUControlE\[3\]
+ VGND VGND VPWR VPWR _05723_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_135_3724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30636_ clknet_leaf_198_clk _02371_ VGND VGND VPWR VPWR datamem.data_ram\[51\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_135_3735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_3746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17309_ _04917_ VGND VGND VPWR VPWR _01390_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18289_ _05653_ VGND VGND VPWR VPWR _05654_ sky130_fd_sc_hd__buf_2
X_30567_ clknet_leaf_147_clk _02302_ VGND VGND VPWR VPWR datamem.data_ram\[54\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_25_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20320_ datamem.data_ram\[26\]\[4\] _06989_ _06921_ datamem.data_ram\[29\]\[4\] VGND
+ VGND VPWR VPWR _07612_ sky130_fd_sc_hd__a22o_1
XFILLER_0_160_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32306_ clknet_leaf_273_clk _03728_ VGND VGND VPWR VPWR datamem.data_ram\[32\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_22996__702 clknet_1_1__leaf__10084_ VGND VGND VPWR VPWR net828 sky130_fd_sc_hd__inv_2
XFILLER_0_86_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30498_ clknet_leaf_140_clk _02233_ VGND VGND VPWR VPWR datamem.data_ram\[57\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_23319__959 clknet_1_0__leaf__10134_ VGND VGND VPWR VPWR net1085 sky130_fd_sc_hd__inv_2
XFILLER_0_86_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold901 rvcpu.dp.rf.reg_file_arr\[30\]\[17\] VGND VGND VPWR VPWR net2051 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold912 rvcpu.dp.pcreg.q\[14\] VGND VGND VPWR VPWR net2062 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20251_ _06967_ _07541_ _07543_ VGND VGND VPWR VPWR _07544_ sky130_fd_sc_hd__or3_1
XFILLER_0_114_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold923 rvcpu.dp.rf.reg_file_arr\[16\]\[7\] VGND VGND VPWR VPWR net2073 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32237_ clknet_leaf_242_clk _03659_ VGND VGND VPWR VPWR datamem.data_ram\[35\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_38_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold934 datamem.data_ram\[33\]\[14\] VGND VGND VPWR VPWR net2084 sky130_fd_sc_hd__dlygate4sd3_1
Xhold945 datamem.data_ram\[42\]\[14\] VGND VGND VPWR VPWR net2095 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold956 rvcpu.dp.rf.reg_file_arr\[5\]\[17\] VGND VGND VPWR VPWR net2106 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold967 datamem.data_ram\[43\]\[14\] VGND VGND VPWR VPWR net2117 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3003 rvcpu.dp.rf.reg_file_arr\[13\]\[23\] VGND VGND VPWR VPWR net4153 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20182_ datamem.data_ram\[10\]\[11\] _06692_ _07473_ _07474_ VGND VGND VPWR VPWR
+ _07475_ sky130_fd_sc_hd__o211a_1
X_32168_ clknet_leaf_277_clk _03590_ VGND VGND VPWR VPWR datamem.data_ram\[38\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold978 rvcpu.dp.rf.reg_file_arr\[27\]\[1\] VGND VGND VPWR VPWR net2128 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3014 datamem.data_ram\[0\]\[23\] VGND VGND VPWR VPWR net4164 sky130_fd_sc_hd__dlygate4sd3_1
Xhold989 datamem.data_ram\[33\]\[31\] VGND VGND VPWR VPWR net2139 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3025 datamem.data_ram\[18\]\[17\] VGND VGND VPWR VPWR net4175 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3036 datamem.data_ram\[15\]\[10\] VGND VGND VPWR VPWR net4186 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_228_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31119_ clknet_leaf_110_clk _02854_ VGND VGND VPWR VPWR datamem.data_ram\[35\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_196_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2302 datamem.data_ram\[36\]\[25\] VGND VGND VPWR VPWR net3452 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3047 datamem.data_ram\[48\]\[29\] VGND VGND VPWR VPWR net4197 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32099_ clknet_leaf_107_clk _03521_ VGND VGND VPWR VPWR datamem.data_ram\[23\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2313 datamem.data_ram\[53\]\[22\] VGND VGND VPWR VPWR net3463 sky130_fd_sc_hd__dlygate4sd3_1
X_24990_ _10439_ net3291 _10715_ VGND VGND VPWR VPWR _10716_ sky130_fd_sc_hd__mux2_1
Xhold3058 rvcpu.dp.rf.reg_file_arr\[14\]\[16\] VGND VGND VPWR VPWR net4208 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3069 rvcpu.dp.rf.reg_file_arr\[25\]\[25\] VGND VGND VPWR VPWR net4219 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2324 rvcpu.dp.rf.reg_file_arr\[12\]\[18\] VGND VGND VPWR VPWR net3474 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2335 datamem.data_ram\[28\]\[11\] VGND VGND VPWR VPWR net3485 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1601 datamem.data_ram\[15\]\[26\] VGND VGND VPWR VPWR net2751 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2346 rvcpu.dp.rf.reg_file_arr\[28\]\[9\] VGND VGND VPWR VPWR net3496 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2357 datamem.data_ram\[4\]\[11\] VGND VGND VPWR VPWR net3507 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1612 datamem.data_ram\[7\]\[26\] VGND VGND VPWR VPWR net2762 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1623 datamem.data_ram\[45\]\[22\] VGND VGND VPWR VPWR net2773 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2368 rvcpu.dp.rf.reg_file_arr\[21\]\[3\] VGND VGND VPWR VPWR net3518 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2379 datamem.data_ram\[22\]\[17\] VGND VGND VPWR VPWR net3529 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1634 rvcpu.dp.rf.reg_file_arr\[23\]\[2\] VGND VGND VPWR VPWR net2784 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1645 datamem.data_ram\[36\]\[21\] VGND VGND VPWR VPWR net2795 sky130_fd_sc_hd__dlygate4sd3_1
X_26660_ _11679_ _11677_ VGND VGND VPWR VPWR _11680_ sky130_fd_sc_hd__and2_1
Xhold1656 rvcpu.dp.rf.reg_file_arr\[13\]\[27\] VGND VGND VPWR VPWR net2806 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1667 datamem.data_ram\[16\]\[19\] VGND VGND VPWR VPWR net2817 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1678 datamem.data_ram\[9\]\[21\] VGND VGND VPWR VPWR net2828 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1689 rvcpu.dp.rf.reg_file_arr\[20\]\[21\] VGND VGND VPWR VPWR net2839 sky130_fd_sc_hd__dlygate4sd3_1
X_25611_ _10731_ net3048 net53 VGND VGND VPWR VPWR _11070_ sky130_fd_sc_hd__mux2_1
Xclkbuf_0__10260_ _10260_ VGND VGND VPWR VPWR clknet_0__10260_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_169_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__10160_ clknet_0__10160_ VGND VGND VPWR VPWR clknet_1_1__leaf__10160_
+ sky130_fd_sc_hd__clkbuf_16
X_22823_ rvcpu.dp.rf.reg_file_arr\[4\]\[27\] rvcpu.dp.rf.reg_file_arr\[5\]\[27\] rvcpu.dp.rf.reg_file_arr\[6\]\[27\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[27\] _09416_ _09716_ VGND VGND VPWR VPWR _09962_
+ sky130_fd_sc_hd__mux4_1
X_26591_ _11618_ net1701 _11639_ _11642_ VGND VGND VPWR VPWR _03238_ sky130_fd_sc_hd__a31o_1
XFILLER_0_17_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28330_ _12369_ net2909 _12632_ VGND VGND VPWR VPWR _12639_ sky130_fd_sc_hd__mux2_1
X_25542_ _10739_ net3613 _11021_ VGND VGND VPWR VPWR _11029_ sky130_fd_sc_hd__mux2_1
Xclkbuf_0__10191_ _10191_ VGND VGND VPWR VPWR clknet_0__10191_ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_1__f__10091_ clknet_0__10091_ VGND VGND VPWR VPWR clknet_1_1__leaf__10091_
+ sky130_fd_sc_hd__clkbuf_16
X_22754_ rvcpu.dp.rf.reg_file_arr\[8\]\[23\] rvcpu.dp.rf.reg_file_arr\[10\]\[23\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[23\] rvcpu.dp.rf.reg_file_arr\[11\]\[23\] _09483_
+ _09656_ VGND VGND VPWR VPWR _09897_ sky130_fd_sc_hd__mux4_1
XFILLER_0_17_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21705_ _08565_ _08948_ _08950_ _08576_ VGND VGND VPWR VPWR _08951_ sky130_fd_sc_hd__o211a_1
X_28261_ _12600_ VGND VGND VPWR VPWR _03950_ sky130_fd_sc_hd__clkbuf_1
X_25473_ _10418_ _10985_ VGND VGND VPWR VPWR _10993_ sky130_fd_sc_hd__and2_1
X_22685_ _09831_ VGND VGND VPWR VPWR _01143_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_212_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27212_ _11980_ _12008_ VGND VGND VPWR VPWR _12016_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24424_ _09281_ VGND VGND VPWR VPWR _10394_ sky130_fd_sc_hd__buf_2
XFILLER_0_212_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28192_ _12563_ VGND VGND VPWR VPWR _03918_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_922 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21636_ _08798_ _08884_ VGND VGND VPWR VPWR _08885_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_229_6009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27143_ _11918_ VGND VGND VPWR VPWR _11974_ sky130_fd_sc_hd__buf_2
X_24355_ _09288_ net3578 _10348_ VGND VGND VPWR VPWR _10355_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_211_5570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21567_ rvcpu.dp.rf.reg_file_arr\[12\]\[9\] rvcpu.dp.rf.reg_file_arr\[13\]\[9\] rvcpu.dp.rf.reg_file_arr\[14\]\[9\]
+ rvcpu.dp.rf.reg_file_arr\[15\]\[9\] _08696_ _08568_ VGND VGND VPWR VPWR _08820_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_35_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27074_ _11833_ _11924_ VGND VGND VPWR VPWR _11930_ sky130_fd_sc_hd__and2_1
X_20518_ datamem.data_ram\[30\]\[21\] _07028_ _07808_ datamem.data_ram\[25\]\[21\]
+ VGND VGND VPWR VPWR _07809_ sky130_fd_sc_hd__o22a_1
X_24286_ _10297_ _09269_ _10269_ VGND VGND VPWR VPWR _10316_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_16_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21498_ _08542_ _08753_ VGND VGND VPWR VPWR _08754_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26025_ _11109_ _10980_ VGND VGND VPWR VPWR _11338_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20449_ datamem.data_ram\[3\]\[20\] _06738_ _06700_ datamem.data_ram\[1\]\[20\] _07740_
+ VGND VGND VPWR VPWR _07741_ sky130_fd_sc_hd__o221a_1
XFILLER_0_127_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22119_ _09326_ net3380 _09302_ VGND VGND VPWR VPWR _09327_ sky130_fd_sc_hd__mux2_1
X_27976_ _12444_ VGND VGND VPWR VPWR _03821_ sky130_fd_sc_hd__clkbuf_1
X_15990_ _14332_ VGND VGND VPWR VPWR _02032_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_206_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14941_ _13488_ _13489_ VGND VGND VPWR VPWR _13490_ sky130_fd_sc_hd__nor2_1
X_26927_ _11831_ net1529 _11841_ _11843_ VGND VGND VPWR VPWR _03373_ sky130_fd_sc_hd__a31o_1
X_29715_ net1061 _01450_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[22\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_202_Right_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_215_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2880 rvcpu.dp.rf.reg_file_arr\[26\]\[6\] VGND VGND VPWR VPWR net4030 sky130_fd_sc_hd__dlygate4sd3_1
X_17660_ net3633 _13240_ _05093_ VGND VGND VPWR VPWR _05103_ sky130_fd_sc_hd__mux2_1
X_26858_ _11676_ _11798_ VGND VGND VPWR VPWR _11799_ sky130_fd_sc_hd__and2_1
X_14872_ _13281_ _13414_ VGND VGND VPWR VPWR _13424_ sky130_fd_sc_hd__nor2_1
X_29646_ net992 _01381_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[24\]\[9\] sky130_fd_sc_hd__dfxtp_1
Xhold2891 datamem.data_ram\[46\]\[8\] VGND VGND VPWR VPWR net4041 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_214_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16611_ _14143_ net3446 _04540_ VGND VGND VPWR VPWR _04547_ sky130_fd_sc_hd__mux2_1
XFILLER_0_203_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25809_ _11197_ _11198_ _11149_ VGND VGND VPWR VPWR _11199_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_218_5724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17591_ _05066_ VGND VGND VPWR VPWR _01241_ sky130_fd_sc_hd__clkbuf_1
X_29577_ net931 _01312_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[26\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26789_ _11687_ _11749_ VGND VGND VPWR VPWR _11757_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_207_Left_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_218_5735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28528_ _09235_ VGND VGND VPWR VPWR _12754_ sky130_fd_sc_hd__buf_2
X_19330_ _06625_ VGND VGND VPWR VPWR _06626_ sky130_fd_sc_hd__clkbuf_8
X_16542_ _14143_ net3757 _04503_ VGND VGND VPWR VPWR _04510_ sky130_fd_sc_hd__mux2_1
XFILLER_0_211_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_171_4603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19261_ _06562_ rvcpu.dp.plde.ImmExtE\[31\] rvcpu.dp.plde.luiE VGND VGND VPWR VPWR
+ _06563_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28459_ _12711_ VGND VGND VPWR VPWR _04037_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16473_ _04473_ VGND VGND VPWR VPWR _01806_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18212_ _05575_ _05389_ _05576_ _05394_ VGND VGND VPWR VPWR _05577_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15424_ _13368_ _13948_ _13952_ _13955_ VGND VGND VPWR VPWR _13956_ sky130_fd_sc_hd__a211o_1
XFILLER_0_38_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19192_ _06501_ _06502_ VGND VGND VPWR VPWR _06503_ sky130_fd_sc_hd__nand2_1
X_31470_ clknet_leaf_7_clk rvcpu.dp.SrcBFW_Mux.y\[28\] VGND VGND VPWR VPWR rvcpu.dp.plem.WriteDataM\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23577__199 clknet_1_1__leaf__10176_ VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__inv_2
XFILLER_0_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18143_ _05508_ VGND VGND VPWR VPWR rvcpu.dp.SrcBFW_Mux.y\[16\] sky130_fd_sc_hd__buf_1
XFILLER_0_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30421_ net759 _02156_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[29\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15355_ _13665_ _13668_ _13610_ VGND VGND VPWR VPWR _13890_ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18074_ _05441_ _05430_ VGND VGND VPWR VPWR _05442_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_3610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_854 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30352_ net698 _02087_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[3\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_15286_ _13392_ _13523_ VGND VGND VPWR VPWR _13824_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_130_3621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_216_Left_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_169_4543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold208 datamem.data_ram\[40\]\[1\] VGND VGND VPWR VPWR net1358 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_169_4554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__10180_ clknet_0__10180_ VGND VGND VPWR VPWR clknet_1_0__leaf__10180_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_41_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold219 datamem.data_ram\[7\]\[7\] VGND VGND VPWR VPWR net1369 sky130_fd_sc_hd__dlygate4sd3_1
X_17025_ _04766_ VGND VGND VPWR VPWR _01523_ sky130_fd_sc_hd__clkbuf_1
X_30283_ clknet_leaf_140_clk _02018_ VGND VGND VPWR VPWR datamem.data_ram\[58\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32022_ clknet_leaf_129_clk _03444_ VGND VGND VPWR VPWR datamem.data_ram\[51\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18976_ _06202_ _06311_ _05698_ VGND VGND VPWR VPWR _06312_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_128_3561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17927_ rvcpu.dp.plde.RD1E\[28\] _05291_ _05294_ _13189_ _05299_ VGND VGND VPWR VPWR
+ _05300_ sky130_fd_sc_hd__o221a_2
XTAP_TAPCELL_ROW_128_3572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32924_ clknet_leaf_258_clk _04346_ VGND VGND VPWR VPWR datamem.data_ram\[0\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_17858_ _05233_ VGND VGND VPWR VPWR rvcpu.dp.SrcBFW_Mux.y\[7\] sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_225_Left_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_124_3469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16809_ net1908 _14428_ _04648_ VGND VGND VPWR VPWR _04652_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32855_ clknet_leaf_185_clk _04277_ VGND VGND VPWR VPWR datamem.data_ram\[11\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17789_ net122 VGND VGND VPWR VPWR _05185_ sky130_fd_sc_hd__inv_2
XFILLER_0_191_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31806_ clknet_leaf_73_clk _03260_ VGND VGND VPWR VPWR datamem.data_ram\[46\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19528_ datamem.data_ram\[42\]\[24\] _06802_ _06669_ datamem.data_ram\[47\]\[24\]
+ VGND VGND VPWR VPWR _06824_ sky130_fd_sc_hd__o22a_1
XFILLER_0_49_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_5_22__f_clk clknet_2_2_0_clk VGND VGND VPWR VPWR clknet_5_22__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_113_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32786_ clknet_leaf_259_clk _04208_ VGND VGND VPWR VPWR datamem.data_ram\[14\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19459_ datamem.data_ram\[58\]\[16\] _06754_ _06671_ datamem.data_ram\[63\]\[16\]
+ VGND VGND VPWR VPWR _06755_ sky130_fd_sc_hd__o22a_1
XFILLER_0_118_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31737_ net186 _03195_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[9\]\[23\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_27_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22470_ rvcpu.dp.rf.reg_file_arr\[8\]\[8\] rvcpu.dp.rf.reg_file_arr\[10\]\[8\] rvcpu.dp.rf.reg_file_arr\[9\]\[8\]
+ rvcpu.dp.rf.reg_file_arr\[11\]\[8\] _09608_ _09532_ VGND VGND VPWR VPWR _09628_
+ sky130_fd_sc_hd__mux4_1
X_31668_ clknet_leaf_47_clk net1298 VGND VGND VPWR VPWR rvcpu.dp.plmw.ALUResultW\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21421_ _08678_ _08679_ _08514_ VGND VGND VPWR VPWR _08680_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_98_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30619_ clknet_leaf_136_clk _02354_ VGND VGND VPWR VPWR datamem.data_ram\[52\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31599_ clknet_leaf_47_clk net1229 VGND VGND VPWR VPWR rvcpu.dp.plmw.PCPlus4W\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21352_ rvcpu.dp.plde.funct3E\[0\] rvcpu.dp.plde.funct3E\[1\] rvcpu.ALUResultE\[31\]
+ rvcpu.dp.plde.funct3E\[2\] VGND VGND VPWR VPWR _08614_ sky130_fd_sc_hd__or4bb_1
X_24140_ clknet_1_0__leaf__10244_ VGND VGND VPWR VPWR _10262_ sky130_fd_sc_hd__buf_1
XFILLER_0_86_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20303_ _06916_ _07579_ _07584_ _07595_ _06985_ VGND VGND VPWR VPWR _07596_ sky130_fd_sc_hd__o311a_1
XFILLER_0_130_824 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21283_ _08513_ _08521_ _08530_ _08539_ _08544_ VGND VGND VPWR VPWR _08545_ sky130_fd_sc_hd__o32a_1
Xhold720 datamem.data_ram\[52\]\[6\] VGND VGND VPWR VPWR net1870 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold731 rvcpu.dp.rf.reg_file_arr\[6\]\[12\] VGND VGND VPWR VPWR net1881 sky130_fd_sc_hd__dlygate4sd3_1
Xhold742 rvcpu.dp.plfd.PCPlus4D\[25\] VGND VGND VPWR VPWR net1892 sky130_fd_sc_hd__dlygate4sd3_1
X_20234_ datamem.data_ram\[2\]\[3\] _07000_ _07523_ _07526_ VGND VGND VPWR VPWR _07527_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_188_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold753 datamem.data_ram\[46\]\[14\] VGND VGND VPWR VPWR net1903 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23022_ clknet_1_0__leaf__10087_ VGND VGND VPWR VPWR _10088_ sky130_fd_sc_hd__buf_1
XFILLER_0_40_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_57_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold764 rvcpu.dp.rf.reg_file_arr\[6\]\[30\] VGND VGND VPWR VPWR net1914 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold775 datamem.data_ram\[36\]\[22\] VGND VGND VPWR VPWR net1925 sky130_fd_sc_hd__dlygate4sd3_1
Xhold786 datamem.data_ram\[32\]\[23\] VGND VGND VPWR VPWR net1936 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27830_ _12359_ net3505 _12357_ VGND VGND VPWR VPWR _12360_ sky130_fd_sc_hd__mux2_1
Xhold797 rvcpu.dp.rf.reg_file_arr\[7\]\[30\] VGND VGND VPWR VPWR net1947 sky130_fd_sc_hd__dlygate4sd3_1
X_20165_ datamem.data_ram\[17\]\[27\] _06657_ _07454_ _07457_ VGND VGND VPWR VPWR
+ _07458_ sky130_fd_sc_hd__o211a_1
XFILLER_0_228_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2110 datamem.data_ram\[44\]\[25\] VGND VGND VPWR VPWR net3260 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_200_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2121 datamem.data_ram\[57\]\[12\] VGND VGND VPWR VPWR net3271 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2132 rvcpu.dp.rf.reg_file_arr\[21\]\[5\] VGND VGND VPWR VPWR net3282 sky130_fd_sc_hd__dlygate4sd3_1
X_27761_ _12320_ VGND VGND VPWR VPWR _03730_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24973_ _10465_ net3839 net101 VGND VGND VPWR VPWR _10707_ sky130_fd_sc_hd__mux2_1
X_20096_ _06715_ _07378_ _07389_ _06712_ VGND VGND VPWR VPWR _07390_ sky130_fd_sc_hd__o211a_1
Xhold2143 datamem.data_ram\[48\]\[12\] VGND VGND VPWR VPWR net3293 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2154 datamem.data_ram\[30\]\[26\] VGND VGND VPWR VPWR net3304 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2165 datamem.data_ram\[1\]\[20\] VGND VGND VPWR VPWR net3315 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1420 datamem.data_ram\[33\]\[20\] VGND VGND VPWR VPWR net2570 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2176 datamem.data_ram\[35\]\[10\] VGND VGND VPWR VPWR net3326 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1431 datamem.data_ram\[7\]\[11\] VGND VGND VPWR VPWR net2581 sky130_fd_sc_hd__dlygate4sd3_1
X_26712_ _10824_ net3503 _11704_ VGND VGND VPWR VPWR _11711_ sky130_fd_sc_hd__mux2_1
X_29500_ net862 _01235_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[28\]\[7\] sky130_fd_sc_hd__dfxtp_1
Xhold1442 rvcpu.dp.rf.reg_file_arr\[7\]\[26\] VGND VGND VPWR VPWR net2592 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27692_ _12132_ net2486 _12280_ VGND VGND VPWR VPWR _12284_ sky130_fd_sc_hd__mux2_1
Xhold2187 datamem.data_ram\[18\]\[24\] VGND VGND VPWR VPWR net3337 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1453 rvcpu.dp.rf.reg_file_arr\[17\]\[9\] VGND VGND VPWR VPWR net2603 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2198 datamem.data_ram\[62\]\[26\] VGND VGND VPWR VPWR net3348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1464 rvcpu.dp.rf.reg_file_arr\[22\]\[21\] VGND VGND VPWR VPWR net2614 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1475 rvcpu.dp.rf.reg_file_arr\[31\]\[19\] VGND VGND VPWR VPWR net2625 sky130_fd_sc_hd__dlygate4sd3_1
X_29431_ net793 _01166_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[30\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_26643_ _11665_ net1700 _11662_ _11668_ VGND VGND VPWR VPWR _03264_ sky130_fd_sc_hd__a31o_1
XFILLER_0_196_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1486 rvcpu.dp.rf.reg_file_arr\[17\]\[23\] VGND VGND VPWR VPWR net2636 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1497 datamem.data_ram\[30\]\[11\] VGND VGND VPWR VPWR net2647 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_200_5293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__10243_ _10243_ VGND VGND VPWR VPWR clknet_0__10243_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_197_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29362_ clknet_leaf_268_clk _01097_ VGND VGND VPWR VPWR datamem.data_ram\[61\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_22806_ rvcpu.dp.rf.reg_file_arr\[0\]\[26\] rvcpu.dp.rf.reg_file_arr\[1\]\[26\] rvcpu.dp.rf.reg_file_arr\[2\]\[26\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[26\] _09463_ _09637_ VGND VGND VPWR VPWR _09946_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_0_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26574_ _11632_ VGND VGND VPWR VPWR _03231_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_212_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20998_ datamem.data_ram\[24\]\[15\] _06643_ _06616_ datamem.data_ram\[28\]\[15\]
+ _08286_ VGND VGND VPWR VPWR _08287_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_0_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28313_ _12460_ net3276 net72 VGND VGND VPWR VPWR _12630_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25525_ _11018_ net1582 _11009_ _11019_ VGND VGND VPWR VPWR _02795_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_0_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__10174_ _10174_ VGND VGND VPWR VPWR clknet_0__10174_ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_192_5094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29293_ clknet_leaf_0_clk _01028_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD1E\[0\] sky130_fd_sc_hd__dfxtp_1
X_22737_ rvcpu.dp.rf.reg_file_arr\[0\]\[22\] rvcpu.dp.rf.reg_file_arr\[1\]\[22\] rvcpu.dp.rf.reg_file_arr\[2\]\[22\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[22\] _09477_ _09466_ VGND VGND VPWR VPWR _09881_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_213_5610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28244_ _12591_ VGND VGND VPWR VPWR _03942_ sky130_fd_sc_hd__clkbuf_1
X_23496__142 clknet_1_1__leaf__10160_ VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__inv_2
X_25456_ _10783_ _10981_ _10982_ net1294 VGND VGND VPWR VPWR _02763_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_211_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22668_ rvcpu.dp.rf.reg_file_arr\[16\]\[19\] rvcpu.dp.rf.reg_file_arr\[17\]\[19\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[19\] rvcpu.dp.rf.reg_file_arr\[19\]\[19\] _09384_
+ _09430_ VGND VGND VPWR VPWR _09815_ sky130_fd_sc_hd__mux4_1
XFILLER_0_164_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24407_ _09288_ net2658 _10376_ VGND VGND VPWR VPWR _10383_ sky130_fd_sc_hd__mux2_1
X_28175_ _12554_ VGND VGND VPWR VPWR _03910_ sky130_fd_sc_hd__clkbuf_1
X_21619_ _08673_ _08868_ VGND VGND VPWR VPWR _08869_ sky130_fd_sc_hd__or2_1
X_25387_ _10938_ net1378 _10934_ _10945_ VGND VGND VPWR VPWR _02731_ sky130_fd_sc_hd__a31o_1
XFILLER_0_168_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22599_ _09412_ _09745_ _09747_ _09749_ _09413_ VGND VGND VPWR VPWR _09750_ sky130_fd_sc_hd__a221o_1
XFILLER_0_180_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15140_ _13573_ _13472_ _13546_ VGND VGND VPWR VPWR _13684_ sky130_fd_sc_hd__or3_1
X_27126_ _11837_ _11953_ VGND VGND VPWR VPWR _11962_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_11_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24338_ _10345_ VGND VGND VPWR VPWR _02282_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_11_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15071_ _13470_ _13614_ _13616_ VGND VGND VPWR VPWR _13617_ sky130_fd_sc_hd__or3_1
X_27057_ _11835_ _11911_ VGND VGND VPWR VPWR _11920_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_205_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24269_ _10297_ _09229_ _10269_ VGND VGND VPWR VPWR _10307_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_205_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26008_ _11143_ VGND VGND VPWR VPWR _11329_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_207_5458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_207_5469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_4440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18830_ _05990_ _06047_ _06174_ _06109_ _06175_ VGND VGND VPWR VPWR _06176_ sky130_fd_sc_hd__o221a_1
XFILLER_0_219_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_4326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_4337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18761_ _05960_ _06022_ _06110_ VGND VGND VPWR VPWR _06111_ sky130_fd_sc_hd__o21ai_1
X_15973_ net2427 _13217_ _14322_ VGND VGND VPWR VPWR _14324_ sky130_fd_sc_hd__mux2_1
X_27959_ _09235_ VGND VGND VPWR VPWR _12433_ sky130_fd_sc_hd__clkbuf_2
X_14924_ _13402_ _13472_ VGND VGND VPWR VPWR _13473_ sky130_fd_sc_hd__nor2_2
X_17712_ _13217_ net3906 _05129_ VGND VGND VPWR VPWR _05131_ sky130_fd_sc_hd__mux2_1
X_30970_ clknet_leaf_216_clk _02705_ VGND VGND VPWR VPWR datamem.data_ram\[39\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_222_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18692_ _05966_ _06045_ _05705_ VGND VGND VPWR VPWR _06046_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold80 rvcpu.dp.plde.PCPlus4E\[11\] VGND VGND VPWR VPWR net1230 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold91 rvcpu.dp.plem.PCPlus4M\[3\] VGND VGND VPWR VPWR net1241 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14855_ _13341_ _13294_ VGND VGND VPWR VPWR _13407_ sky130_fd_sc_hd__nand2_1
X_29629_ clknet_leaf_142_clk _01364_ VGND VGND VPWR VPWR datamem.data_ram\[5\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_17643_ _05094_ VGND VGND VPWR VPWR _01217_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23348__985 clknet_1_1__leaf__10137_ VGND VGND VPWR VPWR net1111 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_63_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_188_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32640_ clknet_leaf_3_clk _04062_ VGND VGND VPWR VPWR datamem.data_ram\[1\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_17574_ _13213_ net2532 _05057_ VGND VGND VPWR VPWR _05058_ sky130_fd_sc_hd__mux2_1
XFILLER_0_212_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14786_ _13328_ _13330_ _13338_ VGND VGND VPWR VPWR _13339_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_203_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_367 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_4277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_4288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16525_ _04500_ VGND VGND VPWR VPWR _01781_ sky130_fd_sc_hd__clkbuf_1
X_19313_ _06608_ VGND VGND VPWR VPWR _06609_ sky130_fd_sc_hd__buf_6
X_32571_ clknet_leaf_252_clk _03993_ VGND VGND VPWR VPWR datamem.data_ram\[22\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_158_4299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_70_clk clknet_5_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_70_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_133_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31522_ clknet_leaf_47_clk net1224 VGND VGND VPWR VPWR rvcpu.dp.plem.PCPlus4M\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_19244_ rvcpu.dp.plde.ImmExtE\[29\] rvcpu.dp.plde.PCE\[29\] VGND VGND VPWR VPWR _06548_
+ sky130_fd_sc_hd__or2_1
X_16456_ net4258 _14486_ _14560_ VGND VGND VPWR VPWR _04463_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_730 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15407_ _13933_ _13935_ _13938_ _13466_ VGND VGND VPWR VPWR _13939_ sky130_fd_sc_hd__o2bb2a_1
X_19175_ _06486_ _06487_ VGND VGND VPWR VPWR _06488_ sky130_fd_sc_hd__nand2_1
XFILLER_0_171_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31453_ clknet_leaf_5_clk rvcpu.dp.SrcBFW_Mux.y\[11\] VGND VGND VPWR VPWR rvcpu.dp.plem.WriteDataM\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_22_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16387_ _14558_ VGND VGND VPWR VPWR _01845_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18126_ _05492_ VGND VGND VPWR VPWR rvcpu.dp.SrcBFW_Mux.y\[18\] sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_42_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30404_ net742 _02139_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[31\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_15338_ _13696_ _13873_ VGND VGND VPWR VPWR _13874_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31384_ clknet_leaf_39_clk _03087_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCE\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_3295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18057_ _05421_ _05424_ VGND VGND VPWR VPWR _05425_ sky130_fd_sc_hd__and2_1
X_30335_ net681 _02070_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[4\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_15269_ _13463_ _13728_ _13807_ _13428_ _13412_ VGND VGND VPWR VPWR _13808_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_188_4996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17008_ net2549 _14420_ _04757_ VGND VGND VPWR VPWR _04758_ sky130_fd_sc_hd__mux2_1
X_30266_ net620 _02001_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[6\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32005_ clknet_leaf_135_clk _03427_ VGND VGND VPWR VPWR datamem.data_ram\[52\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30197_ net551 _01932_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[8\]\[16\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_126_3509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18959_ _05543_ _06295_ VGND VGND VPWR VPWR _06296_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_207_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_225_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_1246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21970_ _09199_ _09200_ rvcpu.dp.plfd.InstrD\[17\] VGND VGND VPWR VPWR _09201_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20921_ datamem.data_ram\[46\]\[22\] datamem.data_ram\[47\]\[22\] _07829_ VGND VGND
+ VPWR VPWR _08211_ sky130_fd_sc_hd__mux2_1
X_32907_ clknet_leaf_262_clk _04329_ VGND VGND VPWR VPWR datamem.data_ram\[7\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_221_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23640_ _10186_ VGND VGND VPWR VPWR _01743_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_194_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32838_ clknet_leaf_283_clk _04260_ VGND VGND VPWR VPWR datamem.data_ram\[12\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_20852_ _07851_ _08141_ VGND VGND VPWR VPWR _08142_ sky130_fd_sc_hd__or2_1
XFILLER_0_166_507 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_221_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32769_ clknet_leaf_234_clk _04191_ VGND VGND VPWR VPWR datamem.data_ram\[14\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_20783_ datamem.data_ram\[0\]\[30\] _06779_ _06783_ datamem.data_ram\[1\]\[30\] VGND
+ VGND VPWR VPWR _08073_ sky130_fd_sc_hd__o22a_1
XFILLER_0_92_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_193_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_61_clk clknet_5_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_61_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_14_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25310_ _10811_ net3398 _10899_ VGND VGND VPWR VPWR _10900_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22522_ _09495_ _09676_ _09472_ VGND VGND VPWR VPWR _09677_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26290_ _11477_ VGND VGND VPWR VPWR _03102_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_174_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25241_ _10860_ VGND VGND VPWR VPWR _02670_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22453_ _09429_ _09609_ _09611_ _09438_ VGND VGND VPWR VPWR _09612_ sky130_fd_sc_hd__a211o_1
XFILLER_0_88_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21404_ rvcpu.dp.rf.reg_file_arr\[12\]\[2\] rvcpu.dp.rf.reg_file_arr\[13\]\[2\] rvcpu.dp.rf.reg_file_arr\[14\]\[2\]
+ rvcpu.dp.rf.reg_file_arr\[15\]\[2\] _08551_ _08555_ VGND VGND VPWR VPWR _08664_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_32_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25172_ _10821_ VGND VGND VPWR VPWR _02640_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_59_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22384_ _09540_ _09542_ _09545_ _09412_ _09413_ VGND VGND VPWR VPWR _09546_ sky130_fd_sc_hd__a221o_1
XFILLER_0_161_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21335_ _08591_ _08594_ _08596_ VGND VGND VPWR VPWR _08597_ sky130_fd_sc_hd__and3b_2
XFILLER_0_163_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29980_ net350 _01715_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[14\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28931_ _12971_ VGND VGND VPWR VPWR _04249_ sky130_fd_sc_hd__clkbuf_1
Xhold550 datamem.data_ram\[17\]\[3\] VGND VGND VPWR VPWR net1700 sky130_fd_sc_hd__dlygate4sd3_1
X_21266_ _08527_ VGND VGND VPWR VPWR _08528_ sky130_fd_sc_hd__clkbuf_8
Xhold561 datamem.data_ram\[54\]\[6\] VGND VGND VPWR VPWR net1711 sky130_fd_sc_hd__dlygate4sd3_1
Xhold572 datamem.data_ram\[14\]\[6\] VGND VGND VPWR VPWR net1722 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold583 datamem.data_ram\[27\]\[5\] VGND VGND VPWR VPWR net1733 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20217_ datamem.data_ram\[29\]\[3\] _06920_ _06937_ datamem.data_ram\[24\]\[3\] _07509_
+ VGND VGND VPWR VPWR _07510_ sky130_fd_sc_hd__a221o_1
Xhold594 datamem.data_ram\[25\]\[3\] VGND VGND VPWR VPWR net1744 sky130_fd_sc_hd__dlygate4sd3_1
X_21197_ _07277_ _07737_ _07691_ _06915_ VGND VGND VPWR VPWR _08480_ sky130_fd_sc_hd__o22ai_1
X_28862_ _12692_ net2794 _12932_ VGND VGND VPWR VPWR _12935_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27813_ _12349_ VGND VGND VPWR VPWR _03753_ sky130_fd_sc_hd__clkbuf_1
X_22974__682 clknet_1_0__leaf__10082_ VGND VGND VPWR VPWR net808 sky130_fd_sc_hd__inv_2
X_20148_ datamem.data_ram\[62\]\[27\] _06627_ _06600_ _07440_ VGND VGND VPWR VPWR
+ _07441_ sky130_fd_sc_hd__o211a_1
XFILLER_0_218_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_202_5333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28793_ _12898_ VGND VGND VPWR VPWR _04184_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_202_5344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_202_5355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27744_ _12311_ VGND VGND VPWR VPWR _03722_ sky130_fd_sc_hd__clkbuf_1
X_20079_ datamem.data_ram\[38\]\[10\] _06717_ _06812_ datamem.data_ram\[35\]\[10\]
+ VGND VGND VPWR VPWR _07373_ sky130_fd_sc_hd__o22a_1
X_24956_ _10697_ VGND VGND VPWR VPWR _02548_ sky130_fd_sc_hd__clkbuf_1
Xhold1250 rvcpu.dp.plfd.PCPlus4D\[4\] VGND VGND VPWR VPWR net2400 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1261 rvcpu.dp.rf.reg_file_arr\[6\]\[15\] VGND VGND VPWR VPWR net2411 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_197_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23907_ clknet_1_0__leaf__10224_ VGND VGND VPWR VPWR _10225_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_194_5145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1272 rvcpu.dp.rf.reg_file_arr\[14\]\[18\] VGND VGND VPWR VPWR net2422 sky130_fd_sc_hd__dlygate4sd3_1
X_27675_ _12274_ VGND VGND VPWR VPWR _03690_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_213_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1283 datamem.data_ram\[10\]\[21\] VGND VGND VPWR VPWR net2433 sky130_fd_sc_hd__dlygate4sd3_1
X_24887_ _10660_ VGND VGND VPWR VPWR _02516_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_194_5156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_401 _06619_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1294 rvcpu.dp.rf.reg_file_arr\[20\]\[23\] VGND VGND VPWR VPWR net2444 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_412 _06667_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26626_ _10061_ _11659_ _11660_ net1338 VGND VGND VPWR VPWR _03255_ sky130_fd_sc_hd__a22o_1
X_29414_ clknet_leaf_11_clk _01149_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD2E\[25\] sky130_fd_sc_hd__dfxtp_1
X_14640_ net2299 _13213_ _13214_ VGND VGND VPWR VPWR _13215_ sky130_fd_sc_hd__mux2_1
XANTENNA_423 _06780_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23838_ _10215_ VGND VGND VPWR VPWR _01912_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_434 _06821_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_200_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_196_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_445 _07077_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_456 _08144_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_0__10226_ _10226_ VGND VGND VPWR VPWR clknet_0__10226_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_185_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_467 _08843_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_184_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29345_ clknet_leaf_204_clk _01080_ VGND VGND VPWR VPWR datamem.data_ram\[61\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_26557_ _11623_ VGND VGND VPWR VPWR _03223_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1__f__10126_ clknet_0__10126_ VGND VGND VPWR VPWR clknet_1_1__leaf__10126_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_67_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_478 _09317_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_52_clk clknet_5_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_52_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_196_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_489 _09728_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16310_ net2228 _14476_ _14511_ VGND VGND VPWR VPWR _14518_ sky130_fd_sc_hd__mux2_1
X_25508_ _09226_ _10921_ _10922_ VGND VGND VPWR VPWR _11010_ sky130_fd_sc_hd__and3_2
Xclkbuf_0__10157_ _10157_ VGND VGND VPWR VPWR clknet_0__10157_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_211_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17290_ _04907_ VGND VGND VPWR VPWR _01399_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29276_ _09225_ _09301_ _09230_ VGND VGND VPWR VPWR _13159_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_12_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_153_4163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_4174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16241_ _14479_ VGND VGND VPWR VPWR _01920_ sky130_fd_sc_hd__clkbuf_1
X_28227_ _12582_ VGND VGND VPWR VPWR _03934_ sky130_fd_sc_hd__clkbuf_1
X_25439_ _10762_ net2837 _10970_ VGND VGND VPWR VPWR _10976_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__10088_ _10088_ VGND VGND VPWR VPWR clknet_0__10088_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_125_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23732__324 clknet_1_1__leaf__10198_ VGND VGND VPWR VPWR net450 sky130_fd_sc_hd__inv_2
X_16172_ net2074 _14432_ _14422_ VGND VGND VPWR VPWR _14433_ sky130_fd_sc_hd__mux2_1
X_28158_ _12545_ VGND VGND VPWR VPWR _03902_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_209_5509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15123_ _13298_ _13349_ VGND VGND VPWR VPWR _13668_ sky130_fd_sc_hd__nand2_2
X_27109_ _11951_ VGND VGND VPWR VPWR _11952_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_23_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_149_Left_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28089_ _12445_ net2009 _12501_ VGND VGND VPWR VPWR _12509_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23847__411 clknet_1_1__leaf__10208_ VGND VGND VPWR VPWR net537 sky130_fd_sc_hd__inv_2
X_30120_ net482 _01855_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[10\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_15054_ _13598_ _13546_ _13600_ VGND VGND VPWR VPWR _13601_ sky130_fd_sc_hd__o21ai_1
X_19931_ _06797_ _07190_ _07202_ _07225_ VGND VGND VPWR VPWR _07226_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_220_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput2 net2 VGND VGND VPWR VPWR Instr[0] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_112_3181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30051_ net413 _01786_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[12\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_19862_ datamem.data_ram\[6\]\[1\] _07127_ _06977_ datamem.data_ram\[4\]\[1\] VGND
+ VGND VPWR VPWR _07157_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_183_4882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_4893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18813_ _05990_ _06026_ _06159_ _06109_ VGND VGND VPWR VPWR _06160_ sky130_fd_sc_hd__o22a_1
XFILLER_0_37_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19793_ datamem.data_ram\[53\]\[9\] _06703_ _07031_ _07087_ VGND VGND VPWR VPWR _07088_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_208_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_207_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18744_ _06093_ _06094_ _05706_ VGND VGND VPWR VPWR _06095_ sky130_fd_sc_hd__mux2_1
X_15956_ net3710 _13190_ _14311_ VGND VGND VPWR VPWR _14315_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_121_3406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_158_Left_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14907_ _13445_ _13457_ _13406_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__o21a_1
XFILLER_0_222_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18675_ _05693_ _05719_ VGND VGND VPWR VPWR _06030_ sky130_fd_sc_hd__nand2_1
X_30953_ clknet_leaf_255_clk _02688_ VGND VGND VPWR VPWR datamem.data_ram\[3\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_86_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15887_ _14278_ VGND VGND VPWR VPWR _02081_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_86_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17626_ _05085_ VGND VGND VPWR VPWR _01225_ sky130_fd_sc_hd__clkbuf_1
X_14838_ _13389_ _13390_ VGND VGND VPWR VPWR _13391_ sky130_fd_sc_hd__nand2_4
X_26487__41 clknet_1_1__leaf__10267_ VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__inv_2
X_30884_ clknet_leaf_3_clk _02619_ VGND VGND VPWR VPWR datamem.data_ram\[42\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_82_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_188_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23893__453 clknet_1_0__leaf__10222_ VGND VGND VPWR VPWR net579 sky130_fd_sc_hd__inv_2
XFILLER_0_187_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_82_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32623_ clknet_leaf_274_clk _04045_ VGND VGND VPWR VPWR datamem.data_ram\[20\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_14769_ _13286_ _13280_ VGND VGND VPWR VPWR _13322_ sky130_fd_sc_hd__nor2b_4
XFILLER_0_169_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17557_ _13187_ net3857 _05046_ VGND VGND VPWR VPWR _05049_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_43_clk clknet_5_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_43_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16508_ net2374 _14468_ _04489_ VGND VGND VPWR VPWR _04492_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17488_ _05012_ VGND VGND VPWR VPWR _01298_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_15_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32554_ clknet_leaf_239_clk _03976_ VGND VGND VPWR VPWR datamem.data_ram\[22\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_190_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19227_ rvcpu.dp.plde.ImmExtE\[26\] rvcpu.dp.plde.PCE\[26\] VGND VGND VPWR VPWR _06533_
+ sky130_fd_sc_hd__nor2_1
X_31505_ clknet_leaf_26_clk rvcpu.dp.lAuiPCE\[31\] VGND VGND VPWR VPWR rvcpu.dp.plem.lAuiPCM\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_16439_ _04454_ VGND VGND VPWR VPWR _01821_ sky130_fd_sc_hd__clkbuf_1
X_32485_ clknet_leaf_231_clk _03907_ VGND VGND VPWR VPWR datamem.data_ram\[25\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_167_Left_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31436_ clknet_leaf_102_clk _03139_ VGND VGND VPWR VPWR datamem.data_ram\[14\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_19158_ rvcpu.dp.plde.ImmExtE\[18\] rvcpu.dp.plde.PCE\[18\] VGND VGND VPWR VPWR _06473_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_171_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18109_ rvcpu.dp.plem.ALUResultM\[20\] _05476_ _05177_ VGND VGND VPWR VPWR _05477_
+ sky130_fd_sc_hd__mux2_1
X_31367_ clknet_leaf_17_clk _03070_ VGND VGND VPWR VPWR rvcpu.dp.plde.ImmExtE\[16\]
+ sky130_fd_sc_hd__dfxtp_2
X_19089_ _06412_ VGND VGND VPWR VPWR rvcpu.dp.lAuiPCE\[9\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_169_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21120_ datamem.data_ram\[44\]\[23\] datamem.data_ram\[45\]\[23\] _07874_ VGND VGND
+ VPWR VPWR _08409_ sky130_fd_sc_hd__mux2_1
X_30318_ net664 _02053_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[4\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31298_ clknet_leaf_65_clk _03001_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCPlus4E\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_54_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1099 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21051_ datamem.data_ram\[32\]\[31\] datamem.data_ram\[33\]\[31\] _07911_ VGND VGND
+ VPWR VPWR _08340_ sky130_fd_sc_hd__mux2_1
X_30249_ net603 _01984_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[6\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20002_ datamem.data_ram\[24\]\[2\] _06936_ _07294_ _07295_ VGND VGND VPWR VPWR _07296_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_185_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24810_ _10618_ VGND VGND VPWR VPWR _02481_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25790_ net1676 _11181_ _11177_ _11184_ VGND VGND VPWR VPWR _02895_ sky130_fd_sc_hd__o211a_1
XFILLER_0_119_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24741_ _10579_ VGND VGND VPWR VPWR _02451_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_2_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21953_ _08626_ _09180_ _09182_ _09184_ _08808_ VGND VGND VPWR VPWR _09185_ sky130_fd_sc_hd__a221o_1
XFILLER_0_55_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_179_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20904_ _07840_ _08192_ _08193_ VGND VGND VPWR VPWR _08194_ sky130_fd_sc_hd__or3_1
XFILLER_0_55_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27460_ _10113_ _10898_ _11713_ VGND VGND VPWR VPWR _12159_ sky130_fd_sc_hd__a21oi_2
X_24672_ _07123_ VGND VGND VPWR VPWR _10542_ sky130_fd_sc_hd__buf_8
XFILLER_0_90_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21884_ _08835_ _09119_ VGND VGND VPWR VPWR _09120_ sky130_fd_sc_hd__or2_1
XFILLER_0_132_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26411_ _11548_ _11549_ _11550_ _11551_ VGND VGND VPWR VPWR _03149_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_221_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20835_ _08124_ _06797_ VGND VGND VPWR VPWR _08125_ sky130_fd_sc_hd__nand2_8
X_27391_ _10739_ net2333 net86 VGND VGND VPWR VPWR _12115_ sky130_fd_sc_hd__mux2_1
XFILLER_0_178_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23143__818 clknet_1_1__leaf__10107_ VGND VGND VPWR VPWR net944 sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_34_clk clknet_5_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_34_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_132_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29130_ _09247_ net3185 _13076_ VGND VGND VPWR VPWR _13081_ sky130_fd_sc_hd__mux2_1
X_26342_ _11501_ net1522 _11496_ _11506_ VGND VGND VPWR VPWR _03125_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_13_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20766_ datamem.data_ram\[48\]\[6\] _07138_ _07123_ datamem.data_ram\[52\]\[6\] VGND
+ VGND VPWR VPWR _08056_ sky130_fd_sc_hd__a22o_1
XFILLER_0_175_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31746__123 VGND VGND VPWR VPWR _31746__123/HI net123 sky130_fd_sc_hd__conb_1
XFILLER_0_147_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29061_ _13044_ VGND VGND VPWR VPWR _04306_ sky130_fd_sc_hd__clkbuf_1
X_22505_ _09457_ _09653_ _09655_ _09658_ _09660_ VGND VGND VPWR VPWR _09661_ sky130_fd_sc_hd__o32a_1
X_26273_ net1593 _11467_ VGND VGND VPWR VPWR _11469_ sky130_fd_sc_hd__and2_1
XFILLER_0_162_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20697_ datamem.data_ram\[2\]\[5\] _07000_ _06927_ datamem.data_ram\[7\]\[5\] VGND
+ VGND VPWR VPWR _07988_ sky130_fd_sc_hd__a22o_1
XFILLER_0_220_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28012_ _12363_ net4404 net97 VGND VGND VPWR VPWR _12468_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25224_ _10851_ VGND VGND VPWR VPWR _02662_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22436_ rvcpu.dp.rf.reg_file_arr\[24\]\[7\] rvcpu.dp.rf.reg_file_arr\[25\]\[7\] rvcpu.dp.rf.reg_file_arr\[26\]\[7\]
+ rvcpu.dp.rf.reg_file_arr\[27\]\[7\] _09393_ _09395_ VGND VGND VPWR VPWR _09595_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_165_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25155_ _10766_ net2393 _10802_ VGND VGND VPWR VPWR _10810_ sky130_fd_sc_hd__mux2_1
X_22367_ _09528_ _09529_ _09426_ VGND VGND VPWR VPWR _09530_ sky130_fd_sc_hd__a21o_1
X_21318_ rvcpu.dp.plfd.InstrD\[15\] VGND VGND VPWR VPWR _08580_ sky130_fd_sc_hd__inv_2
XFILLER_0_206_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29963_ net333 _01698_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[15\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_25086_ _10774_ VGND VGND VPWR VPWR _02601_ sky130_fd_sc_hd__clkbuf_1
X_22298_ _09462_ VGND VGND VPWR VPWR _09463_ sky130_fd_sc_hd__clkbuf_8
X_28914_ _12962_ VGND VGND VPWR VPWR _04241_ sky130_fd_sc_hd__clkbuf_1
Xhold380 datamem.data_ram\[29\]\[2\] VGND VGND VPWR VPWR net1530 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21249_ _08510_ VGND VGND VPWR VPWR _08511_ sky130_fd_sc_hd__buf_2
XFILLER_0_229_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold391 datamem.data_ram\[4\]\[3\] VGND VGND VPWR VPWR net1541 sky130_fd_sc_hd__dlygate4sd3_1
X_29894_ net272 _01629_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[17\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28845_ _12739_ net3508 net69 VGND VGND VPWR VPWR _12926_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_196_5207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15810_ _14235_ VGND VGND VPWR VPWR _14236_ sky130_fd_sc_hd__buf_4
X_16790_ _04641_ VGND VGND VPWR VPWR _01649_ sky130_fd_sc_hd__clkbuf_1
X_25988_ net4422 _11315_ _11312_ _11318_ VGND VGND VPWR VPWR _02959_ sky130_fd_sc_hd__o211a_1
X_28776_ _12889_ VGND VGND VPWR VPWR _04176_ sky130_fd_sc_hd__clkbuf_1
X_23230__879 clknet_1_1__leaf__10125_ VGND VGND VPWR VPWR net1005 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_221_5797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15741_ _14198_ VGND VGND VPWR VPWR _14199_ sky130_fd_sc_hd__clkbuf_4
X_24939_ _10688_ VGND VGND VPWR VPWR _02540_ sky130_fd_sc_hd__clkbuf_1
X_27727_ _12302_ VGND VGND VPWR VPWR _03714_ sky130_fd_sc_hd__clkbuf_1
Xhold1080 datamem.data_ram\[17\]\[14\] VGND VGND VPWR VPWR net2230 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_172_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1091 datamem.data_ram\[56\]\[30\] VGND VGND VPWR VPWR net2241 sky130_fd_sc_hd__dlygate4sd3_1
X_18460_ _05625_ _05621_ _05633_ _05626_ _05579_ _05662_ VGND VGND VPWR VPWR _05823_
+ sky130_fd_sc_hd__mux4_1
X_15672_ _14130_ VGND VGND VPWR VPWR _14152_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_213_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27658_ _12265_ VGND VGND VPWR VPWR _03682_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_220 _09822_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_231 _10142_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_242 _11086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_212_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_184_101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_4214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17411_ _14193_ net2464 _04937_ VGND VGND VPWR VPWR _04971_ sky130_fd_sc_hd__mux2_1
X_14623_ net2323 _13201_ _13181_ VGND VGND VPWR VPWR _13202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_212_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_4225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18391_ _05642_ _05662_ VGND VGND VPWR VPWR _05755_ sky130_fd_sc_hd__nand2_1
XANTENNA_253 _13198_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26609_ _11652_ VGND VGND VPWR VPWR _03246_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27589_ _12228_ VGND VGND VPWR VPWR _03650_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_264 _13217_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_25_clk clknet_5_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_25_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_275 _13244_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_185_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_286 _13275_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_200_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17342_ _04934_ VGND VGND VPWR VPWR _01374_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_297 _13638_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29328_ clknet_leaf_144_clk _01063_ VGND VGND VPWR VPWR datamem.data_ram\[62\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__10109_ clknet_0__10109_ VGND VGND VPWR VPWR clknet_1_1__leaf__10109_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_184_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23656__255 clknet_1_1__leaf__10191_ VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__inv_2
X_17273_ _04897_ VGND VGND VPWR VPWR _01406_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29259_ _07125_ _09269_ _09230_ VGND VGND VPWR VPWR _13150_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_55_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_181_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19012_ _05300_ _05539_ _05666_ VGND VGND VPWR VPWR _06346_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16224_ _13250_ VGND VGND VPWR VPWR _14468_ sky130_fd_sc_hd__buf_4
XFILLER_0_141_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32270_ clknet_leaf_215_clk _03692_ VGND VGND VPWR VPWR datamem.data_ram\[33\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_114_3221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload206 clknet_leaf_200_clk VGND VGND VPWR VPWR clkload206/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_114_3232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload217 clknet_leaf_168_clk VGND VGND VPWR VPWR clkload217/Y sky130_fd_sc_hd__clkinv_1
XTAP_TAPCELL_ROW_114_3243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31221_ clknet_leaf_40_clk _02924_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCD\[10\] sky130_fd_sc_hd__dfxtp_1
Xclkload228 clknet_leaf_92_clk VGND VGND VPWR VPWR clkload228/Y sky130_fd_sc_hd__inv_6
XFILLER_0_24_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload239 clknet_leaf_119_clk VGND VGND VPWR VPWR clkload239/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_141_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16155_ _13177_ _14273_ VGND VGND VPWR VPWR _14421_ sky130_fd_sc_hd__nor2_2
XFILLER_0_12_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_185_4933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15106_ _13648_ _13650_ _13429_ VGND VGND VPWR VPWR _13651_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_110_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_185_4944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31152_ clknet_leaf_67_clk rvcpu.ALUResultE\[11\] VGND VGND VPWR VPWR rvcpu.dp.plem.ALUResultM\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_16086_ _14090_ _14271_ VGND VGND VPWR VPWR _14384_ sky130_fd_sc_hd__nor2_2
XFILLER_0_45_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30103_ net465 _01838_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[11\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_24142__646 clknet_1_0__leaf__10262_ VGND VGND VPWR VPWR net772 sky130_fd_sc_hd__inv_2
XFILLER_0_224_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15037_ _13581_ _13582_ _13583_ _13533_ VGND VGND VPWR VPWR _13584_ sky130_fd_sc_hd__o22a_1
X_19914_ datamem.data_ram\[38\]\[17\] _06630_ _06621_ datamem.data_ram\[36\]\[17\]
+ VGND VGND VPWR VPWR _07209_ sky130_fd_sc_hd__o22a_1
XFILLER_0_20_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31083_ clknet_leaf_95_clk _02818_ VGND VGND VPWR VPWR datamem.data_ram\[20\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2709 datamem.data_ram\[51\]\[24\] VGND VGND VPWR VPWR net3859 sky130_fd_sc_hd__dlygate4sd3_1
X_30034_ net396 _01769_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[13\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_19845_ datamem.data_ram\[42\]\[1\] _07136_ _07137_ datamem.data_ram\[43\]\[1\] _07139_
+ VGND VGND VPWR VPWR _07140_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_88_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_3951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19776_ _06716_ VGND VGND VPWR VPWR _07071_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_144_3962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16988_ _04746_ VGND VGND VPWR VPWR _01548_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_147_Right_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_218_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18727_ _06006_ _06078_ _05706_ VGND VGND VPWR VPWR _06079_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_84_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15939_ _14305_ VGND VGND VPWR VPWR _02056_ sky130_fd_sc_hd__clkbuf_1
X_31985_ clknet_leaf_117_clk _03407_ VGND VGND VPWR VPWR datamem.data_ram\[37\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_140_3848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23901__460 clknet_1_0__leaf__10223_ VGND VGND VPWR VPWR net586 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_140_3859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire36 _07964_ VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_189_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18658_ _05238_ _06000_ _06003_ _06013_ VGND VGND VPWR VPWR _06014_ sky130_fd_sc_hd__a211o_1
X_30936_ clknet_leaf_258_clk _02671_ VGND VGND VPWR VPWR datamem.data_ram\[40\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire47 _12403_ VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_4
Xwire58 _10812_ VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_4
XFILLER_0_87_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17609_ _13266_ net3453 _05068_ VGND VGND VPWR VPWR _05076_ sky130_fd_sc_hd__mux2_1
XFILLER_0_175_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18589_ _05676_ _05800_ VGND VGND VPWR VPWR _05948_ sky130_fd_sc_hd__nor2_1
X_30867_ clknet_leaf_280_clk _02602_ VGND VGND VPWR VPWR datamem.data_ram\[43\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_16_clk clknet_5_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_16_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_4_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20620_ _06652_ VGND VGND VPWR VPWR _07911_ sky130_fd_sc_hd__buf_6
X_32606_ clknet_leaf_243_clk _04028_ VGND VGND VPWR VPWR datamem.data_ram\[20\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_43_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30798_ clknet_leaf_227_clk _02533_ VGND VGND VPWR VPWR datamem.data_ram\[45\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_43_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_175_Left_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20551_ _07822_ _07830_ _07834_ _07841_ VGND VGND VPWR VPWR _07842_ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32537_ clknet_leaf_79_clk _03959_ VGND VGND VPWR VPWR datamem.data_ram\[23\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_138_3799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32468_ clknet_leaf_80_clk _03890_ VGND VGND VPWR VPWR datamem.data_ram\[26\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_20482_ datamem.data_ram\[62\]\[20\] _06627_ _06815_ datamem.data_ram\[61\]\[20\]
+ VGND VGND VPWR VPWR _07774_ sky130_fd_sc_hd__o22a_1
XFILLER_0_172_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22221_ rvcpu.dp.plfd.InstrD\[24\] rvcpu.dp.plfd.InstrD\[23\] VGND VGND VPWR VPWR
+ _09387_ sky130_fd_sc_hd__or2_2
X_31419_ clknet_leaf_53_clk _03122_ VGND VGND VPWR VPWR datamem.data_ram\[15\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32399_ clknet_leaf_75_clk _03821_ VGND VGND VPWR VPWR datamem.data_ram\[29\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23446__96 clknet_1_1__leaf__10156_ VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__inv_2
X_22152_ _09282_ net3721 net62 VGND VGND VPWR VPWR _09346_ sky130_fd_sc_hd__mux2_1
XFILLER_0_203_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21103_ _06623_ _08388_ _08390_ _08391_ VGND VGND VPWR VPWR _08392_ sky130_fd_sc_hd__a211o_1
XFILLER_0_2_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26960_ _11837_ _11854_ VGND VGND VPWR VPWR _11862_ sky130_fd_sc_hd__and2_1
X_22083_ rvcpu.dp.plem.WriteDataM\[24\] _09296_ _09215_ VGND VGND VPWR VPWR _09297_
+ sky130_fd_sc_hd__mux2_8
XFILLER_0_1_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__10129_ clknet_0__10129_ VGND VGND VPWR VPWR clknet_1_0__leaf__10129_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_22_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_184_Left_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25911_ net2171 _11256_ _11273_ _11274_ VGND VGND VPWR VPWR _02926_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_7_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21034_ datamem.data_ram\[22\]\[31\] _06625_ _06684_ datamem.data_ram\[20\]\[31\]
+ VGND VGND VPWR VPWR _08323_ sky130_fd_sc_hd__o22a_1
X_26891_ _11689_ _11810_ VGND VGND VPWR VPWR _11818_ sky130_fd_sc_hd__and2_1
XFILLER_0_201_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_227_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25842_ _11225_ VGND VGND VPWR VPWR _02906_ sky130_fd_sc_hd__clkbuf_1
X_28630_ _12811_ VGND VGND VPWR VPWR _04108_ sky130_fd_sc_hd__clkbuf_1
X_23761__350 clknet_1_0__leaf__10201_ VGND VGND VPWR VPWR net476 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_114_Right_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_214_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25773_ rvcpu.dp.pcreg.q\[10\] _11168_ VGND VGND VPWR VPWR _11171_ sky130_fd_sc_hd__and2_1
X_28561_ _12774_ VGND VGND VPWR VPWR _04076_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_215_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24724_ _06997_ VGND VGND VPWR VPWR _10570_ sky130_fd_sc_hd__buf_8
X_27512_ _12187_ VGND VGND VPWR VPWR _03614_ sky130_fd_sc_hd__clkbuf_1
X_28492_ _10782_ _12723_ _12730_ VGND VGND VPWR VPWR _04051_ sky130_fd_sc_hd__o21a_1
X_21936_ _08510_ _09168_ VGND VGND VPWR VPWR _09169_ sky130_fd_sc_hd__nor2_1
X_27443_ _12147_ net3196 net84 VGND VGND VPWR VPWR _12148_ sky130_fd_sc_hd__mux2_1
XFILLER_0_194_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24655_ _10405_ _10532_ VGND VGND VPWR VPWR _10533_ sky130_fd_sc_hd__and2_1
XFILLER_0_167_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21867_ _08682_ _09101_ _09103_ _08558_ VGND VGND VPWR VPWR _09104_ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_193_Left_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20818_ _06715_ _08101_ _08107_ _06712_ VGND VGND VPWR VPWR _08108_ sky130_fd_sc_hd__o211a_1
X_27374_ _12105_ VGND VGND VPWR VPWR _03558_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24586_ _10390_ net2848 _10491_ VGND VGND VPWR VPWR _10494_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21798_ _09030_ _09034_ _09038_ _08624_ VGND VGND VPWR VPWR _01049_ sky130_fd_sc_hd__o31a_1
XFILLER_0_132_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26325_ _10325_ _10935_ _10052_ VGND VGND VPWR VPWR _11497_ sky130_fd_sc_hd__and3_2
XFILLER_0_154_329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_4100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29113_ _09281_ net3403 _13067_ VGND VGND VPWR VPWR _13072_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_189_5022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20749_ datamem.data_ram\[9\]\[6\] _07833_ VGND VGND VPWR VPWR _08039_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_189_5033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29044_ _13018_ net1766 _13030_ _13035_ VGND VGND VPWR VPWR _04298_ sky130_fd_sc_hd__a31o_1
X_26256_ net1863 _11432_ VGND VGND VPWR VPWR _11460_ sky130_fd_sc_hd__and2_1
X_25207_ _10842_ VGND VGND VPWR VPWR _02654_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22419_ _09516_ _09578_ VGND VGND VPWR VPWR _09579_ sky130_fd_sc_hd__or2_1
X_26187_ _11430_ VGND VGND VPWR VPWR _03046_ sky130_fd_sc_hd__clkbuf_1
X_23399_ _10150_ VGND VGND VPWR VPWR _01538_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_227_5940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25138_ _10480_ net1999 _10793_ VGND VGND VPWR VPWR _10801_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_227_5951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_148_4040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_4051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_308 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25069_ _10764_ net2308 _10752_ VGND VGND VPWR VPWR _10765_ sky130_fd_sc_hd__mux2_1
X_17960_ _05327_ _05330_ VGND VGND VPWR VPWR _05331_ sky130_fd_sc_hd__and2_1
X_29946_ net316 _01681_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[15\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_223_5837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_223_5848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_223_5859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16911_ _04705_ VGND VGND VPWR VPWR _01584_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_217_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17891_ _05252_ _05263_ VGND VGND VPWR VPWR _05264_ sky130_fd_sc_hd__and2_1
X_29877_ net255 _01612_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[17\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19630_ _06925_ VGND VGND VPWR VPWR _06926_ sky130_fd_sc_hd__buf_4
X_28828_ _12756_ net3111 _12914_ VGND VGND VPWR VPWR _12917_ sky130_fd_sc_hd__mux2_1
X_16842_ net2452 _14461_ _04659_ VGND VGND VPWR VPWR _04669_ sky130_fd_sc_hd__mux2_1
X_23011__715 clknet_1_1__leaf__10086_ VGND VGND VPWR VPWR net841 sky130_fd_sc_hd__inv_2
X_19561_ datamem.data_ram\[5\]\[24\] _06823_ _06855_ _06856_ VGND VGND VPWR VPWR _06857_
+ sky130_fd_sc_hd__o211a_1
X_16773_ _04632_ VGND VGND VPWR VPWR _01657_ sky130_fd_sc_hd__clkbuf_1
X_28759_ _12692_ net2751 _12877_ VGND VGND VPWR VPWR _12880_ sky130_fd_sc_hd__mux2_1
XFILLER_0_176_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_5_3__f_clk clknet_2_0_0_clk VGND VGND VPWR VPWR clknet_5_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_18512_ _05865_ _05867_ _05869_ _05873_ VGND VGND VPWR VPWR _05874_ sky130_fd_sc_hd__a211o_1
X_15724_ _13265_ VGND VGND VPWR VPWR _14187_ sky130_fd_sc_hd__clkbuf_8
X_19492_ datamem.data_ram\[30\]\[16\] _06629_ _06620_ datamem.data_ram\[28\]\[16\]
+ VGND VGND VPWR VPWR _06788_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_17_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31770_ clknet_leaf_228_clk _03224_ VGND VGND VPWR VPWR datamem.data_ram\[1\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_178_4770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_624 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18443_ _05720_ _05805_ VGND VGND VPWR VPWR _05806_ sky130_fd_sc_hd__nor2_1
X_30721_ clknet_leaf_178_clk _02456_ VGND VGND VPWR VPWR datamem.data_ram\[49\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_197_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15655_ _14140_ VGND VGND VPWR VPWR _02183_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_4667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14606_ _13188_ VGND VGND VPWR VPWR _03201_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_174_4678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18374_ _05651_ _05657_ _05738_ VGND VGND VPWR VPWR _05739_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_139_860 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30652_ clknet_leaf_190_clk _02387_ VGND VGND VPWR VPWR datamem.data_ram\[51\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_15586_ _14100_ VGND VGND VPWR VPWR _02212_ sky130_fd_sc_hd__clkbuf_1
X_17325_ net4268 _13247_ _04924_ VGND VGND VPWR VPWR _04926_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30583_ clknet_leaf_189_clk _02318_ VGND VGND VPWR VPWR datamem.data_ram\[53\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32322_ clknet_leaf_81_clk _03744_ VGND VGND VPWR VPWR datamem.data_ram\[31\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17256_ _14175_ net4088 _04887_ VGND VGND VPWR VPWR _04889_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_226_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23931__486 clknet_1_0__leaf__10227_ VGND VGND VPWR VPWR net612 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_77_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16207_ _14456_ VGND VGND VPWR VPWR _01931_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32253_ clknet_leaf_167_clk _03675_ VGND VGND VPWR VPWR datamem.data_ram\[34\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_17187_ _04852_ VGND VGND VPWR VPWR _01447_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_226_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_3685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_3696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_1086 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31204_ clknet_leaf_27_clk _02907_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCPlus4D\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_579 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16138_ net4376 _13257_ _14407_ VGND VGND VPWR VPWR _14412_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_216_Right_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32184_ clknet_leaf_168_clk _03606_ VGND VGND VPWR VPWR datamem.data_ram\[37\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_23630__247 clknet_1_0__leaf__10181_ VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__inv_2
XFILLER_0_84_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23172__844 clknet_1_0__leaf__10110_ VGND VGND VPWR VPWR net970 sky130_fd_sc_hd__inv_2
Xhold3207 datamem.data_ram\[63\]\[10\] VGND VGND VPWR VPWR net4357 sky130_fd_sc_hd__dlygate4sd3_1
X_31135_ clknet_leaf_211_clk _02870_ VGND VGND VPWR VPWR datamem.data_ram\[4\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_16069_ _14375_ VGND VGND VPWR VPWR _01988_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_227_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold3218 datamem.data_ram\[52\]\[3\] VGND VGND VPWR VPWR net4368 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_5_clk clknet_5_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3229 datamem.data_ram\[54\]\[22\] VGND VGND VPWR VPWR net4379 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2506 datamem.data_ram\[41\]\[12\] VGND VGND VPWR VPWR net3656 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_36_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31066_ clknet_leaf_283_clk _02801_ VGND VGND VPWR VPWR datamem.data_ram\[8\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2517 datamem.data_ram\[29\]\[11\] VGND VGND VPWR VPWR net3667 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2528 rvcpu.dp.rf.reg_file_arr\[7\]\[4\] VGND VGND VPWR VPWR net3678 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2539 datamem.data_ram\[23\]\[11\] VGND VGND VPWR VPWR net3689 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_75_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_224_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30017_ net379 _01752_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[13\]\[4\] sky130_fd_sc_hd__dfxtp_1
Xhold1805 datamem.data_ram\[47\]\[24\] VGND VGND VPWR VPWR net2955 sky130_fd_sc_hd__dlygate4sd3_1
X_19828_ _06976_ VGND VGND VPWR VPWR _07123_ sky130_fd_sc_hd__buf_4
Xhold1816 datamem.data_ram\[1\]\[27\] VGND VGND VPWR VPWR net2966 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_209_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1827 datamem.data_ram\[19\]\[17\] VGND VGND VPWR VPWR net2977 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1838 datamem.data_ram\[16\]\[27\] VGND VGND VPWR VPWR net2988 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1849 datamem.data_ram\[21\]\[18\] VGND VGND VPWR VPWR net2999 sky130_fd_sc_hd__dlygate4sd3_1
X_19759_ datamem.data_ram\[50\]\[25\] _06803_ _06696_ datamem.data_ram\[48\]\[25\]
+ VGND VGND VPWR VPWR _07054_ sky130_fd_sc_hd__o22a_1
XFILLER_0_155_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_189_760 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23973__509 clknet_1_1__leaf__10238_ VGND VGND VPWR VPWR net635 sky130_fd_sc_hd__inv_2
X_22770_ _09433_ _09911_ _09789_ VGND VGND VPWR VPWR _09912_ sky130_fd_sc_hd__a21o_1
X_31968_ clknet_leaf_130_clk _03390_ VGND VGND VPWR VPWR datamem.data_ram\[54\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_911 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21721_ rvcpu.dp.rf.reg_file_arr\[8\]\[17\] rvcpu.dp.rf.reg_file_arr\[10\]\[17\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[17\] rvcpu.dp.rf.reg_file_arr\[11\]\[17\] _08649_
+ _08537_ VGND VGND VPWR VPWR _08966_ sky130_fd_sc_hd__mux4_2
XFILLER_0_56_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30919_ clknet_leaf_201_clk _02654_ VGND VGND VPWR VPWR datamem.data_ram\[40\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_101_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_646 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31899_ _04441_ net118 VGND VGND VPWR VPWR datamem.rd_data_mem\[4\] sky130_fd_sc_hd__dlxtn_1
XFILLER_0_17_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24440_ _09299_ _08059_ _10052_ VGND VGND VPWR VPWR _10406_ sky130_fd_sc_hd__and3_1
XFILLER_0_177_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21652_ rvcpu.dp.rf.reg_file_arr\[24\]\[14\] rvcpu.dp.rf.reg_file_arr\[25\]\[14\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[14\] rvcpu.dp.rf.reg_file_arr\[27\]\[14\] _08524_
+ _08527_ VGND VGND VPWR VPWR _08900_ sky130_fd_sc_hd__mux4_1
XFILLER_0_136_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20603_ datamem.data_ram\[61\]\[13\] _06723_ _06731_ datamem.data_ram\[59\]\[13\]
+ VGND VGND VPWR VPWR _07894_ sky130_fd_sc_hd__o22a_1
XFILLER_0_117_521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24371_ _10363_ VGND VGND VPWR VPWR _02297_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_62_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23791__376 clknet_1_0__leaf__10205_ VGND VGND VPWR VPWR net502 sky130_fd_sc_hd__inv_2
XFILLER_0_75_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21583_ _08673_ VGND VGND VPWR VPWR _08835_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_191_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26110_ _11390_ VGND VGND VPWR VPWR _03008_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_191_468 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27090_ _10402_ _11075_ VGND VGND VPWR VPWR _11941_ sky130_fd_sc_hd__nor2_1
X_20534_ _07824_ VGND VGND VPWR VPWR _07825_ sky130_fd_sc_hd__buf_6
X_24010__543 clknet_1_1__leaf__10241_ VGND VGND VPWR VPWR net669 sky130_fd_sc_hd__inv_2
XFILLER_0_117_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26041_ _11121_ net1799 _11339_ _11347_ VGND VGND VPWR VPWR _02983_ sky130_fd_sc_hd__a31o_1
XFILLER_0_162_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20465_ datamem.data_ram\[19\]\[20\] _06635_ _07753_ _07756_ VGND VGND VPWR VPWR
+ _07757_ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22204_ _09279_ net3251 _09371_ VGND VGND VPWR VPWR _09375_ sky130_fd_sc_hd__mux2_1
X_23184_ clknet_1_1__leaf__10108_ VGND VGND VPWR VPWR _10112_ sky130_fd_sc_hd__buf_1
X_20396_ _06741_ _07685_ _07687_ VGND VGND VPWR VPWR _07688_ sky130_fd_sc_hd__and3_1
X_29800_ clknet_leaf_203_clk _01535_ VGND VGND VPWR VPWR datamem.data_ram\[59\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22135_ _09248_ net3907 _09332_ VGND VGND VPWR VPWR _09337_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27992_ _12455_ VGND VGND VPWR VPWR _03826_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29731_ net1077 _01466_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[22\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26943_ _07182_ _11109_ _11839_ VGND VGND VPWR VPWR _11852_ sky130_fd_sc_hd__or3_1
X_22066_ _09283_ VGND VGND VPWR VPWR _01072_ sky130_fd_sc_hd__clkbuf_1
X_23685__281 clknet_1_1__leaf__10194_ VGND VGND VPWR VPWR net407 sky130_fd_sc_hd__inv_2
X_24164__6 clknet_1_1__leaf__10264_ VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__inv_2
X_21017_ datamem.data_ram\[50\]\[31\] datamem.data_ram\[51\]\[31\] _06652_ VGND VGND
+ VPWR VPWR _08306_ sky130_fd_sc_hd__mux2_1
X_29662_ net1008 _01397_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[24\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_26874_ _11795_ net1551 _11797_ _11807_ VGND VGND VPWR VPWR _03356_ sky130_fd_sc_hd__a31o_1
XFILLER_0_57_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28613_ _12802_ VGND VGND VPWR VPWR _04100_ sky130_fd_sc_hd__clkbuf_1
X_25825_ _11206_ _11207_ _11211_ VGND VGND VPWR VPWR _11212_ sky130_fd_sc_hd__and3_1
XFILLER_0_57_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29593_ net947 _01328_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[26\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_23149__824 clknet_1_1__leaf__10107_ VGND VGND VPWR VPWR net950 sky130_fd_sc_hd__inv_2
X_25756_ net1594 _11144_ _11147_ _11158_ VGND VGND VPWR VPWR _02887_ sky130_fd_sc_hd__o211a_1
X_28544_ _12764_ net2695 _12752_ VGND VGND VPWR VPWR _12765_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24707_ _10268_ _10327_ _10501_ VGND VGND VPWR VPWR _10561_ sky130_fd_sc_hd__a21oi_2
X_21919_ rvcpu.dp.rf.reg_file_arr\[4\]\[28\] rvcpu.dp.rf.reg_file_arr\[5\]\[28\] rvcpu.dp.rf.reg_file_arr\[6\]\[28\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[28\] _08628_ _08856_ VGND VGND VPWR VPWR _09153_
+ sky130_fd_sc_hd__mux4_1
X_25687_ _11105_ net1749 _11111_ _11115_ VGND VGND VPWR VPWR _02861_ sky130_fd_sc_hd__a31o_1
XFILLER_0_195_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28475_ _12460_ net4020 _12713_ VGND VGND VPWR VPWR _12720_ sky130_fd_sc_hd__mux2_1
X_22899_ _09433_ _10033_ _09789_ VGND VGND VPWR VPWR _10034_ sky130_fd_sc_hd__a21o_1
XFILLER_0_38_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15440_ _13358_ _13450_ _13489_ _13758_ _13893_ VGND VGND VPWR VPWR _13971_ sky130_fd_sc_hd__a32o_1
XFILLER_0_167_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_214_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27426_ _09251_ VGND VGND VPWR VPWR _12136_ sky130_fd_sc_hd__buf_2
X_24638_ _10388_ net3019 _10521_ VGND VGND VPWR VPWR _10523_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_216_5674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_216_5685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_194_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15371_ _13528_ _13553_ _13514_ VGND VGND VPWR VPWR _13905_ sky130_fd_sc_hd__o21ai_1
X_24569_ _10444_ net3569 _10482_ VGND VGND VPWR VPWR _10485_ sky130_fd_sc_hd__mux2_1
X_27357_ _12096_ VGND VGND VPWR VPWR _03550_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17110_ _04811_ VGND VGND VPWR VPWR _01483_ sky130_fd_sc_hd__clkbuf_1
X_26308_ net1847 _11478_ VGND VGND VPWR VPWR _11487_ sky130_fd_sc_hd__and2_1
X_18090_ _05456_ _05457_ VGND VGND VPWR VPWR _05458_ sky130_fd_sc_hd__or2_1
X_27288_ _11970_ _12054_ VGND VGND VPWR VPWR _12057_ sky130_fd_sc_hd__and2_1
XFILLER_0_135_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17041_ net2472 _14455_ _04768_ VGND VGND VPWR VPWR _04775_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26239_ _11379_ _03045_ _11454_ VGND VGND VPWR VPWR _03072_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29027_ _13025_ VGND VGND VPWR VPWR _04291_ sky130_fd_sc_hd__clkbuf_1
X_23121__798 clknet_1_0__leaf__10105_ VGND VGND VPWR VPWR net924 sky130_fd_sc_hd__inv_2
XFILLER_0_80_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap109 net110 VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_61_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_72_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23768__356 clknet_1_1__leaf__10202_ VGND VGND VPWR VPWR net482 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_72_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23425__77 clknet_1_0__leaf__10154_ VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__inv_2
XFILLER_0_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_221_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18992_ _05561_ _05728_ _06108_ _05556_ _06326_ VGND VGND VPWR VPWR _06327_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_167_4493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17943_ _05313_ _05314_ VGND VGND VPWR VPWR _05315_ sky130_fd_sc_hd__nand2_1
X_29929_ net299 _01664_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[16\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_225_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_221_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32940_ clknet_leaf_154_clk _04362_ VGND VGND VPWR VPWR datamem.data_ram\[6\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_17874_ rvcpu.dp.plde.Rs1E\[0\] _05162_ _05245_ rvcpu.dp.plde.Rs1E\[3\] _05246_ VGND
+ VGND VPWR VPWR _05247_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_105_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19613_ _06596_ _06875_ _06908_ VGND VGND VPWR VPWR _06909_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_105_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16825_ _04660_ VGND VGND VPWR VPWR _01625_ sky130_fd_sc_hd__clkbuf_1
X_32871_ clknet_leaf_282_clk _04293_ VGND VGND VPWR VPWR datamem.data_ram\[11\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_31822_ clknet_leaf_104_clk _03276_ VGND VGND VPWR VPWR datamem.data_ram\[9\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_176_4718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19544_ datamem.data_ram\[29\]\[24\] _06815_ _06670_ datamem.data_ram\[31\]\[24\]
+ _06839_ VGND VGND VPWR VPWR _06840_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_176_4729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16756_ net3217 _14442_ _04623_ VGND VGND VPWR VPWR _04624_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15707_ _14175_ net3164 _14173_ VGND VGND VPWR VPWR _14176_ sky130_fd_sc_hd__mux2_1
X_31753_ clknet_leaf_58_clk _03207_ VGND VGND VPWR VPWR datamem.data_ram\[45\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_19475_ datamem.data_ram\[54\]\[16\] _06764_ _06767_ _06770_ VGND VGND VPWR VPWR
+ _06771_ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16687_ _04575_ VGND VGND VPWR VPWR _04587_ sky130_fd_sc_hd__buf_4
XFILLER_0_186_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18426_ _05789_ _05775_ VGND VGND VPWR VPWR _05790_ sky130_fd_sc_hd__nand2_1
X_30704_ clknet_leaf_219_clk _02439_ VGND VGND VPWR VPWR datamem.data_ram\[49\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15638_ rvcpu.dp.plmw.RdW\[1\] _13178_ VGND VGND VPWR VPWR _14128_ sky130_fd_sc_hd__nor2_4
XFILLER_0_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31684_ clknet_leaf_37_clk _03142_ VGND VGND VPWR VPWR rvcpu.dp.pcreg.q\[2\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_150_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_174_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_1047 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18357_ rvcpu.dp.plde.ALUControlE\[3\] rvcpu.dp.plde.ALUControlE\[2\] VGND VGND VPWR
+ VPWR _05722_ sky130_fd_sc_hd__or2b_1
X_30635_ clknet_leaf_194_clk _02370_ VGND VGND VPWR VPWR datamem.data_ram\[51\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_3725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15569_ _14089_ _14090_ VGND VGND VPWR VPWR _14091_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_135_3736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_3747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17308_ net4384 _13222_ _04913_ VGND VGND VPWR VPWR _04917_ sky130_fd_sc_hd__mux2_1
XFILLER_0_185_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30566_ clknet_leaf_142_clk _02301_ VGND VGND VPWR VPWR datamem.data_ram\[54\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_18288_ _05652_ _00003_ VGND VGND VPWR VPWR _05653_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_25_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32305_ clknet_leaf_240_clk _03727_ VGND VGND VPWR VPWR datamem.data_ram\[32\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_24148__652 clknet_1_0__leaf__10262_ VGND VGND VPWR VPWR net778 sky130_fd_sc_hd__inv_2
XFILLER_0_226_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17239_ _14158_ net4234 _04876_ VGND VGND VPWR VPWR _04880_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23554__178 clknet_1_0__leaf__10174_ VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__inv_2
X_30497_ clknet_leaf_145_clk _02232_ VGND VGND VPWR VPWR datamem.data_ram\[57\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_568 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold902 rvcpu.dp.rf.reg_file_arr\[4\]\[7\] VGND VGND VPWR VPWR net2052 sky130_fd_sc_hd__dlygate4sd3_1
Xhold913 datamem.data_ram\[36\]\[23\] VGND VGND VPWR VPWR net2063 sky130_fd_sc_hd__dlygate4sd3_1
X_20250_ datamem.data_ram\[32\]\[3\] _06937_ _06961_ datamem.data_ram\[35\]\[3\] _07542_
+ VGND VGND VPWR VPWR _07543_ sky130_fd_sc_hd__a221o_1
XFILLER_0_12_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32236_ clknet_leaf_257_clk _03658_ VGND VGND VPWR VPWR datamem.data_ram\[35\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold924 rvcpu.dp.rf.reg_file_arr\[8\]\[26\] VGND VGND VPWR VPWR net2074 sky130_fd_sc_hd__dlygate4sd3_1
X_23096__775 clknet_1_0__leaf__10103_ VGND VGND VPWR VPWR net901 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_38_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold935 rvcpu.dp.rf.reg_file_arr\[12\]\[29\] VGND VGND VPWR VPWR net2085 sky130_fd_sc_hd__dlygate4sd3_1
Xhold946 rvcpu.dp.rf.reg_file_arr\[13\]\[0\] VGND VGND VPWR VPWR net2096 sky130_fd_sc_hd__dlygate4sd3_1
Xhold957 datamem.data_ram\[44\]\[14\] VGND VGND VPWR VPWR net2107 sky130_fd_sc_hd__dlygate4sd3_1
X_20181_ datamem.data_ram\[14\]\[11\] _06763_ _06737_ datamem.data_ram\[11\]\[11\]
+ _06741_ VGND VGND VPWR VPWR _07474_ sky130_fd_sc_hd__o221a_1
Xhold968 rvcpu.dp.rf.reg_file_arr\[2\]\[26\] VGND VGND VPWR VPWR net2118 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3004 rvcpu.dp.rf.reg_file_arr\[21\]\[23\] VGND VGND VPWR VPWR net4154 sky130_fd_sc_hd__dlygate4sd3_1
X_32167_ clknet_leaf_180_clk _03589_ VGND VGND VPWR VPWR datamem.data_ram\[38\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3015 datamem.data_ram\[39\]\[17\] VGND VGND VPWR VPWR net4165 sky130_fd_sc_hd__dlygate4sd3_1
Xhold979 rvcpu.dp.rf.reg_file_arr\[10\]\[6\] VGND VGND VPWR VPWR net2129 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3026 rvcpu.dp.rf.reg_file_arr\[14\]\[0\] VGND VGND VPWR VPWR net4176 sky130_fd_sc_hd__dlygate4sd3_1
X_31118_ clknet_leaf_109_clk _02853_ VGND VGND VPWR VPWR datamem.data_ram\[35\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3037 rvcpu.dp.rf.reg_file_arr\[15\]\[2\] VGND VGND VPWR VPWR net4187 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold3048 datamem.data_ram\[44\]\[11\] VGND VGND VPWR VPWR net4198 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2303 rvcpu.dp.rf.reg_file_arr\[28\]\[4\] VGND VGND VPWR VPWR net3453 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32098_ clknet_leaf_114_clk _03520_ VGND VGND VPWR VPWR datamem.data_ram\[23\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3059 rvcpu.dp.rf.reg_file_arr\[23\]\[8\] VGND VGND VPWR VPWR net4209 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2314 datamem.data_ram\[26\]\[30\] VGND VGND VPWR VPWR net3464 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2325 datamem.data_ram\[62\]\[11\] VGND VGND VPWR VPWR net3475 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23940_ clknet_1_0__leaf__10224_ VGND VGND VPWR VPWR _10228_ sky130_fd_sc_hd__buf_1
Xhold2336 datamem.data_ram\[55\]\[31\] VGND VGND VPWR VPWR net3486 sky130_fd_sc_hd__dlygate4sd3_1
X_31049_ clknet_leaf_236_clk _02784_ VGND VGND VPWR VPWR datamem.data_ram\[9\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2347 datamem.data_ram\[21\]\[25\] VGND VGND VPWR VPWR net3497 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1602 datamem.data_ram\[21\]\[9\] VGND VGND VPWR VPWR net2752 sky130_fd_sc_hd__dlygate4sd3_1
X_24040__569 clknet_1_0__leaf__10245_ VGND VGND VPWR VPWR net695 sky130_fd_sc_hd__inv_2
Xhold1613 datamem.data_ram\[40\]\[14\] VGND VGND VPWR VPWR net2763 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2358 datamem.data_ram\[14\]\[10\] VGND VGND VPWR VPWR net3508 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1624 datamem.data_ram\[21\]\[8\] VGND VGND VPWR VPWR net2774 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2369 datamem.data_ram\[6\]\[27\] VGND VGND VPWR VPWR net3519 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_196_1288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1635 rvcpu.dp.rf.reg_file_arr\[11\]\[20\] VGND VGND VPWR VPWR net2785 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1646 datamem.data_ram\[13\]\[29\] VGND VGND VPWR VPWR net2796 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1657 rvcpu.dp.rf.reg_file_arr\[4\]\[1\] VGND VGND VPWR VPWR net2807 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1668 datamem.data_ram\[10\]\[20\] VGND VGND VPWR VPWR net2818 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1679 rvcpu.dp.rf.reg_file_arr\[15\]\[27\] VGND VGND VPWR VPWR net2829 sky130_fd_sc_hd__dlygate4sd3_1
X_25610_ _11069_ VGND VGND VPWR VPWR _02830_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22822_ rvcpu.dp.rf.reg_file_arr\[0\]\[27\] rvcpu.dp.rf.reg_file_arr\[1\]\[27\] rvcpu.dp.rf.reg_file_arr\[2\]\[27\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[27\] _09714_ _09383_ VGND VGND VPWR VPWR _09961_
+ sky130_fd_sc_hd__mux4_1
X_26590_ _11081_ _11640_ VGND VGND VPWR VPWR _11642_ sky130_fd_sc_hd__and2_1
XFILLER_0_168_218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25541_ _11028_ VGND VGND VPWR VPWR _02802_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_189_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22753_ _09622_ _09893_ _09895_ VGND VGND VPWR VPWR _09896_ sky130_fd_sc_hd__a21o_1
Xclkbuf_1_1__f__10090_ clknet_0__10090_ VGND VGND VPWR VPWR clknet_1_1__leaf__10090_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_149_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21704_ _08842_ _08949_ VGND VGND VPWR VPWR _08950_ sky130_fd_sc_hd__or2_1
X_28260_ _12462_ net3076 _12592_ VGND VGND VPWR VPWR _12600_ sky130_fd_sc_hd__mux2_1
X_25472_ _10991_ net1659 _10984_ _10992_ VGND VGND VPWR VPWR _02769_ sky130_fd_sc_hd__a31o_1
XFILLER_0_17_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22684_ _09705_ _09822_ _09826_ _09830_ VGND VGND VPWR VPWR _09831_ sky130_fd_sc_hd__and4_1
XFILLER_0_109_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27211_ _12005_ net1535 _12007_ _12015_ VGND VGND VPWR VPWR _03485_ sky130_fd_sc_hd__a31o_1
X_24423_ _10393_ VGND VGND VPWR VPWR _02319_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_212_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28191_ _12445_ net2524 _12555_ VGND VGND VPWR VPWR _12563_ sky130_fd_sc_hd__mux2_1
X_21635_ rvcpu.dp.rf.reg_file_arr\[20\]\[13\] rvcpu.dp.rf.reg_file_arr\[21\]\[13\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[13\] rvcpu.dp.rf.reg_file_arr\[23\]\[13\] _08799_
+ _08800_ VGND VGND VPWR VPWR _08884_ sky130_fd_sc_hd__mux4_2
XFILLER_0_192_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27142_ _11956_ net1684 _11964_ _11973_ VGND VGND VPWR VPWR _03458_ sky130_fd_sc_hd__a31o_1
XFILLER_0_192_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24354_ _10354_ VGND VGND VPWR VPWR _02289_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_211_5560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21566_ rvcpu.dp.rf.reg_file_arr\[8\]\[9\] rvcpu.dp.rf.reg_file_arr\[10\]\[9\] rvcpu.dp.rf.reg_file_arr\[9\]\[9\]
+ rvcpu.dp.rf.reg_file_arr\[11\]\[9\] _08693_ _08818_ VGND VGND VPWR VPWR _08819_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_63_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_211_5571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23040__741 clknet_1_0__leaf__10089_ VGND VGND VPWR VPWR net867 sky130_fd_sc_hd__inv_2
XFILLER_0_144_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27073_ _11919_ net1673 _11923_ _11929_ VGND VGND VPWR VPWR _03433_ sky130_fd_sc_hd__a31o_1
X_20517_ _06659_ VGND VGND VPWR VPWR _07808_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_133_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24285_ _10315_ VGND VGND VPWR VPWR _02259_ sky130_fd_sc_hd__clkbuf_1
X_21497_ rvcpu.dp.rf.reg_file_arr\[8\]\[6\] rvcpu.dp.rf.reg_file_arr\[10\]\[6\] rvcpu.dp.rf.reg_file_arr\[9\]\[6\]
+ rvcpu.dp.rf.reg_file_arr\[11\]\[6\] _08560_ _08561_ VGND VGND VPWR VPWR _08753_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_90_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26024_ net1909 _11329_ _11146_ _11337_ VGND VGND VPWR VPWR _02976_ sky130_fd_sc_hd__o211a_1
X_23236_ clknet_1_1__leaf__10108_ VGND VGND VPWR VPWR _10126_ sky130_fd_sc_hd__buf_1
X_20448_ datamem.data_ram\[2\]\[20\] _06691_ _06619_ datamem.data_ram\[4\]\[20\] VGND
+ VGND VPWR VPWR _07740_ sky130_fd_sc_hd__o22a_1
XFILLER_0_140_1221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20379_ datamem.data_ram\[62\]\[28\] _06625_ _06684_ datamem.data_ram\[60\]\[28\]
+ _07670_ VGND VGND VPWR VPWR _07671_ sky130_fd_sc_hd__o221a_1
XFILLER_0_219_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22118_ _09325_ VGND VGND VPWR VPWR _09326_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_101_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27975_ _12443_ net2337 _12431_ VGND VGND VPWR VPWR _12444_ sky130_fd_sc_hd__mux2_1
X_29714_ net1060 _01449_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[22\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_14940_ _13303_ _13393_ VGND VGND VPWR VPWR _13489_ sky130_fd_sc_hd__nand2_4
X_26926_ _11822_ _11842_ VGND VGND VPWR VPWR _11843_ sky130_fd_sc_hd__and2_1
XFILLER_0_140_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22049_ _09267_ net3759 _09270_ VGND VGND VPWR VPWR _09271_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_162_4390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2870 datamem.data_ram\[20\]\[14\] VGND VGND VPWR VPWR net4020 sky130_fd_sc_hd__dlygate4sd3_1
X_29645_ net991 _01380_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[24\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14871_ _13422_ VGND VGND VPWR VPWR _13423_ sky130_fd_sc_hd__clkbuf_4
X_26857_ _11725_ _11039_ VGND VGND VPWR VPWR _11798_ sky130_fd_sc_hd__nor2_2
Xhold2881 datamem.data_ram\[49\]\[24\] VGND VGND VPWR VPWR net4031 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2892 rvcpu.dp.rf.reg_file_arr\[14\]\[14\] VGND VGND VPWR VPWR net4042 sky130_fd_sc_hd__dlygate4sd3_1
X_16610_ _04546_ VGND VGND VPWR VPWR _01734_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_214_163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25808_ rvcpu.dp.pcreg.q\[17\] _11191_ rvcpu.dp.pcreg.q\[18\] VGND VGND VPWR VPWR
+ _11198_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_187_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29576_ net930 _01311_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[26\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_17590_ _13238_ net2718 _05057_ VGND VGND VPWR VPWR _05066_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_218_5725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26788_ _11753_ net1654 _11748_ _11756_ VGND VGND VPWR VPWR _03321_ sky130_fd_sc_hd__a31o_1
XFILLER_0_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_218_5736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28527_ _12753_ VGND VGND VPWR VPWR _04063_ sky130_fd_sc_hd__clkbuf_1
X_16541_ _04509_ VGND VGND VPWR VPWR _01774_ sky130_fd_sc_hd__clkbuf_1
X_25739_ _08620_ _08621_ VGND VGND VPWR VPWR _11145_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_1182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24017__549 clknet_1_1__leaf__10242_ VGND VGND VPWR VPWR net675 sky130_fd_sc_hd__inv_2
XFILLER_0_214_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_4604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19260_ _06560_ _06561_ VGND VGND VPWR VPWR _06562_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28458_ _12443_ net3478 _12704_ VGND VGND VPWR VPWR _12711_ sky130_fd_sc_hd__mux2_1
X_16472_ net3205 _14432_ _04467_ VGND VGND VPWR VPWR _04473_ sky130_fd_sc_hd__mux2_1
XFILLER_0_214_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_1079 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18211_ _05390_ _05392_ VGND VGND VPWR VPWR _05576_ sky130_fd_sc_hd__nand2_1
X_15423_ _13940_ _13764_ _13954_ _13327_ VGND VGND VPWR VPWR _13955_ sky130_fd_sc_hd__o211a_1
X_27409_ _12124_ VGND VGND VPWR VPWR _03574_ sky130_fd_sc_hd__clkbuf_1
X_19191_ rvcpu.dp.plde.ImmExtE\[22\] rvcpu.dp.plde.PCE\[22\] VGND VGND VPWR VPWR _06502_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_155_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28389_ _12433_ net4174 _12669_ VGND VGND VPWR VPWR _12671_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15354_ _13528_ _13359_ _13634_ _13463_ VGND VGND VPWR VPWR _13889_ sky130_fd_sc_hd__o31ai_1
X_18142_ rvcpu.dp.plem.ALUResultM\[16\] _05507_ _05177_ VGND VGND VPWR VPWR _05508_
+ sky130_fd_sc_hd__mux2_1
X_30420_ net758 _02155_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[31\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23473__121 clknet_1_1__leaf__10158_ VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__inv_2
XFILLER_0_110_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15285_ _13599_ VGND VGND VPWR VPWR _13823_ sky130_fd_sc_hd__clkbuf_4
X_18073_ rvcpu.dp.plde.RD1E\[9\] _05267_ _05271_ _13250_ _05428_ VGND VGND VPWR VPWR
+ _05441_ sky130_fd_sc_hd__a221o_2
X_30351_ net697 _02086_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[3\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_3611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_3622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_169_4544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_680 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold209 datamem.data_ram\[0\]\[5\] VGND VGND VPWR VPWR net1359 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_169_4555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17024_ net2444 _14438_ _04757_ VGND VGND VPWR VPWR _04766_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30282_ clknet_leaf_140_clk _02017_ VGND VGND VPWR VPWR datamem.data_ram\[58\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32021_ clknet_leaf_129_clk _03443_ VGND VGND VPWR VPWR datamem.data_ram\[51\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_91_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xload_slew112 _09268_ VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__buf_8
X_23017__721 clknet_1_1__leaf__10086_ VGND VGND VPWR VPWR net847 sky130_fd_sc_hd__inv_2
X_18975_ _06255_ _06310_ _05707_ VGND VGND VPWR VPWR _06311_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17926_ rvcpu.dp.plem.ALUResultM\[28\] _05252_ VGND VGND VPWR VPWR _05299_ sky130_fd_sc_hd__or2_1
XFILLER_0_147_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_3562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_128_3573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32923_ clknet_leaf_262_clk _04345_ VGND VGND VPWR VPWR datamem.data_ram\[0\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_68_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17857_ rvcpu.dp.plem.ALUResultM\[7\] _05232_ _05176_ VGND VGND VPWR VPWR _05233_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_50_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16808_ _04651_ VGND VGND VPWR VPWR _01633_ sky130_fd_sc_hd__clkbuf_1
X_32854_ clknet_leaf_237_clk _04276_ VGND VGND VPWR VPWR datamem.data_ram\[11\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_17788_ _05154_ _05161_ rvcpu.dp.plde.RD2E\[2\] VGND VGND VPWR VPWR _05184_ sky130_fd_sc_hd__a21o_1
X_31805_ clknet_leaf_83_clk _03259_ VGND VGND VPWR VPWR datamem.data_ram\[46\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_1136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19527_ _06722_ VGND VGND VPWR VPWR _06823_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_191_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16739_ net4314 _14426_ _04612_ VGND VGND VPWR VPWR _04615_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32785_ clknet_leaf_254_clk _04207_ VGND VGND VPWR VPWR datamem.data_ram\[14\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19458_ _06728_ VGND VGND VPWR VPWR _06754_ sky130_fd_sc_hd__buf_8
X_31736_ net185 _03194_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[9\]\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_27_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23937__492 clknet_1_0__leaf__10227_ VGND VGND VPWR VPWR net618 sky130_fd_sc_hd__inv_2
X_18409_ _05388_ _05666_ _05772_ _05671_ VGND VGND VPWR VPWR _05773_ sky130_fd_sc_hd__a211o_1
X_31667_ clknet_leaf_70_clk net1264 VGND VGND VPWR VPWR rvcpu.dp.plmw.ALUResultW\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19389_ _06684_ VGND VGND VPWR VPWR _06685_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_98_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21420_ rvcpu.dp.rf.reg_file_arr\[20\]\[3\] rvcpu.dp.rf.reg_file_arr\[21\]\[3\] rvcpu.dp.rf.reg_file_arr\[22\]\[3\]
+ rvcpu.dp.rf.reg_file_arr\[23\]\[3\] _08524_ _08527_ VGND VGND VPWR VPWR _08679_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_98_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30618_ clknet_leaf_136_clk _02353_ VGND VGND VPWR VPWR datamem.data_ram\[52\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_228_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31598_ clknet_leaf_48_clk net1161 VGND VGND VPWR VPWR rvcpu.dp.plmw.PCPlus4W\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21351_ rvcpu.dp.plde.funct3E\[2\] rvcpu.dp.plde.funct3E\[0\] rvcpu.dp.plde.funct3E\[1\]
+ VGND VGND VPWR VPWR _08613_ sky130_fd_sc_hd__or3_1
XFILLER_0_154_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30549_ clknet_leaf_181_clk _02284_ VGND VGND VPWR VPWR datamem.data_ram\[55\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_20302_ _06716_ _07589_ _07594_ VGND VGND VPWR VPWR _07595_ sky130_fd_sc_hd__or3_1
Xhold710 rvcpu.dp.pcreg.q\[28\] VGND VGND VPWR VPWR net1860 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21282_ _08542_ _08543_ _08513_ VGND VGND VPWR VPWR _08544_ sky130_fd_sc_hd__o21ai_1
Xhold721 rvcpu.dp.plfd.PCD\[26\] VGND VGND VPWR VPWR net1871 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_229_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_188_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold732 rvcpu.dp.rf.reg_file_arr\[9\]\[15\] VGND VGND VPWR VPWR net1882 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23021_ clknet_1_0__leaf__10079_ VGND VGND VPWR VPWR _10087_ sky130_fd_sc_hd__buf_1
X_20233_ datamem.data_ram\[6\]\[3\] _06952_ _07524_ _07525_ VGND VGND VPWR VPWR _07526_
+ sky130_fd_sc_hd__a211o_1
Xhold743 rvcpu.dp.rf.reg_file_arr\[11\]\[18\] VGND VGND VPWR VPWR net1893 sky130_fd_sc_hd__dlygate4sd3_1
X_32219_ clknet_leaf_210_clk _03641_ VGND VGND VPWR VPWR datamem.data_ram\[35\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold754 rvcpu.dp.pcreg.q\[15\] VGND VGND VPWR VPWR net1904 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold765 rvcpu.dp.rf.reg_file_arr\[4\]\[9\] VGND VGND VPWR VPWR net1915 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold776 rvcpu.dp.rf.reg_file_arr\[1\]\[11\] VGND VGND VPWR VPWR net1926 sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 datamem.data_ram\[29\]\[23\] VGND VGND VPWR VPWR net1937 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_228_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20164_ datamem.data_ram\[22\]\[27\] _06718_ _07455_ _07456_ VGND VGND VPWR VPWR
+ _07457_ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold798 datamem.data_ram\[39\]\[31\] VGND VGND VPWR VPWR net1948 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2100 rvcpu.dp.rf.reg_file_arr\[26\]\[15\] VGND VGND VPWR VPWR net3250 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2111 datamem.data_ram\[27\]\[20\] VGND VGND VPWR VPWR net3261 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2122 datamem.data_ram\[53\]\[27\] VGND VGND VPWR VPWR net3272 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2133 datamem.data_ram\[43\]\[28\] VGND VGND VPWR VPWR net3283 sky130_fd_sc_hd__dlygate4sd3_1
X_27760_ _12149_ net3547 net48 VGND VGND VPWR VPWR _12320_ sky130_fd_sc_hd__mux2_1
Xhold2144 datamem.data_ram\[20\]\[21\] VGND VGND VPWR VPWR net3294 sky130_fd_sc_hd__dlygate4sd3_1
X_20095_ _06751_ _07383_ _07388_ VGND VGND VPWR VPWR _07389_ sky130_fd_sc_hd__or3_1
X_24972_ _10542_ _10601_ _10705_ VGND VGND VPWR VPWR _10706_ sky130_fd_sc_hd__a21oi_1
Xhold1410 datamem.data_ram\[45\]\[30\] VGND VGND VPWR VPWR net2560 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2155 datamem.data_ram\[1\]\[19\] VGND VGND VPWR VPWR net3305 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2166 datamem.data_ram\[37\]\[20\] VGND VGND VPWR VPWR net3316 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1421 rvcpu.dp.rf.reg_file_arr\[17\]\[6\] VGND VGND VPWR VPWR net2571 sky130_fd_sc_hd__dlygate4sd3_1
X_26711_ _11710_ VGND VGND VPWR VPWR _03290_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_207_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2177 datamem.data_ram\[8\]\[23\] VGND VGND VPWR VPWR net3327 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1432 rvcpu.dp.rf.reg_file_arr\[0\]\[31\] VGND VGND VPWR VPWR net2582 sky130_fd_sc_hd__dlygate4sd3_1
X_27691_ _12283_ VGND VGND VPWR VPWR _03697_ sky130_fd_sc_hd__clkbuf_1
Xhold2188 datamem.data_ram\[23\]\[27\] VGND VGND VPWR VPWR net3338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1443 datamem.data_ram\[36\]\[12\] VGND VGND VPWR VPWR net2593 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1454 datamem.data_ram\[41\]\[22\] VGND VGND VPWR VPWR net2604 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2199 datamem.data_ram\[20\]\[28\] VGND VGND VPWR VPWR net3349 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1465 datamem.data_ram\[11\]\[10\] VGND VGND VPWR VPWR net2615 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_197_814 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_220_clk clknet_5_21__leaf_clk VGND VGND VPWR VPWR clknet_leaf_220_clk
+ sky130_fd_sc_hd__clkbuf_8
X_29430_ net792 _01165_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[30\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_26642_ _11086_ _11663_ VGND VGND VPWR VPWR _11668_ sky130_fd_sc_hd__and2_1
Xhold1476 rvcpu.dp.rf.reg_file_arr\[22\]\[29\] VGND VGND VPWR VPWR net2626 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1487 datamem.data_ram\[33\]\[22\] VGND VGND VPWR VPWR net2637 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_200_5294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1498 rvcpu.dp.rf.reg_file_arr\[27\]\[12\] VGND VGND VPWR VPWR net2648 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0__10242_ _10242_ VGND VGND VPWR VPWR clknet_0__10242_ sky130_fd_sc_hd__clkbuf_16
X_22805_ rvcpu.dp.rf.reg_file_arr\[4\]\[26\] rvcpu.dp.rf.reg_file_arr\[5\]\[26\] rvcpu.dp.rf.reg_file_arr\[6\]\[26\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[26\] _09386_ _09419_ VGND VGND VPWR VPWR _09945_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29361_ clknet_leaf_267_clk _01096_ VGND VGND VPWR VPWR datamem.data_ram\[61\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_26573_ _10729_ net3165 _11629_ VGND VGND VPWR VPWR _11632_ sky130_fd_sc_hd__mux2_1
XFILLER_0_200_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_196_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20997_ datamem.data_ram\[25\]\[15\] _06653_ _08285_ _06922_ VGND VGND VPWR VPWR
+ _08286_ sky130_fd_sc_hd__o22a_1
X_23797__382 clknet_1_1__leaf__10205_ VGND VGND VPWR VPWR net508 sky130_fd_sc_hd__inv_2
XFILLER_0_223_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28312_ _12629_ VGND VGND VPWR VPWR _03972_ sky130_fd_sc_hd__clkbuf_1
X_25524_ _10076_ _11010_ VGND VGND VPWR VPWR _11019_ sky130_fd_sc_hd__and2_1
XFILLER_0_165_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0__10173_ _10173_ VGND VGND VPWR VPWR clknet_0__10173_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_67_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22736_ rvcpu.dp.rf.reg_file_arr\[4\]\[22\] rvcpu.dp.rf.reg_file_arr\[5\]\[22\] rvcpu.dp.rf.reg_file_arr\[6\]\[22\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[22\] _09464_ _09467_ VGND VGND VPWR VPWR _09880_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_213_5600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_192_5095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29292_ _13167_ VGND VGND VPWR VPWR _04414_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_213_5611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25455_ _10073_ _10981_ _10982_ net1375 VGND VGND VPWR VPWR _02762_ sky130_fd_sc_hd__a22o_1
X_28243_ _12445_ net2724 _12583_ VGND VGND VPWR VPWR _12591_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_755 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22667_ _09814_ VGND VGND VPWR VPWR _01142_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24406_ _10382_ VGND VGND VPWR VPWR _02313_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21618_ rvcpu.dp.rf.reg_file_arr\[24\]\[12\] rvcpu.dp.rf.reg_file_arr\[25\]\[12\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[12\] rvcpu.dp.rf.reg_file_arr\[27\]\[12\] _08549_
+ _08553_ VGND VGND VPWR VPWR _08868_ sky130_fd_sc_hd__mux4_1
X_25386_ _10076_ _10936_ VGND VGND VPWR VPWR _10945_ sky130_fd_sc_hd__and2_1
XFILLER_0_153_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28174_ _12371_ net3616 _12546_ VGND VGND VPWR VPWR _12554_ sky130_fd_sc_hd__mux2_1
X_22598_ _09399_ _09748_ _09472_ VGND VGND VPWR VPWR _09749_ sky130_fd_sc_hd__o21a_1
XFILLER_0_129_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_287_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_287_clk
+ sky130_fd_sc_hd__clkbuf_8
X_27125_ _11956_ net1647 _11952_ _11961_ VGND VGND VPWR VPWR _03453_ sky130_fd_sc_hd__a31o_1
X_24337_ _09256_ net4327 _10338_ VGND VGND VPWR VPWR _10345_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21549_ _08798_ _08801_ VGND VGND VPWR VPWR _08802_ sky130_fd_sc_hd__or2_1
X_15070_ _13615_ _13447_ VGND VGND VPWR VPWR _13616_ sky130_fd_sc_hd__nor2_1
X_27056_ _11918_ VGND VGND VPWR VPWR _11919_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_181_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24268_ _10306_ VGND VGND VPWR VPWR _02251_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26007_ _09457_ _11315_ _11325_ _11328_ VGND VGND VPWR VPWR _02968_ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24199_ _09230_ VGND VGND VPWR VPWR _10269_ sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_207_5459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_4430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_164_4441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_160_4327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18760_ _06109_ _05971_ _05962_ _05990_ VGND VGND VPWR VPWR _06110_ sky130_fd_sc_hd__o22a_1
XFILLER_0_101_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_160_4338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27958_ _12432_ VGND VGND VPWR VPWR _03815_ sky130_fd_sc_hd__clkbuf_1
X_15972_ _14323_ VGND VGND VPWR VPWR _02041_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_1046 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1272 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17711_ _05130_ VGND VGND VPWR VPWR _01185_ sky130_fd_sc_hd__clkbuf_1
X_14923_ _13303_ _13414_ VGND VGND VPWR VPWR _13472_ sky130_fd_sc_hd__nand2_4
X_26909_ _11813_ net1450 _11821_ _11830_ VGND VGND VPWR VPWR _03368_ sky130_fd_sc_hd__a31o_1
X_18691_ _05606_ _05429_ _05604_ _05596_ _05664_ _05669_ VGND VGND VPWR VPWR _06045_
+ sky130_fd_sc_hd__mux4_1
X_27889_ _12391_ net1436 _12393_ _12395_ VGND VGND VPWR VPWR _03783_ sky130_fd_sc_hd__a31o_1
Xhold70 rvcpu.dp.plem.lAuiPCM\[22\] VGND VGND VPWR VPWR net1220 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 rvcpu.dp.plem.PCPlus4M\[12\] VGND VGND VPWR VPWR net1231 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_211_clk clknet_5_22__leaf_clk VGND VGND VPWR VPWR clknet_leaf_211_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold92 rvcpu.dp.plem.lAuiPCM\[10\] VGND VGND VPWR VPWR net1242 sky130_fd_sc_hd__dlygate4sd3_1
X_29628_ net982 _01363_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[25\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_17642_ net3615 _13212_ _05093_ VGND VGND VPWR VPWR _05094_ sky130_fd_sc_hd__mux2_1
X_14854_ _13316_ _13325_ _13362_ _13406_ VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__o31a_1
XFILLER_0_187_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29559_ net913 _01294_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[27\]\[26\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_63_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17573_ _05045_ VGND VGND VPWR VPWR _05057_ sky130_fd_sc_hd__clkbuf_4
X_14785_ _13333_ _13337_ VGND VGND VPWR VPWR _13338_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19312_ _06605_ _06607_ VGND VGND VPWR VPWR _06608_ sky130_fd_sc_hd__nand2_8
XFILLER_0_187_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_4278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16524_ net3369 _14484_ _04466_ VGND VGND VPWR VPWR _04500_ sky130_fd_sc_hd__mux2_1
X_23047__747 clknet_1_0__leaf__10090_ VGND VGND VPWR VPWR net873 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_158_4289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32570_ clknet_leaf_285_clk _03992_ VGND VGND VPWR VPWR datamem.data_ram\[22\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_355 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31521_ clknet_leaf_48_clk net1240 VGND VGND VPWR VPWR rvcpu.dp.plem.PCPlus4M\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_19243_ _06535_ _06542_ _06543_ _06540_ VGND VGND VPWR VPWR _06547_ sky130_fd_sc_hd__a31o_1
XFILLER_0_42_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16455_ _04462_ VGND VGND VPWR VPWR _01813_ sky130_fd_sc_hd__clkbuf_1
X_15406_ _13429_ _13936_ _13937_ _13353_ VGND VGND VPWR VPWR _13938_ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19174_ rvcpu.dp.plde.ImmExtE\[20\] rvcpu.dp.plde.PCE\[20\] VGND VGND VPWR VPWR _06487_
+ sky130_fd_sc_hd__nand2_1
X_31452_ clknet_leaf_5_clk rvcpu.dp.SrcBFW_Mux.y\[10\] VGND VGND VPWR VPWR rvcpu.dp.plem.WriteDataM\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16386_ net2363 _14484_ _14524_ VGND VGND VPWR VPWR _14558_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_22_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18125_ rvcpu.dp.plem.ALUResultM\[18\] _05491_ _05176_ VGND VGND VPWR VPWR _05492_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30403_ net741 _02138_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[31\]\[14\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_278_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_278_clk
+ sky130_fd_sc_hd__clkbuf_8
X_15337_ _13692_ _13322_ _13872_ _13517_ _13458_ VGND VGND VPWR VPWR _13873_ sky130_fd_sc_hd__a221o_1
X_31383_ clknet_leaf_42_clk _03086_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCE\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_117_3296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18056_ rvcpu.dp.plde.ImmExtE\[8\] rvcpu.dp.SrcBFW_Mux.y\[8\] _05278_ VGND VGND VPWR
+ VPWR _05424_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1 _01038_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_30334_ net680 _02069_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[4\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_15268_ _13449_ _13658_ _13671_ VGND VGND VPWR VPWR _13807_ sky130_fd_sc_hd__or3_1
XFILLER_0_13_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_188_4997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17007_ _04756_ VGND VGND VPWR VPWR _04757_ sky130_fd_sc_hd__buf_4
X_15199_ _13430_ _13387_ _13320_ VGND VGND VPWR VPWR _13741_ sky130_fd_sc_hd__and3_1
X_30265_ net619 _02000_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[6\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_32004_ clknet_leaf_134_clk _03426_ VGND VGND VPWR VPWR datamem.data_ram\[52\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_30196_ net550 _01931_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[8\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18958_ _05549_ _06280_ _05638_ VGND VGND VPWR VPWR _06295_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_52_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17909_ _05275_ _05280_ VGND VGND VPWR VPWR _05282_ sky130_fd_sc_hd__nand2_1
XFILLER_0_206_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18889_ _06171_ _06230_ _05707_ VGND VGND VPWR VPWR _06231_ sky130_fd_sc_hd__mux2_1
XFILLER_0_193_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_202_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_202_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_222_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20920_ _08198_ _08203_ _08209_ _06916_ VGND VGND VPWR VPWR _08210_ sky130_fd_sc_hd__a211o_1
X_32906_ clknet_leaf_260_clk _04328_ VGND VGND VPWR VPWR datamem.data_ram\[7\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32837_ clknet_leaf_287_clk _04259_ VGND VGND VPWR VPWR datamem.data_ram\[12\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_20851_ datamem.data_ram\[2\]\[14\] datamem.data_ram\[3\]\[14\] _07835_ VGND VGND
+ VPWR VPWR _08141_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20782_ _07840_ _08070_ _08071_ rvcpu.dp.plem.ALUResultM\[3\] _07845_ VGND VGND VPWR
+ VPWR _08072_ sky130_fd_sc_hd__a221o_1
X_32768_ clknet_leaf_283_clk _04190_ VGND VGND VPWR VPWR datamem.data_ram\[15\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22521_ rvcpu.dp.rf.reg_file_arr\[28\]\[11\] rvcpu.dp.rf.reg_file_arr\[30\]\[11\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[11\] rvcpu.dp.rf.reg_file_arr\[31\]\[11\] _09558_
+ _09417_ VGND VGND VPWR VPWR _09676_ sky130_fd_sc_hd__mux4_1
XFILLER_0_174_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31719_ net168 _03177_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[9\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23870__432 clknet_1_0__leaf__10220_ VGND VGND VPWR VPWR net558 sky130_fd_sc_hd__inv_2
X_32699_ clknet_leaf_238_clk _04121_ VGND VGND VPWR VPWR datamem.data_ram\[17\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_25240_ _10729_ net3115 net55 VGND VGND VPWR VPWR _10860_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22452_ _09534_ _09610_ VGND VGND VPWR VPWR _09611_ sky130_fd_sc_hd__and2_1
XFILLER_0_174_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21403_ _08532_ VGND VGND VPWR VPWR _08663_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_269_clk clknet_5_19__leaf_clk VGND VGND VPWR VPWR clknet_leaf_269_clk
+ sky130_fd_sc_hd__clkbuf_8
X_25171_ _10820_ net4334 net58 VGND VGND VPWR VPWR _10821_ sky130_fd_sc_hd__mux2_1
XFILLER_0_199_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22383_ _09543_ _09544_ _09380_ VGND VGND VPWR VPWR _09545_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_59_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_1302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_59_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21334_ _08595_ rvcpu.dp.plde.RdE\[1\] VGND VGND VPWR VPWR _08596_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_199_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_791 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28930_ _12756_ net2770 _12968_ VGND VGND VPWR VPWR _12971_ sky130_fd_sc_hd__mux2_1
Xhold540 rvcpu.dp.pcreg.q\[10\] VGND VGND VPWR VPWR net1690 sky130_fd_sc_hd__dlygate4sd3_1
X_21265_ _08526_ VGND VGND VPWR VPWR _08527_ sky130_fd_sc_hd__clkbuf_8
Xhold551 datamem.data_ram\[8\]\[1\] VGND VGND VPWR VPWR net1701 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold562 datamem.data_ram\[25\]\[4\] VGND VGND VPWR VPWR net1712 sky130_fd_sc_hd__dlygate4sd3_1
X_20216_ datamem.data_ram\[27\]\[3\] _06941_ _06925_ datamem.data_ram\[31\]\[3\] VGND
+ VGND VPWR VPWR _07509_ sky130_fd_sc_hd__a22o_1
Xhold573 datamem.data_ram\[37\]\[1\] VGND VGND VPWR VPWR net1723 sky130_fd_sc_hd__dlygate4sd3_1
Xhold584 datamem.data_ram\[26\]\[4\] VGND VGND VPWR VPWR net1734 sky130_fd_sc_hd__dlygate4sd3_1
X_28861_ _12934_ VGND VGND VPWR VPWR _04216_ sky130_fd_sc_hd__clkbuf_1
Xhold595 datamem.data_ram\[62\]\[2\] VGND VGND VPWR VPWR net1745 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1070 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21196_ _08479_ VGND VGND VPWR VPWR _04417_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27812_ _12147_ net3382 net78 VGND VGND VPWR VPWR _12349_ sky130_fd_sc_hd__mux2_1
X_20147_ datamem.data_ram\[56\]\[27\] _06820_ _06617_ datamem.data_ram\[60\]\[27\]
+ _07439_ VGND VGND VPWR VPWR _07440_ sky130_fd_sc_hd__o221a_1
X_28792_ _12737_ net3527 net70 VGND VGND VPWR VPWR _12898_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_202_5334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_202_5345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27743_ _12132_ net3538 _12307_ VGND VGND VPWR VPWR _12311_ sky130_fd_sc_hd__mux2_1
X_20078_ datamem.data_ram\[43\]\[10\] _06829_ _06806_ datamem.data_ram\[44\]\[10\]
+ _07371_ VGND VGND VPWR VPWR _07372_ sky130_fd_sc_hd__o221a_1
X_24955_ _10385_ net2710 _10696_ VGND VGND VPWR VPWR _10697_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1240 datamem.data_ram\[33\]\[13\] VGND VGND VPWR VPWR net2390 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1251 datamem.data_ram\[59\]\[27\] VGND VGND VPWR VPWR net2401 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1262 rvcpu.dp.rf.reg_file_arr\[17\]\[13\] VGND VGND VPWR VPWR net2412 sky130_fd_sc_hd__dlygate4sd3_1
X_23906_ clknet_1_1__leaf__10078_ VGND VGND VPWR VPWR _10224_ sky130_fd_sc_hd__buf_1
Xhold1273 datamem.data_ram\[32\]\[16\] VGND VGND VPWR VPWR net2423 sky130_fd_sc_hd__dlygate4sd3_1
X_27674_ _12087_ net3784 net51 VGND VGND VPWR VPWR _12274_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_194_5146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24886_ _10439_ net3211 _10659_ VGND VGND VPWR VPWR _10660_ sky130_fd_sc_hd__mux2_1
Xhold1284 rvcpu.dp.rf.reg_file_arr\[7\]\[11\] VGND VGND VPWR VPWR net2434 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_194_5157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_402 _06619_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29413_ clknet_leaf_290_clk _01148_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD2E\[24\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1295 rvcpu.dp.rf.reg_file_arr\[4\]\[17\] VGND VGND VPWR VPWR net2445 sky130_fd_sc_hd__dlygate4sd3_1
X_26625_ _10058_ _11659_ _11660_ net1325 VGND VGND VPWR VPWR _03254_ sky130_fd_sc_hd__a22o_1
XANTENNA_413 _06667_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_424 _06783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23837_ _09318_ net3002 _10210_ VGND VGND VPWR VPWR _10215_ sky130_fd_sc_hd__mux2_1
XFILLER_0_213_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_435 _06922_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_212_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_446 _07832_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_0__10225_ _10225_ VGND VGND VPWR VPWR clknet_0__10225_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_196_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_184_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_457 _08361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_1_1__f__10125_ clknet_0__10125_ VGND VGND VPWR VPWR clknet_1_1__leaf__10125_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_36_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29344_ clknet_leaf_204_clk _01079_ VGND VGND VPWR VPWR datamem.data_ram\[61\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_468 _08848_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26556_ _10816_ net2944 _11620_ VGND VGND VPWR VPWR _11623_ sky130_fd_sc_hd__mux2_1
XANTENNA_479 _09317_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_211_1041 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25507_ _11008_ VGND VGND VPWR VPWR _11009_ sky130_fd_sc_hd__buf_2
XFILLER_0_177_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0__10156_ _10156_ VGND VGND VPWR VPWR clknet_0__10156_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_165_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29275_ _13158_ VGND VGND VPWR VPWR _04406_ sky130_fd_sc_hd__clkbuf_1
X_22719_ rvcpu.dp.rf.reg_file_arr\[0\]\[21\] rvcpu.dp.rf.reg_file_arr\[1\]\[21\] rvcpu.dp.rf.reg_file_arr\[2\]\[21\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[21\] _09477_ _09466_ VGND VGND VPWR VPWR _09864_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_193_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_4164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16240_ net2071 _14478_ _14464_ VGND VGND VPWR VPWR _14479_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28226_ _12371_ net3329 _12574_ VGND VGND VPWR VPWR _12582_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_153_4175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25438_ _10975_ VGND VGND VPWR VPWR _02752_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__10087_ _10087_ VGND VGND VPWR VPWR clknet_0__10087_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_165_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25369_ _07131_ _07154_ VGND VGND VPWR VPWR _10935_ sky130_fd_sc_hd__nor2_2
XFILLER_0_152_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28157_ _12462_ net3983 _12537_ VGND VGND VPWR VPWR _12545_ sky130_fd_sc_hd__mux2_1
X_16171_ _13197_ VGND VGND VPWR VPWR _14432_ sky130_fd_sc_hd__buf_4
XFILLER_0_51_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_959 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15122_ _13425_ _13428_ _13494_ _13666_ VGND VGND VPWR VPWR _13667_ sky130_fd_sc_hd__and4_1
X_27108_ _11109_ _10778_ VGND VGND VPWR VPWR _11951_ sky130_fd_sc_hd__or2_1
XFILLER_0_105_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28088_ _12508_ VGND VGND VPWR VPWR _03869_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_1113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15053_ _13599_ _13473_ VGND VGND VPWR VPWR _13600_ sky130_fd_sc_hd__nor2_1
X_19930_ _07071_ _07208_ _07213_ _07224_ VGND VGND VPWR VPWR _07225_ sky130_fd_sc_hd__o31a_1
X_27039_ _11904_ net1726 _11897_ _11908_ VGND VGND VPWR VPWR _03420_ sky130_fd_sc_hd__a31o_1
Xoutput3 net3 VGND VGND VPWR VPWR Instr[10] sky130_fd_sc_hd__buf_2
XFILLER_0_142_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_128_Right_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_3182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_3193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30050_ net412 _01785_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[12\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_19861_ datamem.data_ram\[5\]\[1\] _07132_ _07125_ datamem.data_ram\[7\]\[1\] _07155_
+ VGND VGND VPWR VPWR _07156_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_183_4883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_4894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18812_ _06158_ VGND VGND VPWR VPWR _06159_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19792_ datamem.data_ram\[48\]\[9\] _06778_ _06766_ datamem.data_ram\[52\]\[9\] _07086_
+ VGND VGND VPWR VPWR _07087_ sky130_fd_sc_hd__o221a_1
XFILLER_0_207_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18743_ _05437_ _05610_ _05408_ _05606_ _05665_ _05670_ VGND VGND VPWR VPWR _06094_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15955_ _14314_ VGND VGND VPWR VPWR _02049_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_222_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14906_ _13413_ _13453_ _13456_ _13325_ VGND VGND VPWR VPWR _13457_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_121_3407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18674_ _05696_ _05862_ VGND VGND VPWR VPWR _06029_ sky130_fd_sc_hd__nand2_1
X_30952_ clknet_leaf_257_clk _02687_ VGND VGND VPWR VPWR datamem.data_ram\[3\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_86_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15886_ net3215 _13187_ _14275_ VGND VGND VPWR VPWR _14278_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_86_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17625_ net4223 _13186_ _05082_ VGND VGND VPWR VPWR _05085_ sky130_fd_sc_hd__mux2_1
X_14837_ _13288_ _13280_ VGND VGND VPWR VPWR _13390_ sky130_fd_sc_hd__nand2_4
XFILLER_0_203_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30883_ clknet_leaf_280_clk _02618_ VGND VGND VPWR VPWR datamem.data_ram\[42\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32622_ clknet_leaf_271_clk _04044_ VGND VGND VPWR VPWR datamem.data_ram\[20\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17556_ _05048_ VGND VGND VPWR VPWR _01258_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_82_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14768_ _13280_ _13286_ VGND VGND VPWR VPWR _13321_ sky130_fd_sc_hd__nor2b_4
XFILLER_0_187_187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16507_ _04491_ VGND VGND VPWR VPWR _01790_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32553_ clknet_leaf_244_clk _03975_ VGND VGND VPWR VPWR datamem.data_ram\[22\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17487_ _13184_ net4089 _05010_ VGND VGND VPWR VPWR _05012_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14699_ rvcpu.dp.plmw.ALUResultW\[6\] rvcpu.dp.plmw.ReadDataW\[6\] rvcpu.dp.plmw.PCPlus4W\[6\]
+ rvcpu.dp.plmw.lAuiPCW\[6\] _13192_ _13193_ VGND VGND VPWR VPWR _13259_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_119_3347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19226_ _06532_ VGND VGND VPWR VPWR rvcpu.dp.lAuiPCE\[26\] sky130_fd_sc_hd__clkbuf_1
X_31504_ clknet_leaf_24_clk rvcpu.dp.lAuiPCE\[30\] VGND VGND VPWR VPWR rvcpu.dp.plem.lAuiPCM\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_119_3358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16438_ net2457 _14468_ _04451_ VGND VGND VPWR VPWR _04454_ sky130_fd_sc_hd__mux2_1
X_32484_ clknet_leaf_232_clk _03906_ VGND VGND VPWR VPWR datamem.data_ram\[25\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_229_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31435_ clknet_leaf_53_clk _03138_ VGND VGND VPWR VPWR datamem.data_ram\[14\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_19157_ _06445_ _06459_ _06465_ _06449_ _06466_ VGND VGND VPWR VPWR _06472_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_171_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16369_ _14549_ VGND VGND VPWR VPWR _01854_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_41_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18108_ _13216_ rvcpu.dp.plde.RD2E\[20\] _05196_ VGND VGND VPWR VPWR _05476_ sky130_fd_sc_hd__mux2_1
X_19088_ _06411_ rvcpu.dp.plde.ImmExtE\[9\] _06355_ VGND VGND VPWR VPWR _06412_ sky130_fd_sc_hd__mux2_1
X_31366_ clknet_leaf_13_clk _03069_ VGND VGND VPWR VPWR rvcpu.dp.plde.ImmExtE\[15\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_14_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18039_ rvcpu.dp.plde.ImmExtE\[11\] rvcpu.dp.SrcBFW_Mux.y\[11\] _05277_ VGND VGND
+ VPWR VPWR _05409_ sky130_fd_sc_hd__mux2_2
X_30317_ net663 _02052_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[4\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_31297_ clknet_leaf_38_clk _03000_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCPlus4E\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_631 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22958__667 clknet_1_0__leaf__10081_ VGND VGND VPWR VPWR net793 sky130_fd_sc_hd__inv_2
X_21050_ datamem.data_ram\[38\]\[31\] datamem.data_ram\[39\]\[31\] _07826_ VGND VGND
+ VPWR VPWR _08339_ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30248_ net602 _01983_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[6\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20001_ datamem.data_ram\[26\]\[2\] _06930_ _06924_ datamem.data_ram\[31\]\[2\] _06677_
+ VGND VGND VPWR VPWR _07295_ sky130_fd_sc_hd__a221o_1
XFILLER_0_185_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30179_ clknet_leaf_194_clk _01914_ VGND VGND VPWR VPWR datamem.data_ram\[58\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_226_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24740_ _10454_ net2114 _10571_ VGND VGND VPWR VPWR _10579_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21952_ _08531_ _09183_ _08806_ VGND VGND VPWR VPWR _09184_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_2_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20903_ _07635_ datamem.data_ram\[14\]\[22\] datamem.data_ram\[15\]\[22\] _07832_
+ _07867_ VGND VGND VPWR VPWR _08193_ sky130_fd_sc_hd__o221a_1
X_24671_ _10538_ net1342 _10531_ _10541_ VGND VGND VPWR VPWR _02419_ sky130_fd_sc_hd__a31o_1
XFILLER_0_210_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21883_ rvcpu.dp.rf.reg_file_arr\[8\]\[26\] rvcpu.dp.rf.reg_file_arr\[10\]\[26\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[26\] rvcpu.dp.rf.reg_file_arr\[11\]\[26\] _08635_
+ _08637_ VGND VGND VPWR VPWR _09119_ sky130_fd_sc_hd__mux4_1
X_26410_ _13539_ _11152_ _10780_ VGND VGND VPWR VPWR _11551_ sky130_fd_sc_hd__a21o_1
XFILLER_0_167_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20834_ rvcpu.dp.plem.ALUResultM\[5\] VGND VGND VPWR VPWR _08124_ sky130_fd_sc_hd__clkbuf_8
X_27390_ _12114_ VGND VGND VPWR VPWR _03565_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_193_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26341_ _11064_ _11497_ VGND VGND VPWR VPWR _11506_ sky130_fd_sc_hd__and2_1
X_20765_ datamem.data_ram\[54\]\[6\] _07159_ _07137_ datamem.data_ram\[51\]\[6\] VGND
+ VGND VPWR VPWR _08055_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23716__309 clknet_1_1__leaf__10197_ VGND VGND VPWR VPWR net435 sky130_fd_sc_hd__inv_2
XFILLER_0_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_175_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22504_ _09469_ _09659_ _09457_ VGND VGND VPWR VPWR _09660_ sky130_fd_sc_hd__o21ai_1
X_26272_ _11468_ VGND VGND VPWR VPWR _03093_ sky130_fd_sc_hd__clkbuf_1
X_29060_ _09278_ net4280 net65 VGND VGND VPWR VPWR _13044_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20696_ _06916_ _07970_ _07975_ _07986_ VGND VGND VPWR VPWR _07987_ sky130_fd_sc_hd__a31o_1
XFILLER_0_52_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25223_ _10756_ net3444 _10848_ VGND VGND VPWR VPWR _10851_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28011_ _12467_ VGND VGND VPWR VPWR _03833_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_220_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22435_ _09594_ VGND VGND VPWR VPWR _01130_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_190_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25154_ _10809_ VGND VGND VPWR VPWR _02634_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22366_ rvcpu.dp.rf.reg_file_arr\[4\]\[3\] rvcpu.dp.rf.reg_file_arr\[5\]\[3\] rvcpu.dp.rf.reg_file_arr\[6\]\[3\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[3\] _09423_ _09424_ VGND VGND VPWR VPWR _09529_ sky130_fd_sc_hd__mux4_1
XFILLER_0_60_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21317_ rvcpu.dp.plfd.InstrD\[19\] rvcpu.dp.plfd.InstrD\[18\] VGND VGND VPWR VPWR
+ _08579_ sky130_fd_sc_hd__or2_2
XFILLER_0_130_441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29962_ net332 _01697_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[15\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_25085_ _10735_ net3245 net89 VGND VGND VPWR VPWR _10774_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22297_ _09392_ VGND VGND VPWR VPWR _09462_ sky130_fd_sc_hd__buf_4
X_28913_ _12692_ net3549 _12959_ VGND VGND VPWR VPWR _12962_ sky130_fd_sc_hd__mux2_1
Xhold370 datamem.data_ram\[49\]\[1\] VGND VGND VPWR VPWR net1520 sky130_fd_sc_hd__dlygate4sd3_1
X_21248_ _08509_ VGND VGND VPWR VPWR _08510_ sky130_fd_sc_hd__buf_2
Xhold381 datamem.data_ram\[50\]\[2\] VGND VGND VPWR VPWR net1531 sky130_fd_sc_hd__dlygate4sd3_1
X_29893_ net271 _01628_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[17\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_229_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold392 datamem.data_ram\[55\]\[6\] VGND VGND VPWR VPWR net1542 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_225_5890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28844_ _12925_ VGND VGND VPWR VPWR _04208_ sky130_fd_sc_hd__clkbuf_1
X_21179_ _06582_ VGND VGND VPWR VPWR _08468_ sky130_fd_sc_hd__buf_2
XFILLER_0_102_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_196_5208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28775_ _12754_ net3256 _12887_ VGND VGND VPWR VPWR _12889_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25987_ net7 _11317_ VGND VGND VPWR VPWR _11318_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_221_5798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_204_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27726_ _12087_ net3660 net49 VGND VGND VPWR VPWR _12302_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15740_ _14197_ _14129_ VGND VGND VPWR VPWR _14198_ sky130_fd_sc_hd__nand2_2
X_24938_ _10439_ net3517 _10687_ VGND VGND VPWR VPWR _10688_ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_942 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1070 rvcpu.dp.rf.reg_file_arr\[16\]\[4\] VGND VGND VPWR VPWR net2220 sky130_fd_sc_hd__dlygate4sd3_1
X_24192__32 clknet_1_1__leaf__10266_ VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__inv_2
XFILLER_0_213_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1081 rvcpu.dp.rf.reg_file_arr\[9\]\[20\] VGND VGND VPWR VPWR net2231 sky130_fd_sc_hd__dlygate4sd3_1
X_23877__438 clknet_1_0__leaf__10221_ VGND VGND VPWR VPWR net564 sky130_fd_sc_hd__inv_2
XFILLER_0_73_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_197_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1092 rvcpu.dp.rf.reg_file_arr\[19\]\[20\] VGND VGND VPWR VPWR net2242 sky130_fd_sc_hd__dlygate4sd3_1
X_27657_ _12149_ net3712 net79 VGND VGND VPWR VPWR _12265_ sky130_fd_sc_hd__mux2_1
X_15671_ _13212_ VGND VGND VPWR VPWR _14151_ sky130_fd_sc_hd__buf_4
X_24869_ _10465_ net3543 net92 VGND VGND VPWR VPWR _10651_ sky130_fd_sc_hd__mux2_1
XANTENNA_210 _09560_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_221 _09822_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_232 _10142_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_4204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17410_ _04970_ VGND VGND VPWR VPWR _01334_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_243 _11089_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14622_ _13200_ VGND VGND VPWR VPWR _13201_ sky130_fd_sc_hd__buf_4
X_26608_ _10814_ net2352 _11650_ VGND VGND VPWR VPWR _11652_ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_4215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18390_ _05751_ _05753_ _05676_ VGND VGND VPWR VPWR _05754_ sky130_fd_sc_hd__mux2_1
XANTENNA_254 _13198_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_184_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_4226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27588_ _12132_ net3592 _12224_ VGND VGND VPWR VPWR _12228_ sky130_fd_sc_hd__mux2_1
XANTENNA_265 _13217_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_0__10208_ _10208_ VGND VGND VPWR VPWR clknet_0__10208_ sky130_fd_sc_hd__clkbuf_16
XANTENNA_276 _13244_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29327_ clknet_leaf_144_clk _01062_ VGND VGND VPWR VPWR datamem.data_ram\[62\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_17341_ net4443 _13271_ _04924_ VGND VGND VPWR VPWR _04934_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__10108_ clknet_0__10108_ VGND VGND VPWR VPWR clknet_1_1__leaf__10108_
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_287 _13275_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26539_ _11517_ net1620 _11608_ _11613_ VGND VGND VPWR VPWR _03215_ sky130_fd_sc_hd__a31o_1
XANTENNA_298 _13759_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__10139_ _10139_ VGND VGND VPWR VPWR clknet_0__10139_ sky130_fd_sc_hd__clkbuf_16
X_29258_ _13149_ VGND VGND VPWR VPWR _04398_ sky130_fd_sc_hd__clkbuf_1
X_17272_ _14191_ net2784 _04887_ VGND VGND VPWR VPWR _04897_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19011_ _05671_ _05757_ VGND VGND VPWR VPWR _06345_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16223_ _14467_ VGND VGND VPWR VPWR _01926_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28209_ _12572_ VGND VGND VPWR VPWR _03926_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29189_ _09225_ _11123_ _09230_ VGND VGND VPWR VPWR _13112_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_114_3233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload207 clknet_leaf_201_clk VGND VGND VPWR VPWR clkload207/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_180_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload218 clknet_leaf_173_clk VGND VGND VPWR VPWR clkload218/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_0_3_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload229 clknet_leaf_108_clk VGND VGND VPWR VPWR clkload229/Y sky130_fd_sc_hd__clkinv_1
X_31220_ clknet_leaf_37_clk _02923_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCD\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_588 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16154_ _13172_ VGND VGND VPWR VPWR _14420_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15105_ _13324_ _13649_ VGND VGND VPWR VPWR _13650_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_185_4934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_185_4945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31151_ clknet_leaf_69_clk rvcpu.ALUResultE\[10\] VGND VGND VPWR VPWR rvcpu.dp.plem.ALUResultM\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_16085_ _14383_ VGND VGND VPWR VPWR _01980_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_210_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30102_ net464 _01837_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[11\]\[25\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_75_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15036_ _13559_ _13561_ _13550_ VGND VGND VPWR VPWR _13583_ sky130_fd_sc_hd__a21oi_1
X_19913_ datamem.data_ram\[42\]\[17\] _07203_ _07204_ _07207_ VGND VGND VPWR VPWR
+ _07208_ sky130_fd_sc_hd__o211a_1
X_31082_ clknet_leaf_107_clk _02817_ VGND VGND VPWR VPWR datamem.data_ram\[20\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19844_ datamem.data_ram\[46\]\[1\] _06978_ _07138_ datamem.data_ram\[40\]\[1\] VGND
+ VGND VPWR VPWR _07139_ sky130_fd_sc_hd__a22o_1
X_30033_ net395 _01768_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[13\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_88_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23821__404 clknet_1_0__leaf__10207_ VGND VGND VPWR VPWR net530 sky130_fd_sc_hd__inv_2
X_19775_ _06596_ _07035_ _07069_ VGND VGND VPWR VPWR _07070_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_78_1136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_3952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16987_ net2355 _14470_ _04742_ VGND VGND VPWR VPWR _04746_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_144_3963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18726_ _05610_ _05408_ _05606_ _05429_ _05665_ _05670_ VGND VGND VPWR VPWR _06078_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_155_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15938_ net2510 _13266_ _14297_ VGND VGND VPWR VPWR _14305_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31984_ clknet_leaf_119_clk _03406_ VGND VGND VPWR VPWR datamem.data_ram\[37\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_223_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_3849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_204_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18657_ _05693_ _05820_ _06010_ _05658_ _06012_ VGND VGND VPWR VPWR _06013_ sky130_fd_sc_hd__a221o_1
X_30935_ clknet_leaf_263_clk _02670_ VGND VGND VPWR VPWR datamem.data_ram\[40\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
Xwire37 _07505_ VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_2
X_15869_ net2869 _13269_ _14258_ VGND VGND VPWR VPWR _14267_ sky130_fd_sc_hd__mux2_1
XFILLER_0_204_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17608_ _05075_ VGND VGND VPWR VPWR _01233_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_176_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18588_ _05705_ _05831_ VGND VGND VPWR VPWR _05947_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30866_ clknet_leaf_269_clk _02601_ VGND VGND VPWR VPWR datamem.data_ram\[43\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_32605_ clknet_leaf_240_clk _04027_ VGND VGND VPWR VPWR datamem.data_ram\[20\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_103_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17539_ _13263_ net2504 _05032_ VGND VGND VPWR VPWR _05039_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30797_ clknet_leaf_224_clk _02532_ VGND VGND VPWR VPWR datamem.data_ram\[45\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_43_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20550_ datamem.data_ram\[4\]\[21\] _07837_ _07840_ VGND VGND VPWR VPWR _07841_ sky130_fd_sc_hd__o21a_1
XFILLER_0_62_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32536_ clknet_leaf_183_clk _03958_ VGND VGND VPWR VPWR datamem.data_ram\[23\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_190_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19209_ _06516_ _06517_ VGND VGND VPWR VPWR _06518_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_144_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32467_ clknet_leaf_77_clk _03889_ VGND VGND VPWR VPWR datamem.data_ram\[26\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_20481_ datamem.data_ram\[49\]\[20\] _06782_ _07769_ _07772_ VGND VGND VPWR VPWR
+ _07773_ sky130_fd_sc_hd__o211a_1
XFILLER_0_7_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_717 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22220_ _09385_ VGND VGND VPWR VPWR _09386_ sky130_fd_sc_hd__buf_6
X_31418_ clknet_leaf_103_clk _03121_ VGND VGND VPWR VPWR datamem.data_ram\[15\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_32398_ clknet_leaf_82_clk _03820_ VGND VGND VPWR VPWR datamem.data_ram\[29\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22151_ _09345_ VGND VGND VPWR VPWR _01095_ sky130_fd_sc_hd__clkbuf_1
X_31349_ clknet_leaf_24_clk _03052_ VGND VGND VPWR VPWR rvcpu.dp.hu.ResultSrcE0 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21102_ _06666_ datamem.data_ram\[10\]\[7\] datamem.data_ram\[11\]\[7\] _06944_ _07636_
+ VGND VGND VPWR VPWR _08391_ sky130_fd_sc_hd__o221a_1
XFILLER_0_11_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22082_ rvcpu.dp.plem.WriteDataM\[0\] _08488_ _09293_ _09295_ rvcpu.dp.plem.WriteDataM\[8\]
+ VGND VGND VPWR VPWR _09296_ sky130_fd_sc_hd__a32o_1
XFILLER_0_112_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__10128_ clknet_0__10128_ VGND VGND VPWR VPWR clknet_1_0__leaf__10128_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_1_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25910_ net1838 _11263_ VGND VGND VPWR VPWR _11274_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_1293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21033_ datamem.data_ram\[21\]\[31\] _06721_ _06667_ datamem.data_ram\[23\]\[31\]
+ _06676_ VGND VGND VPWR VPWR _08322_ sky130_fd_sc_hd__o221a_1
XFILLER_0_199_1275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26890_ _11813_ net1395 _11809_ _11817_ VGND VGND VPWR VPWR _03362_ sky130_fd_sc_hd__a31o_1
XFILLER_0_96_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25841_ _11206_ _11207_ _11224_ VGND VGND VPWR VPWR _11225_ sky130_fd_sc_hd__and3_1
XFILLER_0_214_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28560_ _12698_ net3067 _12768_ VGND VGND VPWR VPWR _12774_ sky130_fd_sc_hd__mux2_1
X_25772_ net1890 _11144_ _11147_ _11170_ VGND VGND VPWR VPWR _02891_ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23264__910 clknet_1_1__leaf__10128_ VGND VGND VPWR VPWR net1036 sky130_fd_sc_hd__inv_2
X_27511_ _12157_ net3708 _12179_ VGND VGND VPWR VPWR _12187_ sky130_fd_sc_hd__mux2_1
X_24723_ _10569_ VGND VGND VPWR VPWR _02443_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_215_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28491_ _09231_ net1857 _12724_ VGND VGND VPWR VPWR _12730_ sky130_fd_sc_hd__or3_1
X_21935_ _08795_ _09163_ _09165_ _09167_ VGND VGND VPWR VPWR _09168_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_97_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_222_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_179_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_210_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27442_ _09275_ VGND VGND VPWR VPWR _12147_ sky130_fd_sc_hd__clkbuf_2
X_24654_ _09351_ _10049_ _10052_ VGND VGND VPWR VPWR _10532_ sky130_fd_sc_hd__and3_2
X_21866_ _08835_ _09102_ VGND VGND VPWR VPWR _09103_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20817_ _07829_ _08103_ _08106_ _06751_ VGND VGND VPWR VPWR _08107_ sky130_fd_sc_hd__a211o_1
X_23605_ clknet_1_1__leaf__10172_ VGND VGND VPWR VPWR _10179_ sky130_fd_sc_hd__buf_1
XFILLER_0_33_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27373_ _12095_ net2811 _12097_ VGND VGND VPWR VPWR _12105_ sky130_fd_sc_hd__mux2_1
X_24585_ _10493_ VGND VGND VPWR VPWR _02381_ sky130_fd_sc_hd__clkbuf_1
X_21797_ _08547_ _09035_ _09037_ _08576_ VGND VGND VPWR VPWR _09038_ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29112_ _13071_ VGND VGND VPWR VPWR _04330_ sky130_fd_sc_hd__clkbuf_1
X_26324_ _11495_ VGND VGND VPWR VPWR _11496_ sky130_fd_sc_hd__clkbuf_2
X_20748_ datamem.data_ram\[8\]\[6\] _07829_ VGND VGND VPWR VPWR _08038_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_150_4101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_189_5023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_189_5034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29043_ _10063_ _13031_ VGND VGND VPWR VPWR _13035_ sky130_fd_sc_hd__and2_1
X_26255_ _11458_ VGND VGND VPWR VPWR _03085_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_208_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20679_ _07131_ _07967_ _07969_ VGND VGND VPWR VPWR _07970_ sky130_fd_sc_hd__or3_1
X_22418_ rvcpu.dp.rf.reg_file_arr\[20\]\[6\] rvcpu.dp.rf.reg_file_arr\[21\]\[6\] rvcpu.dp.rf.reg_file_arr\[22\]\[6\]
+ rvcpu.dp.rf.reg_file_arr\[23\]\[6\] _09517_ _09577_ VGND VGND VPWR VPWR _09578_
+ sky130_fd_sc_hd__mux4_2
X_25206_ _10816_ net2268 net56 VGND VGND VPWR VPWR _10842_ sky130_fd_sc_hd__mux2_1
X_26186_ rvcpu.dp.plfd.InstrD\[19\] _11362_ VGND VGND VPWR VPWR _11430_ sky130_fd_sc_hd__and2_1
X_23398_ _09326_ net3585 _10143_ VGND VGND VPWR VPWR _10150_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22349_ _08592_ VGND VGND VPWR VPWR _09512_ sky130_fd_sc_hd__clkbuf_8
X_25137_ _10800_ VGND VGND VPWR VPWR _02626_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_227_5941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_227_5952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_4041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_148_4052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25068_ _09255_ VGND VGND VPWR VPWR _10764_ sky130_fd_sc_hd__buf_2
XFILLER_0_131_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29945_ net315 _01680_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[15\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_223_5838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_223_5849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_4820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16910_ net2766 _14461_ _04695_ VGND VGND VPWR VPWR _04705_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17890_ _05253_ _05258_ _05262_ VGND VGND VPWR VPWR _05263_ sky130_fd_sc_hd__or3b_4
X_29876_ net254 _01611_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[17\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_70_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28827_ _12916_ VGND VGND VPWR VPWR _04200_ sky130_fd_sc_hd__clkbuf_1
X_16841_ _04668_ VGND VGND VPWR VPWR _01617_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_218_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_219_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19560_ datamem.data_ram\[2\]\[24\] _06802_ _06655_ datamem.data_ram\[1\]\[24\] _06732_
+ VGND VGND VPWR VPWR _06856_ sky130_fd_sc_hd__o221a_1
X_16772_ net2265 _14459_ _04623_ VGND VGND VPWR VPWR _04632_ sky130_fd_sc_hd__mux2_1
X_28758_ _12879_ VGND VGND VPWR VPWR _04168_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_107_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18511_ _05789_ _05775_ _05872_ VGND VGND VPWR VPWR _05873_ sky130_fd_sc_hd__and3_1
XFILLER_0_137_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27709_ _12149_ net4000 net50 VGND VGND VPWR VPWR _12293_ sky130_fd_sc_hd__mux2_1
X_15723_ _14186_ VGND VGND VPWR VPWR _02161_ sky130_fd_sc_hd__clkbuf_1
X_19491_ datamem.data_ram\[22\]\[16\] _06630_ _06777_ _06786_ VGND VGND VPWR VPWR
+ _06787_ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28689_ _12737_ net3058 net42 VGND VGND VPWR VPWR _12843_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_178_4760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_178_4771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_940 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_198_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18442_ _05724_ _05733_ VGND VGND VPWR VPWR _05805_ sky130_fd_sc_hd__nor2_2
X_30720_ clknet_leaf_188_clk _02455_ VGND VGND VPWR VPWR datamem.data_ram\[49\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23126__803 clknet_1_0__leaf__10105_ VGND VGND VPWR VPWR net929 sky130_fd_sc_hd__inv_2
X_15654_ _14139_ net3958 _14131_ VGND VGND VPWR VPWR _14140_ sky130_fd_sc_hd__mux2_1
XFILLER_0_185_422 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_197_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_185_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14605_ net2483 _13187_ _13181_ VGND VGND VPWR VPWR _13188_ sky130_fd_sc_hd__mux2_1
XFILLER_0_200_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_174_4668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18373_ _05661_ _05695_ _05718_ _05737_ VGND VGND VPWR VPWR _05738_ sky130_fd_sc_hd__a211o_1
XFILLER_0_139_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30651_ clknet_leaf_178_clk _02386_ VGND VGND VPWR VPWR datamem.data_ram\[51\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_174_4679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15585_ net2148 _13204_ _14092_ VGND VGND VPWR VPWR _14100_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_1278 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17324_ _04925_ VGND VGND VPWR VPWR _01383_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30582_ clknet_leaf_191_clk _02317_ VGND VGND VPWR VPWR datamem.data_ram\[53\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32321_ clknet_leaf_77_clk _03743_ VGND VGND VPWR VPWR datamem.data_ram\[31\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17255_ _04888_ VGND VGND VPWR VPWR _01415_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16206_ net2873 _14455_ _14443_ VGND VGND VPWR VPWR _14456_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32252_ clknet_leaf_168_clk _03674_ VGND VGND VPWR VPWR datamem.data_ram\[34\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_77_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17186_ _14172_ net2534 _04851_ VGND VGND VPWR VPWR _04852_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_180_Right_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_133_3686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31203_ clknet_leaf_27_clk _02906_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCPlus4D\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_133_3697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16137_ _14411_ VGND VGND VPWR VPWR _01956_ sky130_fd_sc_hd__clkbuf_1
X_32183_ clknet_leaf_89_clk _03605_ VGND VGND VPWR VPWR datamem.data_ram\[37\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_31134_ clknet_leaf_211_clk _02869_ VGND VGND VPWR VPWR datamem.data_ram\[4\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3208 datamem.data_ram\[26\]\[14\] VGND VGND VPWR VPWR net4358 sky130_fd_sc_hd__dlygate4sd3_1
X_16068_ net2023 _13254_ _14371_ VGND VGND VPWR VPWR _14375_ sky130_fd_sc_hd__mux2_1
Xhold3219 datamem.data_ram\[57\]\[17\] VGND VGND VPWR VPWR net4369 sky130_fd_sc_hd__dlygate4sd3_1
X_15019_ _13403_ _13523_ _13561_ VGND VGND VPWR VPWR _13567_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2507 datamem.data_ram\[46\]\[9\] VGND VGND VPWR VPWR net3657 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_36_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31065_ clknet_leaf_286_clk _02800_ VGND VGND VPWR VPWR datamem.data_ram\[8\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2518 datamem.data_ram\[47\]\[15\] VGND VGND VPWR VPWR net3668 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_36_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23745__335 clknet_1_1__leaf__10200_ VGND VGND VPWR VPWR net461 sky130_fd_sc_hd__inv_2
Xhold2529 datamem.data_ram\[45\]\[13\] VGND VGND VPWR VPWR net3679 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30016_ net378 _01751_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[13\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19827_ _06990_ VGND VGND VPWR VPWR _07122_ sky130_fd_sc_hd__clkbuf_8
X_23213__864 clknet_1_0__leaf__10112_ VGND VGND VPWR VPWR net990 sky130_fd_sc_hd__inv_2
Xhold1806 rvcpu.dp.rf.reg_file_arr\[22\]\[5\] VGND VGND VPWR VPWR net2956 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1817 datamem.data_ram\[37\]\[16\] VGND VGND VPWR VPWR net2967 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1828 datamem.data_ram\[36\]\[28\] VGND VGND VPWR VPWR net2978 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_16_Left_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1839 rvcpu.dp.rf.reg_file_arr\[19\]\[16\] VGND VGND VPWR VPWR net2989 sky130_fd_sc_hd__dlygate4sd3_1
X_19758_ datamem.data_ram\[54\]\[25\] _06719_ _06671_ datamem.data_ram\[55\]\[25\]
+ VGND VGND VPWR VPWR _07053_ sky130_fd_sc_hd__o22a_1
XFILLER_0_56_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18709_ _05990_ _05903_ _06060_ _06061_ VGND VGND VPWR VPWR _06062_ sky130_fd_sc_hd__o211ai_1
X_31967_ clknet_leaf_130_clk _03389_ VGND VGND VPWR VPWR datamem.data_ram\[54\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_19689_ _06860_ VGND VGND VPWR VPWR _06985_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_56_1242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_189_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24171__13 clknet_1_0__leaf__10264_ VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__inv_2
X_21720_ rvcpu.dp.rf.reg_file_arr\[12\]\[17\] rvcpu.dp.rf.reg_file_arr\[13\]\[17\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[17\] rvcpu.dp.rf.reg_file_arr\[15\]\[17\] _08839_
+ _08840_ VGND VGND VPWR VPWR _08965_ sky130_fd_sc_hd__mux4_2
XFILLER_0_176_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30918_ clknet_leaf_228_clk _02653_ VGND VGND VPWR VPWR datamem.data_ram\[40\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31898_ _04440_ net120 VGND VGND VPWR VPWR datamem.rd_data_mem\[3\] sky130_fd_sc_hd__dlxtn_1
XTAP_TAPCELL_ROW_101_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21651_ _08899_ VGND VGND VPWR VPWR _01041_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_606 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30849_ clknet_leaf_220_clk _02584_ VGND VGND VPWR VPWR datamem.data_ram\[43\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20602_ _07872_ _07879_ _07885_ _07177_ _07892_ VGND VGND VPWR VPWR _07893_ sky130_fd_sc_hd__o221a_1
X_24370_ _09322_ net3311 net61 VGND VGND VPWR VPWR _10363_ sky130_fd_sc_hd__mux2_1
X_21582_ rvcpu.dp.rf.reg_file_arr\[4\]\[10\] rvcpu.dp.rf.reg_file_arr\[5\]\[10\] rvcpu.dp.rf.reg_file_arr\[6\]\[10\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[10\] _08551_ _08555_ VGND VGND VPWR VPWR _08834_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_19_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_25_Left_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20533_ _06652_ VGND VGND VPWR VPWR _07824_ sky130_fd_sc_hd__buf_8
X_32519_ clknet_leaf_74_clk _03941_ VGND VGND VPWR VPWR datamem.data_ram\[24\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23294__936 clknet_1_0__leaf__10132_ VGND VGND VPWR VPWR net1062 sky130_fd_sc_hd__inv_2
XFILLER_0_90_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26040_ _11091_ _11340_ VGND VGND VPWR VPWR _11347_ sky130_fd_sc_hd__and2_1
XFILLER_0_131_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20464_ datamem.data_ram\[20\]\[20\] _07230_ _07755_ _06679_ VGND VGND VPWR VPWR
+ _07756_ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22203_ _09374_ VGND VGND VPWR VPWR _01118_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20395_ datamem.data_ram\[24\]\[28\] _06695_ _06730_ datamem.data_ram\[27\]\[28\]
+ _07686_ VGND VGND VPWR VPWR _07687_ sky130_fd_sc_hd__o221a_1
X_24125__631 clknet_1_0__leaf__10260_ VGND VGND VPWR VPWR net757 sky130_fd_sc_hd__inv_2
X_22134_ _09336_ VGND VGND VPWR VPWR _01087_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_219_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27991_ _12454_ net3667 net76 VGND VGND VPWR VPWR _12455_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29730_ net1076 _01465_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[22\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_26942_ _11849_ net1609 _11841_ _11851_ VGND VGND VPWR VPWR _03380_ sky130_fd_sc_hd__a31o_1
X_22065_ _09282_ net3819 _09270_ VGND VGND VPWR VPWR _09283_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_34_Left_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21016_ datamem.data_ram\[58\]\[31\] _06802_ _06780_ datamem.data_ram\[57\]\[31\]
+ _08304_ VGND VGND VPWR VPWR _08305_ sky130_fd_sc_hd__o221a_1
X_29661_ net1007 _01396_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[24\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26873_ _11672_ _11798_ VGND VGND VPWR VPWR _11807_ sky130_fd_sc_hd__and2_1
XFILLER_0_199_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28612_ _12698_ net3072 _12796_ VGND VGND VPWR VPWR _12802_ sky130_fd_sc_hd__mux2_1
X_25824_ rvcpu.dp.plfd.PCPlus4D\[21\] _11210_ _11142_ VGND VGND VPWR VPWR _11211_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_173_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_199_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29592_ net946 _01327_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[26\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_28543_ _09255_ VGND VGND VPWR VPWR _12764_ sky130_fd_sc_hd__buf_2
X_25755_ _13865_ _11157_ _13758_ VGND VGND VPWR VPWR _11158_ sky130_fd_sc_hd__or3b_1
XFILLER_0_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24706_ _10560_ VGND VGND VPWR VPWR _02435_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21918_ rvcpu.dp.rf.reg_file_arr\[0\]\[28\] rvcpu.dp.rf.reg_file_arr\[1\]\[28\] rvcpu.dp.rf.reg_file_arr\[2\]\[28\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[28\] _08810_ _08811_ VGND VGND VPWR VPWR _09152_
+ sky130_fd_sc_hd__mux4_1
X_28474_ _12719_ VGND VGND VPWR VPWR _04044_ sky130_fd_sc_hd__clkbuf_1
X_25686_ _11081_ _11113_ VGND VGND VPWR VPWR _11115_ sky130_fd_sc_hd__and2_1
XFILLER_0_139_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22898_ rvcpu.dp.rf.reg_file_arr\[4\]\[31\] rvcpu.dp.rf.reg_file_arr\[5\]\[31\] rvcpu.dp.rf.reg_file_arr\[6\]\[31\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[31\] _09416_ _09418_ VGND VGND VPWR VPWR _10033_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_167_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27425_ _12135_ VGND VGND VPWR VPWR _03579_ sky130_fd_sc_hd__clkbuf_1
X_24637_ _10522_ VGND VGND VPWR VPWR _02404_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_214_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21849_ _08682_ _09084_ _09086_ _08558_ VGND VGND VPWR VPWR _09087_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_216_5675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_216_5686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_43_Left_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15370_ _13368_ _13646_ _13793_ _13521_ VGND VGND VPWR VPWR _13904_ sky130_fd_sc_hd__a31oi_1
X_27356_ _12095_ net2700 _12081_ VGND VGND VPWR VPWR _12096_ sky130_fd_sc_hd__mux2_1
X_24568_ _10484_ VGND VGND VPWR VPWR _02373_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26307_ _11486_ VGND VGND VPWR VPWR _03110_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_182_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23519_ _09252_ net2857 _10162_ VGND VGND VPWR VPWR _10168_ sky130_fd_sc_hd__mux2_1
X_27287_ _12036_ net1556 _12053_ _12056_ VGND VGND VPWR VPWR _03520_ sky130_fd_sc_hd__a31o_1
X_24499_ _10439_ net4427 _10440_ VGND VGND VPWR VPWR _10441_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17040_ _04774_ VGND VGND VPWR VPWR _01516_ sky130_fd_sc_hd__clkbuf_1
X_29026_ _12743_ net3449 net66 VGND VGND VPWR VPWR _13025_ sky130_fd_sc_hd__mux2_1
X_26238_ _11379_ _03044_ _11454_ VGND VGND VPWR VPWR _03071_ sky130_fd_sc_hd__a21o_1
XFILLER_0_135_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23156__829 clknet_1_1__leaf__10109_ VGND VGND VPWR VPWR net955 sky130_fd_sc_hd__inv_2
X_26169_ _11421_ VGND VGND VPWR VPWR _03037_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18991_ _05298_ _05785_ VGND VGND VPWR VPWR _06326_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_221_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_4494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_52_Left_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17942_ rvcpu.dp.plde.ImmExtE\[15\] rvcpu.dp.SrcBFW_Mux.y\[15\] _05277_ VGND VGND
+ VPWR VPWR _05314_ sky130_fd_sc_hd__mux2_1
X_29928_ net298 _01663_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[16\]\[19\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_109_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17873_ rvcpu.dp.plde.Rs1E\[2\] rvcpu.dp.plem.RdM\[2\] VGND VGND VPWR VPWR _05246_
+ sky130_fd_sc_hd__xnor2_1
X_29859_ net237 _01594_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[18\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16824_ net1889 _14442_ _04659_ VGND VGND VPWR VPWR _04660_ sky130_fd_sc_hd__mux2_1
X_19612_ _06712_ _06886_ _06897_ _06797_ _06907_ VGND VGND VPWR VPWR _06908_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_105_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32870_ clknet_leaf_282_clk _04292_ VGND VGND VPWR VPWR datamem.data_ram\[11\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_194 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31821_ clknet_leaf_104_clk _03275_ VGND VGND VPWR VPWR datamem.data_ram\[9\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19543_ datamem.data_ram\[30\]\[24\] _06717_ _06812_ datamem.data_ram\[27\]\[24\]
+ VGND VGND VPWR VPWR _06839_ sky130_fd_sc_hd__o22a_1
XFILLER_0_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_176_4708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16755_ _04611_ VGND VGND VPWR VPWR _04623_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_176_4719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_1197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15706_ _13247_ VGND VGND VPWR VPWR _14175_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_66_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31752_ clknet_leaf_61_clk _03206_ VGND VGND VPWR VPWR datamem.data_ram\[45\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_19474_ datamem.data_ram\[50\]\[16\] _06728_ _06768_ datamem.data_ram\[53\]\[16\]
+ _06769_ VGND VGND VPWR VPWR _06770_ sky130_fd_sc_hd__o221a_1
XFILLER_0_76_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16686_ _04586_ VGND VGND VPWR VPWR _01698_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18425_ rvcpu.dp.plde.ALUControlE\[2\] rvcpu.dp.plde.ALUControlE\[3\] rvcpu.dp.plde.ALUControlE\[1\]
+ rvcpu.dp.plde.ALUControlE\[0\] VGND VGND VPWR VPWR _05789_ sky130_fd_sc_hd__and4b_1
X_30703_ clknet_leaf_197_clk _02438_ VGND VGND VPWR VPWR datamem.data_ram\[49\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_61_Left_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15637_ _13172_ VGND VGND VPWR VPWR _14127_ sky130_fd_sc_hd__buf_4
X_31683_ clknet_leaf_8_clk net1303 VGND VGND VPWR VPWR rvcpu.dp.plmw.ALUResultW\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_139_3840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_185_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_1195 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18356_ _05719_ _05720_ VGND VGND VPWR VPWR _05721_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_29_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30634_ clknet_leaf_219_clk _02369_ VGND VGND VPWR VPWR datamem.data_ram\[51\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_15568_ rvcpu.dp.plmw.RegWriteW rvcpu.dp.plmw.RdW\[0\] rvcpu.dp.plmw.RdW\[1\] VGND
+ VGND VPWR VPWR _14090_ sky130_fd_sc_hd__nand3_4
XFILLER_0_51_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_3726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_3737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17307_ _04916_ VGND VGND VPWR VPWR _01391_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18287_ rvcpu.dp.plde.ALUControlE\[0\] VGND VGND VPWR VPWR _05652_ sky130_fd_sc_hd__inv_2
X_30565_ clknet_leaf_143_clk _02300_ VGND VGND VPWR VPWR datamem.data_ram\[54\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15499_ _13370_ _13348_ _13505_ _13425_ _13374_ VGND VGND VPWR VPWR _14027_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_25_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32304_ clknet_leaf_168_clk _03726_ VGND VGND VPWR VPWR datamem.data_ram\[32\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17238_ _04879_ VGND VGND VPWR VPWR _01423_ sky130_fd_sc_hd__clkbuf_1
X_30496_ clknet_leaf_143_clk _02231_ VGND VGND VPWR VPWR datamem.data_ram\[57\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32235_ clknet_leaf_242_clk _03657_ VGND VGND VPWR VPWR datamem.data_ram\[35\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold903 rvcpu.dp.rf.reg_file_arr\[5\]\[19\] VGND VGND VPWR VPWR net2053 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23450__100 clknet_1_0__leaf__10156_ VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__inv_2
X_17169_ _14156_ net4288 _04840_ VGND VGND VPWR VPWR _04843_ sky130_fd_sc_hd__mux2_1
Xhold914 rvcpu.dp.rf.reg_file_arr\[9\]\[24\] VGND VGND VPWR VPWR net2064 sky130_fd_sc_hd__dlygate4sd3_1
Xhold925 rvcpu.dp.rf.reg_file_arr\[18\]\[13\] VGND VGND VPWR VPWR net2075 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold936 rvcpu.dp.rf.reg_file_arr\[7\]\[8\] VGND VGND VPWR VPWR net2086 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold947 rvcpu.dp.rf.reg_file_arr\[30\]\[16\] VGND VGND VPWR VPWR net2097 sky130_fd_sc_hd__dlygate4sd3_1
Xhold958 rvcpu.dp.rf.reg_file_arr\[10\]\[4\] VGND VGND VPWR VPWR net2108 sky130_fd_sc_hd__dlygate4sd3_1
X_20180_ datamem.data_ram\[13\]\[11\] _06702_ _06778_ datamem.data_ram\[8\]\[11\]
+ VGND VGND VPWR VPWR _07473_ sky130_fd_sc_hd__o22a_1
X_32166_ clknet_leaf_277_clk _03588_ VGND VGND VPWR VPWR datamem.data_ram\[38\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold969 rvcpu.dp.rf.reg_file_arr\[6\]\[25\] VGND VGND VPWR VPWR net2119 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3005 datamem.data_ram\[48\]\[17\] VGND VGND VPWR VPWR net4155 sky130_fd_sc_hd__dlygate4sd3_1
X_23669__266 clknet_1_0__leaf__10193_ VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__inv_2
XFILLER_0_177_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3016 rvcpu.dp.rf.reg_file_arr\[26\]\[3\] VGND VGND VPWR VPWR net4166 sky130_fd_sc_hd__dlygate4sd3_1
X_31117_ clknet_leaf_109_clk _02852_ VGND VGND VPWR VPWR datamem.data_ram\[35\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3027 datamem.data_ram\[32\]\[15\] VGND VGND VPWR VPWR net4177 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3038 datamem.data_ram\[15\]\[13\] VGND VGND VPWR VPWR net4188 sky130_fd_sc_hd__dlygate4sd3_1
X_32097_ clknet_leaf_107_clk _03519_ VGND VGND VPWR VPWR datamem.data_ram\[23\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2304 datamem.data_ram\[12\]\[20\] VGND VGND VPWR VPWR net3454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3049 rvcpu.dp.rf.reg_file_arr\[16\]\[3\] VGND VGND VPWR VPWR net4199 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2315 datamem.data_ram\[12\]\[25\] VGND VGND VPWR VPWR net3465 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2326 datamem.data_ram\[36\]\[24\] VGND VGND VPWR VPWR net3476 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2337 rvcpu.dp.rf.reg_file_arr\[13\]\[28\] VGND VGND VPWR VPWR net3487 sky130_fd_sc_hd__dlygate4sd3_1
X_31048_ clknet_leaf_234_clk _02783_ VGND VGND VPWR VPWR datamem.data_ram\[9\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_209_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2348 datamem.data_ram\[16\]\[11\] VGND VGND VPWR VPWR net3498 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1603 datamem.data_ram\[56\]\[24\] VGND VGND VPWR VPWR net2753 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1614 datamem.data_ram\[3\]\[26\] VGND VGND VPWR VPWR net2764 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2359 rvcpu.dp.rf.reg_file_arr\[26\]\[26\] VGND VGND VPWR VPWR net3509 sky130_fd_sc_hd__dlygate4sd3_1
X_26508__60 clknet_1_0__leaf__11602_ VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__inv_2
Xhold1625 rvcpu.dp.rf.reg_file_arr\[5\]\[4\] VGND VGND VPWR VPWR net2775 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1636 rvcpu.dp.rf.reg_file_arr\[1\]\[5\] VGND VGND VPWR VPWR net2786 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1647 datamem.data_ram\[13\]\[20\] VGND VGND VPWR VPWR net2797 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_193_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1658 datamem.data_ram\[32\]\[9\] VGND VGND VPWR VPWR net2808 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1669 datamem.data_ram\[10\]\[18\] VGND VGND VPWR VPWR net2819 sky130_fd_sc_hd__dlygate4sd3_1
X_22821_ _09954_ _09956_ _09959_ _09411_ _09525_ VGND VGND VPWR VPWR _09960_ sky130_fd_sc_hd__a221o_1
XFILLER_0_168_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_196_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25540_ _10737_ net3000 _11021_ VGND VGND VPWR VPWR _11028_ sky130_fd_sc_hd__mux2_1
X_22752_ _09433_ _09894_ _09789_ VGND VGND VPWR VPWR _09895_ sky130_fd_sc_hd__a21o_1
XFILLER_0_17_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21703_ rvcpu.dp.rf.reg_file_arr\[0\]\[16\] rvcpu.dp.rf.reg_file_arr\[1\]\[16\] rvcpu.dp.rf.reg_file_arr\[2\]\[16\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[16\] _08566_ _08569_ VGND VGND VPWR VPWR _08949_
+ sky130_fd_sc_hd__mux4_1
X_25471_ _10416_ _10985_ VGND VGND VPWR VPWR _10992_ sky130_fd_sc_hd__and2_1
XFILLER_0_149_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22683_ _09627_ _09827_ _09829_ _09795_ VGND VGND VPWR VPWR _09830_ sky130_fd_sc_hd__a211o_1
XFILLER_0_137_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27210_ _11978_ _12008_ VGND VGND VPWR VPWR _12015_ sky130_fd_sc_hd__and2_1
XFILLER_0_177_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_176_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_639 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21634_ _08514_ _08882_ VGND VGND VPWR VPWR _08883_ sky130_fd_sc_hd__or2_1
X_24422_ _10392_ net4378 _10386_ VGND VGND VPWR VPWR _10393_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28190_ _12562_ VGND VGND VPWR VPWR _03917_ sky130_fd_sc_hd__clkbuf_1
X_27141_ _11972_ _11966_ VGND VGND VPWR VPWR _11973_ sky130_fd_sc_hd__and2_1
XFILLER_0_191_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_272 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21565_ _08525_ VGND VGND VPWR VPWR _08818_ sky130_fd_sc_hd__buf_4
X_24353_ _09285_ net4356 _10348_ VGND VGND VPWR VPWR _10354_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_211_5550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23914__471 clknet_1_0__leaf__10225_ VGND VGND VPWR VPWR net597 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_211_5561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_191_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20516_ _07071_ _07790_ _07796_ _07801_ _07806_ VGND VGND VPWR VPWR _07807_ sky130_fd_sc_hd__o32a_2
XFILLER_0_133_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27072_ _11803_ _11924_ VGND VGND VPWR VPWR _11929_ sky130_fd_sc_hd__and2_1
XFILLER_0_133_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24284_ _09260_ net2394 _10307_ VGND VGND VPWR VPWR _10315_ sky130_fd_sc_hd__mux2_1
X_21496_ rvcpu.dp.rf.reg_file_arr\[12\]\[6\] rvcpu.dp.rf.reg_file_arr\[13\]\[6\] rvcpu.dp.rf.reg_file_arr\[14\]\[6\]
+ rvcpu.dp.rf.reg_file_arr\[15\]\[6\] _08551_ _08555_ VGND VGND VPWR VPWR _08752_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_160_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26023_ net26 _11152_ VGND VGND VPWR VPWR _11337_ sky130_fd_sc_hd__or2_1
X_23613__232 clknet_1_0__leaf__10179_ VGND VGND VPWR VPWR net358 sky130_fd_sc_hd__inv_2
XFILLER_0_166_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20447_ datamem.data_ram\[6\]\[20\] _06764_ _06779_ datamem.data_ram\[0\]\[20\] _07738_
+ VGND VGND VPWR VPWR _07739_ sky130_fd_sc_hd__o221a_1
XFILLER_0_31_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20378_ datamem.data_ram\[61\]\[28\] _06660_ _06653_ datamem.data_ram\[57\]\[28\]
+ VGND VGND VPWR VPWR _07670_ sky130_fd_sc_hd__o22a_1
X_22117_ rvcpu.dp.plem.WriteDataM\[30\] _09221_ _09295_ rvcpu.dp.plem.WriteDataM\[14\]
+ _09324_ VGND VGND VPWR VPWR _09325_ sky130_fd_sc_hd__a221o_4
X_27974_ _09255_ VGND VGND VPWR VPWR _12443_ sky130_fd_sc_hd__clkbuf_2
X_29713_ net1059 _01448_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[22\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_26925_ _10325_ _08059_ _11609_ VGND VGND VPWR VPWR _11842_ sky130_fd_sc_hd__and3_2
X_22048_ _09226_ _09269_ _09231_ VGND VGND VPWR VPWR _09270_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_162_4380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_4391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29644_ net990 _01379_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[24\]\[7\] sky130_fd_sc_hd__dfxtp_1
Xhold2860 rvcpu.dp.rf.reg_file_arr\[17\]\[19\] VGND VGND VPWR VPWR net4010 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_214_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14870_ _13313_ _13331_ VGND VGND VPWR VPWR _13422_ sky130_fd_sc_hd__or2_2
X_26856_ _11796_ VGND VGND VPWR VPWR _11797_ sky130_fd_sc_hd__buf_2
Xhold2871 datamem.data_ram\[21\]\[21\] VGND VGND VPWR VPWR net4021 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2882 rvcpu.dp.rf.reg_file_arr\[26\]\[28\] VGND VGND VPWR VPWR net4032 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2893 datamem.data_ram\[61\]\[16\] VGND VGND VPWR VPWR net4043 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25807_ rvcpu.dp.pcreg.q\[18\] rvcpu.dp.pcreg.q\[17\] _11191_ VGND VGND VPWR VPWR
+ _11197_ sky130_fd_sc_hd__and3_1
X_29575_ net929 _01310_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[26\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_214_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26787_ _11645_ _11749_ VGND VGND VPWR VPWR _11756_ sky130_fd_sc_hd__and2_1
XFILLER_0_98_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_218_5726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_218_5737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28526_ _12751_ net2850 _12752_ VGND VGND VPWR VPWR _12753_ sky130_fd_sc_hd__mux2_1
X_16540_ _14141_ net3162 _04503_ VGND VGND VPWR VPWR _04509_ sky130_fd_sc_hd__mux2_1
X_25738_ _11143_ VGND VGND VPWR VPWR _11144_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_134_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_731 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28457_ _12710_ VGND VGND VPWR VPWR _04036_ sky130_fd_sc_hd__clkbuf_1
X_16471_ _04472_ VGND VGND VPWR VPWR _01807_ sky130_fd_sc_hd__clkbuf_1
X_25669_ _11047_ _11098_ VGND VGND VPWR VPWR _11103_ sky130_fd_sc_hd__and2_1
XFILLER_0_195_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_171_4605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18210_ _05384_ _05385_ _05388_ VGND VGND VPWR VPWR _05575_ sky130_fd_sc_hd__a21o_1
X_15422_ _13324_ _13649_ _13953_ VGND VGND VPWR VPWR _13954_ sky130_fd_sc_hd__o21ai_1
X_27408_ _12095_ net2305 _12116_ VGND VGND VPWR VPWR _12124_ sky130_fd_sc_hd__mux2_1
X_19190_ rvcpu.dp.plde.ImmExtE\[22\] rvcpu.dp.plde.PCE\[22\] VGND VGND VPWR VPWR _06501_
+ sky130_fd_sc_hd__nand2_1
X_28388_ _12670_ VGND VGND VPWR VPWR _04007_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18141_ _13228_ rvcpu.dp.plde.RD2E\[16\] _05195_ VGND VGND VPWR VPWR _05507_ sky130_fd_sc_hd__mux2_1
X_23242__890 clknet_1_0__leaf__10126_ VGND VGND VPWR VPWR net1016 sky130_fd_sc_hd__inv_2
X_15353_ _13693_ _13780_ _13435_ _13581_ VGND VGND VPWR VPWR _13888_ sky130_fd_sc_hd__a211o_1
X_27339_ _12084_ VGND VGND VPWR VPWR _03544_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18072_ _05439_ VGND VGND VPWR VPWR _05440_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30350_ net696 _02085_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[3\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_15284_ _13419_ _13370_ _13496_ _13469_ VGND VGND VPWR VPWR _13822_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_130_3612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29009_ _12995_ net1610 _13009_ _13015_ VGND VGND VPWR VPWR _04283_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_169_4545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_130_3623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17023_ _04765_ VGND VGND VPWR VPWR _01524_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_169_4556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30281_ clknet_leaf_145_clk _02016_ VGND VGND VPWR VPWR datamem.data_ram\[58\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_1230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32020_ clknet_leaf_129_clk _03442_ VGND VGND VPWR VPWR datamem.data_ram\[51\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_221_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18974_ _05300_ _05539_ _05545_ _05527_ _05666_ _05671_ VGND VGND VPWR VPWR _06310_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_219_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17925_ _05296_ _05297_ VGND VGND VPWR VPWR _05298_ sky130_fd_sc_hd__nor2_2
XFILLER_0_225_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_3563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_3574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17856_ _13256_ rvcpu.dp.plde.RD2E\[7\] _05195_ VGND VGND VPWR VPWR _05232_ sky130_fd_sc_hd__mux2_1
X_32922_ clknet_leaf_272_clk _04344_ VGND VGND VPWR VPWR datamem.data_ram\[0\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_16807_ net1927 _14426_ _04648_ VGND VGND VPWR VPWR _04651_ sky130_fd_sc_hd__mux2_1
X_24074__600 clknet_1_1__leaf__10248_ VGND VGND VPWR VPWR net726 sky130_fd_sc_hd__inv_2
X_17787_ _13271_ _05179_ _05180_ VGND VGND VPWR VPWR _05183_ sky130_fd_sc_hd__nand3b_1
XTAP_TAPCELL_ROW_50_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32853_ clknet_leaf_237_clk _04275_ VGND VGND VPWR VPWR datamem.data_ram\[11\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_14999_ _13303_ _13321_ _13546_ _13331_ VGND VGND VPWR VPWR _13547_ sky130_fd_sc_hd__o31a_1
XFILLER_0_205_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31804_ clknet_leaf_98_clk _03258_ VGND VGND VPWR VPWR datamem.data_ram\[46\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19526_ datamem.data_ram\[40\]\[24\] _06821_ _06805_ datamem.data_ram\[44\]\[24\]
+ VGND VGND VPWR VPWR _06822_ sky130_fd_sc_hd__o22a_1
X_16738_ _04614_ VGND VGND VPWR VPWR _01674_ sky130_fd_sc_hd__clkbuf_1
X_32784_ clknet_leaf_177_clk _04206_ VGND VGND VPWR VPWR datamem.data_ram\[14\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19457_ _06752_ VGND VGND VPWR VPWR _06753_ sky130_fd_sc_hd__buf_6
X_31735_ net184 _03193_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[9\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16669_ _14133_ net2199 _04576_ VGND VGND VPWR VPWR _04578_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18408_ _05666_ _05771_ VGND VGND VPWR VPWR _05772_ sky130_fd_sc_hd__nor2_1
X_31666_ clknet_leaf_66_clk net1281 VGND VGND VPWR VPWR rvcpu.dp.plmw.ALUResultW\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_19388_ _06616_ VGND VGND VPWR VPWR _06684_ sky130_fd_sc_hd__buf_6
XFILLER_0_5_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23024__726 clknet_1_0__leaf__10088_ VGND VGND VPWR VPWR net852 sky130_fd_sc_hd__inv_2
X_18339_ _05398_ VGND VGND VPWR VPWR _05704_ sky130_fd_sc_hd__buf_2
X_30617_ clknet_leaf_147_clk _02352_ VGND VGND VPWR VPWR datamem.data_ram\[52\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31597_ clknet_leaf_48_clk net1233 VGND VGND VPWR VPWR rvcpu.dp.plmw.PCPlus4W\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_21350_ rvcpu.dp.plde.funct3E\[2\] rvcpu.dp.plde.funct3E\[1\] _08611_ rvcpu.dp.plde.funct3E\[0\]
+ VGND VGND VPWR VPWR _08612_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_127_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30548_ clknet_leaf_146_clk _02283_ VGND VGND VPWR VPWR datamem.data_ram\[55\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_23104__783 clknet_1_1__leaf__10103_ VGND VGND VPWR VPWR net909 sky130_fd_sc_hd__inv_2
X_20301_ datamem.data_ram\[0\]\[19\] _06698_ _07590_ _07593_ VGND VGND VPWR VPWR _07594_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_13_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold700 datamem.data_ram\[52\]\[1\] VGND VGND VPWR VPWR net1850 sky130_fd_sc_hd__dlygate4sd3_1
X_21281_ rvcpu.dp.rf.reg_file_arr\[24\]\[0\] rvcpu.dp.rf.reg_file_arr\[25\]\[0\] rvcpu.dp.rf.reg_file_arr\[26\]\[0\]
+ rvcpu.dp.rf.reg_file_arr\[27\]\[0\] _08525_ _08528_ VGND VGND VPWR VPWR _08543_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_4_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30479_ net157 _02214_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[19\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold711 datamem.data_ram\[35\]\[0\] VGND VGND VPWR VPWR net1861 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold722 rvcpu.dp.rf.reg_file_arr\[10\]\[10\] VGND VGND VPWR VPWR net1872 sky130_fd_sc_hd__dlygate4sd3_1
X_20232_ datamem.data_ram\[5\]\[3\] _06919_ _06936_ datamem.data_ram\[0\]\[3\] _06741_
+ VGND VGND VPWR VPWR _07525_ sky130_fd_sc_hd__a221o_1
XFILLER_0_163_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32218_ clknet_leaf_229_clk _03640_ VGND VGND VPWR VPWR datamem.data_ram\[35\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold733 rvcpu.dp.rf.reg_file_arr\[18\]\[4\] VGND VGND VPWR VPWR net1883 sky130_fd_sc_hd__dlygate4sd3_1
Xhold744 datamem.data_ram\[36\]\[31\] VGND VGND VPWR VPWR net1894 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold755 rvcpu.dp.rf.reg_file_arr\[11\]\[11\] VGND VGND VPWR VPWR net1905 sky130_fd_sc_hd__dlygate4sd3_1
Xhold766 datamem.data_ram\[53\]\[4\] VGND VGND VPWR VPWR net1916 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold777 rvcpu.dp.rf.reg_file_arr\[17\]\[29\] VGND VGND VPWR VPWR net1927 sky130_fd_sc_hd__dlygate4sd3_1
Xhold788 datamem.data_ram\[4\]\[15\] VGND VGND VPWR VPWR net1938 sky130_fd_sc_hd__dlygate4sd3_1
X_32149_ clknet_leaf_225_clk _03571_ VGND VGND VPWR VPWR datamem.data_ram\[38\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_20163_ datamem.data_ram\[19\]\[27\] _06730_ _06765_ datamem.data_ram\[20\]\[27\]
+ _06732_ VGND VGND VPWR VPWR _07456_ sky130_fd_sc_hd__o221a_1
Xhold799 datamem.data_ram\[50\]\[30\] VGND VGND VPWR VPWR net1949 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2101 datamem.data_ram\[60\]\[11\] VGND VGND VPWR VPWR net3251 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2112 rvcpu.dp.rf.reg_file_arr\[15\]\[12\] VGND VGND VPWR VPWR net3262 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2123 rvcpu.dp.rf.reg_file_arr\[22\]\[24\] VGND VGND VPWR VPWR net3273 sky130_fd_sc_hd__dlygate4sd3_1
X_24971_ _10500_ VGND VGND VPWR VPWR _10705_ sky130_fd_sc_hd__buf_6
X_20094_ datamem.data_ram\[57\]\[10\] _06790_ _07384_ _07387_ VGND VGND VPWR VPWR
+ _07388_ sky130_fd_sc_hd__o211a_1
XFILLER_0_228_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2134 datamem.data_ram\[53\]\[29\] VGND VGND VPWR VPWR net3284 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2145 datamem.data_ram\[13\]\[23\] VGND VGND VPWR VPWR net3295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1400 datamem.data_ram\[62\]\[25\] VGND VGND VPWR VPWR net2550 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1411 datamem.data_ram\[17\]\[23\] VGND VGND VPWR VPWR net2561 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2156 rvcpu.dp.rf.reg_file_arr\[11\]\[19\] VGND VGND VPWR VPWR net3306 sky130_fd_sc_hd__dlygate4sd3_1
X_26710_ _10822_ net3831 _11704_ VGND VGND VPWR VPWR _11710_ sky130_fd_sc_hd__mux2_1
Xhold2167 datamem.data_ram\[50\]\[21\] VGND VGND VPWR VPWR net3317 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1422 datamem.data_ram\[50\]\[24\] VGND VGND VPWR VPWR net2572 sky130_fd_sc_hd__dlygate4sd3_1
X_27690_ _12130_ net2809 _12280_ VGND VGND VPWR VPWR _12283_ sky130_fd_sc_hd__mux2_1
Xhold1433 rvcpu.dp.rf.reg_file_arr\[6\]\[27\] VGND VGND VPWR VPWR net2583 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2178 datamem.data_ram\[33\]\[30\] VGND VGND VPWR VPWR net3328 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2189 datamem.data_ram\[2\]\[21\] VGND VGND VPWR VPWR net3339 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1444 datamem.data_ram\[55\]\[12\] VGND VGND VPWR VPWR net2594 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1455 datamem.data_ram\[51\]\[19\] VGND VGND VPWR VPWR net2605 sky130_fd_sc_hd__dlygate4sd3_1
X_26641_ _11665_ net1708 _11662_ _11667_ VGND VGND VPWR VPWR _03263_ sky130_fd_sc_hd__a31o_1
Xhold1466 datamem.data_ram\[8\]\[17\] VGND VGND VPWR VPWR net2616 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1477 datamem.data_ram\[38\]\[11\] VGND VGND VPWR VPWR net2627 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1488 datamem.data_ram\[26\]\[12\] VGND VGND VPWR VPWR net2638 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_200_5284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_528 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_200_5295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1499 datamem.data_ram\[19\]\[26\] VGND VGND VPWR VPWR net2649 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__10241_ _10241_ VGND VGND VPWR VPWR clknet_0__10241_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_212_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23185__855 clknet_1_0__leaf__10112_ VGND VGND VPWR VPWR net981 sky130_fd_sc_hd__inv_2
X_29360_ clknet_leaf_261_clk _01095_ VGND VGND VPWR VPWR datamem.data_ram\[61\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_22804_ _09441_ _09943_ VGND VGND VPWR VPWR _09944_ sky130_fd_sc_hd__nor2_1
X_26572_ _11631_ VGND VGND VPWR VPWR _03230_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20996_ datamem.data_ram\[30\]\[15\] datamem.data_ram\[31\]\[15\] _06651_ VGND VGND
+ VPWR VPWR _08285_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28311_ _12458_ net4078 _12623_ VGND VGND VPWR VPWR _12629_ sky130_fd_sc_hd__mux2_1
X_25523_ _10055_ VGND VGND VPWR VPWR _11018_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_0__10172_ _10172_ VGND VGND VPWR VPWR clknet_0__10172_ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_0_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22735_ _09415_ _09876_ _09878_ _09488_ VGND VGND VPWR VPWR _09879_ sky130_fd_sc_hd__o211a_1
X_29291_ _09329_ net1935 _13159_ VGND VGND VPWR VPWR _13167_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_213_5601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_192_5096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_213_5612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28242_ _12590_ VGND VGND VPWR VPWR _03941_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_211_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25454_ _10070_ _10981_ _10982_ net1350 VGND VGND VPWR VPWR _02761_ sky130_fd_sc_hd__a22o_1
XFILLER_0_192_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22666_ _09705_ _09805_ _09809_ _09813_ VGND VGND VPWR VPWR _09814_ sky130_fd_sc_hd__and4_1
XFILLER_0_30_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23457__106 clknet_1_0__leaf__10157_ VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__inv_2
XFILLER_0_211_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24405_ _09285_ net4256 _10376_ VGND VGND VPWR VPWR _10382_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21617_ _08865_ _08866_ _08540_ VGND VGND VPWR VPWR _08867_ sky130_fd_sc_hd__mux2_1
X_28173_ _12553_ VGND VGND VPWR VPWR _03909_ sky130_fd_sc_hd__clkbuf_1
X_25385_ _10938_ net1382 _10934_ _10944_ VGND VGND VPWR VPWR _02730_ sky130_fd_sc_hd__a31o_1
XFILLER_0_146_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_109_Right_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22597_ rvcpu.dp.rf.reg_file_arr\[28\]\[15\] rvcpu.dp.rf.reg_file_arr\[30\]\[15\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[15\] rvcpu.dp.rf.reg_file_arr\[31\]\[15\] _09400_
+ _09484_ VGND VGND VPWR VPWR _09748_ sky130_fd_sc_hd__mux4_1
XFILLER_0_152_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27124_ _11835_ _11953_ VGND VGND VPWR VPWR _11961_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24336_ _10344_ VGND VGND VPWR VPWR _02281_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_11_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21548_ rvcpu.dp.rf.reg_file_arr\[20\]\[9\] rvcpu.dp.rf.reg_file_arr\[21\]\[9\] rvcpu.dp.rf.reg_file_arr\[22\]\[9\]
+ rvcpu.dp.rf.reg_file_arr\[23\]\[9\] _08799_ _08800_ VGND VGND VPWR VPWR _08801_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_16_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27055_ _06587_ VGND VGND VPWR VPWR _11918_ sky130_fd_sc_hd__buf_2
XFILLER_0_132_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24267_ _09330_ net3982 _10298_ VGND VGND VPWR VPWR _10306_ sky130_fd_sc_hd__mux2_1
X_21479_ rvcpu.dp.rf.reg_file_arr\[4\]\[5\] rvcpu.dp.rf.reg_file_arr\[5\]\[5\] rvcpu.dp.rf.reg_file_arr\[6\]\[5\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[5\] _08567_ _08570_ VGND VGND VPWR VPWR _08736_ sky130_fd_sc_hd__mux4_1
XFILLER_0_161_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26006_ net17 _11317_ VGND VGND VPWR VPWR _11328_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24198_ _06997_ VGND VGND VPWR VPWR _10268_ sky130_fd_sc_hd__buf_8
XFILLER_0_222_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_4420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_164_4431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_4442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27957_ _12430_ net3817 _12431_ VGND VGND VPWR VPWR _12432_ sky130_fd_sc_hd__mux2_1
X_15971_ net2167 _13213_ _14322_ VGND VGND VPWR VPWR _14323_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_160_4328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_160_4339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17710_ _13213_ net3104 _05129_ VGND VGND VPWR VPWR _05130_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26908_ _11829_ _11823_ VGND VGND VPWR VPWR _11830_ sky130_fd_sc_hd__and2_1
X_14922_ _13332_ _13462_ VGND VGND VPWR VPWR _13471_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18690_ _05866_ _05697_ _05845_ _06043_ VGND VGND VPWR VPWR _06044_ sky130_fd_sc_hd__a31o_1
X_27888_ _11965_ _12394_ VGND VGND VPWR VPWR _12395_ sky130_fd_sc_hd__and2_1
XFILLER_0_216_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold60 rvcpu.dp.plde.PCPlus4E\[18\] VGND VGND VPWR VPWR net1210 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 rvcpu.dp.plem.lAuiPCM\[30\] VGND VGND VPWR VPWR net1221 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 rvcpu.dp.plde.PCPlus4E\[14\] VGND VGND VPWR VPWR net1232 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2690 datamem.data_ram\[4\]\[12\] VGND VGND VPWR VPWR net3840 sky130_fd_sc_hd__dlygate4sd3_1
X_17641_ _05081_ VGND VGND VPWR VPWR _05093_ sky130_fd_sc_hd__buf_4
X_26839_ _11781_ net1707 _11785_ _11787_ VGND VGND VPWR VPWR _03341_ sky130_fd_sc_hd__a31o_1
X_14853_ _13367_ _13405_ VGND VGND VPWR VPWR _13406_ sky130_fd_sc_hd__or2_1
X_29627_ net981 _01362_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[25\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_216_1123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold93 rvcpu.dp.plem.PCPlus4M\[13\] VGND VGND VPWR VPWR net1243 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_216_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29558_ net912 _01293_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[27\]\[25\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_63_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17572_ _05056_ VGND VGND VPWR VPWR _01250_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_199_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14784_ _13335_ _13336_ VGND VGND VPWR VPWR _13337_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_63_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19311_ rvcpu.dp.plem.ALUResultM\[4\] _06606_ VGND VGND VPWR VPWR _06607_ sky130_fd_sc_hd__nor2_4
X_16523_ _04499_ VGND VGND VPWR VPWR _01782_ sky130_fd_sc_hd__clkbuf_1
X_28509_ _09278_ VGND VGND VPWR VPWR _12741_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_158_4279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29489_ net851 _01224_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[2\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31520_ clknet_leaf_49_clk net1232 VGND VGND VPWR VPWR rvcpu.dp.plem.PCPlus4M\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_19242_ _06546_ VGND VGND VPWR VPWR rvcpu.dp.lAuiPCE\[28\] sky130_fd_sc_hd__clkbuf_1
X_16454_ net2318 _14484_ _14560_ VGND VGND VPWR VPWR _04462_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15405_ _13449_ _13718_ VGND VGND VPWR VPWR _13937_ sky130_fd_sc_hd__or2_1
XFILLER_0_186_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19173_ rvcpu.dp.plde.ImmExtE\[20\] rvcpu.dp.plde.PCE\[20\] VGND VGND VPWR VPWR _06486_
+ sky130_fd_sc_hd__or2_1
X_31451_ clknet_leaf_2_clk rvcpu.dp.SrcBFW_Mux.y\[9\] VGND VGND VPWR VPWR rvcpu.dp.plem.WriteDataM\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_213_82 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16385_ _14557_ VGND VGND VPWR VPWR _01846_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_22_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18124_ _13222_ rvcpu.dp.plde.RD2E\[18\] _05194_ VGND VGND VPWR VPWR _05491_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_22_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30402_ net740 _02137_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[31\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_15336_ _13509_ _13565_ VGND VGND VPWR VPWR _13872_ sky130_fd_sc_hd__or2_1
XFILLER_0_170_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31382_ clknet_leaf_18_clk _03085_ VGND VGND VPWR VPWR rvcpu.dp.plde.ImmExtE\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_117_3297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18055_ _05423_ VGND VGND VPWR VPWR rvcpu.dp.SrcBFW_Mux.y\[8\] sky130_fd_sc_hd__buf_1
X_30333_ net679 _02068_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[4\]\[16\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_93_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15267_ _13805_ _13758_ _13533_ VGND VGND VPWR VPWR _13806_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_93_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2 _01054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__10161_ clknet_0__10161_ VGND VGND VPWR VPWR clknet_1_0__leaf__10161_
+ sky130_fd_sc_hd__clkbuf_16
X_17006_ _04464_ _04755_ VGND VGND VPWR VPWR _04756_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_188_4998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30264_ net618 _01999_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[6\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_15198_ _13639_ _13657_ _13496_ VGND VGND VPWR VPWR _13740_ sky130_fd_sc_hd__o21a_1
XFILLER_0_10_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32003_ clknet_leaf_133_clk _03425_ VGND VGND VPWR VPWR datamem.data_ram\[52\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_30195_ net549 _01930_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[8\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_52_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18957_ _05240_ _06292_ _06293_ VGND VGND VPWR VPWR _06294_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_52_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17908_ _05275_ _05280_ VGND VGND VPWR VPWR _05281_ sky130_fd_sc_hd__or2_1
XFILLER_0_158_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18888_ _05463_ _05469_ _05475_ _05484_ _05666_ _05671_ VGND VGND VPWR VPWR _06230_
+ sky130_fd_sc_hd__mux4_1
X_32905_ clknet_leaf_260_clk _04327_ VGND VGND VPWR VPWR datamem.data_ram\[7\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_17839_ _05220_ VGND VGND VPWR VPWR rvcpu.dp.SrcBFW_Mux.y\[19\] sky130_fd_sc_hd__clkbuf_2
X_20850_ _07823_ datamem.data_ram\[6\]\[14\] datamem.data_ram\[7\]\[14\] _07849_ _07860_
+ VGND VGND VPWR VPWR _08140_ sky130_fd_sc_hd__a221o_1
XFILLER_0_222_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23249__896 clknet_1_1__leaf__10127_ VGND VGND VPWR VPWR net1022 sky130_fd_sc_hd__inv_2
X_32836_ clknet_leaf_254_clk _04258_ VGND VGND VPWR VPWR datamem.data_ram\[12\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19509_ _06685_ VGND VGND VPWR VPWR _06805_ sky130_fd_sc_hd__clkbuf_8
X_20781_ datamem.data_ram\[6\]\[30\] datamem.data_ram\[7\]\[30\] _07836_ VGND VGND
+ VPWR VPWR _08071_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32767_ clknet_leaf_282_clk _04189_ VGND VGND VPWR VPWR datamem.data_ram\[15\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22520_ _09636_ _09674_ VGND VGND VPWR VPWR _09675_ sky130_fd_sc_hd__nor2_1
XFILLER_0_147_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31718_ net167 _03176_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[9\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_32698_ clknet_leaf_266_clk _04120_ VGND VGND VPWR VPWR datamem.data_ram\[17\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31649_ clknet_leaf_25_clk net1192 VGND VGND VPWR VPWR rvcpu.dp.plmw.lAuiPCW\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_22451_ rvcpu.dp.rf.reg_file_arr\[12\]\[7\] rvcpu.dp.rf.reg_file_arr\[13\]\[7\] rvcpu.dp.rf.reg_file_arr\[14\]\[7\]
+ rvcpu.dp.rf.reg_file_arr\[15\]\[7\] _09552_ _09382_ VGND VGND VPWR VPWR _09610_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_146_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21402_ _08511_ _08661_ VGND VGND VPWR VPWR _08662_ sky130_fd_sc_hd__nor2_1
X_22382_ rvcpu.dp.rf.reg_file_arr\[20\]\[4\] rvcpu.dp.rf.reg_file_arr\[21\]\[4\] rvcpu.dp.rf.reg_file_arr\[22\]\[4\]
+ rvcpu.dp.rf.reg_file_arr\[23\]\[4\] _09512_ _09408_ VGND VGND VPWR VPWR _09544_
+ sky130_fd_sc_hd__mux4_1
X_25170_ _09317_ VGND VGND VPWR VPWR _10820_ sky130_fd_sc_hd__buf_2
XFILLER_0_143_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23985__520 clknet_1_0__leaf__10239_ VGND VGND VPWR VPWR net646 sky130_fd_sc_hd__inv_2
X_21333_ rvcpu.dp.plfd.InstrD\[21\] VGND VGND VPWR VPWR _08595_ sky130_fd_sc_hd__buf_4
XFILLER_0_114_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_206_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold530 _02914_ VGND VGND VPWR VPWR net1680 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21264_ rvcpu.dp.plfd.InstrD\[16\] VGND VGND VPWR VPWR _08526_ sky130_fd_sc_hd__buf_4
XFILLER_0_13_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold541 datamem.data_ram\[62\]\[4\] VGND VGND VPWR VPWR net1691 sky130_fd_sc_hd__dlygate4sd3_1
Xhold552 datamem.data_ram\[1\]\[2\] VGND VGND VPWR VPWR net1702 sky130_fd_sc_hd__dlygate4sd3_1
X_20215_ datamem.data_ram\[30\]\[3\] _07127_ _06977_ datamem.data_ram\[28\]\[3\] VGND
+ VGND VPWR VPWR _07508_ sky130_fd_sc_hd__a22o_1
Xhold563 datamem.data_ram\[39\]\[2\] VGND VGND VPWR VPWR net1713 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold574 datamem.data_ram\[15\]\[4\] VGND VGND VPWR VPWR net1724 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28860_ _12690_ net2964 _12932_ VGND VGND VPWR VPWR _12934_ sky130_fd_sc_hd__mux2_1
X_21195_ _08471_ _08478_ VGND VGND VPWR VPWR _08479_ sky130_fd_sc_hd__or2_1
Xhold585 datamem.data_ram\[27\]\[7\] VGND VGND VPWR VPWR net1735 sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 datamem.data_ram\[24\]\[1\] VGND VGND VPWR VPWR net1746 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_8_Left_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27811_ _12348_ VGND VGND VPWR VPWR _03752_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_204_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20146_ datamem.data_ram\[59\]\[27\] _06729_ _06668_ datamem.data_ram\[63\]\[27\]
+ VGND VGND VPWR VPWR _07439_ sky130_fd_sc_hd__o22a_1
XFILLER_0_218_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28791_ _12897_ VGND VGND VPWR VPWR _04183_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_202_5335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_202_5346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27742_ _12310_ VGND VGND VPWR VPWR _03721_ sky130_fd_sc_hd__clkbuf_1
X_24954_ _10113_ _10640_ _10611_ VGND VGND VPWR VPWR _10696_ sky130_fd_sc_hd__a21oi_4
X_20077_ datamem.data_ram\[42\]\[10\] _06803_ _06726_ datamem.data_ram\[47\]\[10\]
+ VGND VGND VPWR VPWR _07371_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_198_5250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1230 rvcpu.dp.rf.reg_file_arr\[19\]\[3\] VGND VGND VPWR VPWR net2380 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1241 rvcpu.dp.rf.reg_file_arr\[9\]\[23\] VGND VGND VPWR VPWR net2391 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1252 rvcpu.dp.rf.reg_file_arr\[3\]\[15\] VGND VGND VPWR VPWR net2402 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27673_ _12273_ VGND VGND VPWR VPWR _03689_ sky130_fd_sc_hd__clkbuf_1
X_24885_ _09226_ _10630_ _10611_ VGND VGND VPWR VPWR _10659_ sky130_fd_sc_hd__a21oi_4
Xhold1263 rvcpu.dp.rf.reg_file_arr\[3\]\[22\] VGND VGND VPWR VPWR net2413 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1274 rvcpu.dp.rf.reg_file_arr\[2\]\[23\] VGND VGND VPWR VPWR net2424 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_194_5147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29412_ clknet_leaf_290_clk _01147_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD2E\[23\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1285 rvcpu.dp.rf.reg_file_arr\[25\]\[16\] VGND VGND VPWR VPWR net2435 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_194_5158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26624_ _10048_ _11659_ _11660_ net1316 VGND VGND VPWR VPWR _03253_ sky130_fd_sc_hd__a22o_1
XANTENNA_403 _06632_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1296 datamem.data_ram\[37\]\[29\] VGND VGND VPWR VPWR net2446 sky130_fd_sc_hd__dlygate4sd3_1
X_23836_ _10214_ VGND VGND VPWR VPWR _01911_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_170_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_414 _06667_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_170_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_425 _06783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_436 _06922_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_0__10224_ _10224_ VGND VGND VPWR VPWR clknet_0__10224_ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_1__f__10124_ clknet_0__10124_ VGND VGND VPWR VPWR clknet_1_1__leaf__10124_
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_447 _07845_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29343_ clknet_leaf_198_clk _01078_ VGND VGND VPWR VPWR datamem.data_ram\[61\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_458 _08634_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26555_ _11622_ VGND VGND VPWR VPWR _03222_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20979_ _07844_ _08264_ _08267_ _06676_ VGND VGND VPWR VPWR _08268_ sky130_fd_sc_hd__a211o_1
XANTENNA_469 _08873_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25506_ _07028_ _10918_ _10897_ VGND VGND VPWR VPWR _11008_ sky130_fd_sc_hd__or3_1
Xclkbuf_0__10155_ _10155_ VGND VGND VPWR VPWR clknet_0__10155_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_71_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29274_ _09290_ net2477 _13150_ VGND VGND VPWR VPWR _13158_ sky130_fd_sc_hd__mux2_1
X_22718_ rvcpu.dp.rf.reg_file_arr\[4\]\[21\] rvcpu.dp.rf.reg_file_arr\[5\]\[21\] rvcpu.dp.rf.reg_file_arr\[6\]\[21\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[21\] _09464_ _09467_ VGND VGND VPWR VPWR _09863_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_211_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28225_ _12581_ VGND VGND VPWR VPWR _03933_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_211_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_153_4165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25437_ _10760_ net3663 _10970_ VGND VGND VPWR VPWR _10975_ sky130_fd_sc_hd__mux2_1
Xclkbuf_0__10086_ _10086_ VGND VGND VPWR VPWR clknet_0__10086_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_125_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22649_ _09797_ VGND VGND VPWR VPWR _01141_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_193_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_4176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22981__688 clknet_1_0__leaf__10083_ VGND VGND VPWR VPWR net814 sky130_fd_sc_hd__inv_2
X_16170_ _14431_ VGND VGND VPWR VPWR _01943_ sky130_fd_sc_hd__clkbuf_1
X_28156_ _12544_ VGND VGND VPWR VPWR _03901_ sky130_fd_sc_hd__clkbuf_1
X_25368_ _10933_ VGND VGND VPWR VPWR _10934_ sky130_fd_sc_hd__buf_2
XFILLER_0_63_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15121_ _13665_ _13294_ VGND VGND VPWR VPWR _13666_ sky130_fd_sc_hd__nand2_1
X_27107_ _11938_ net1774 _11940_ _11950_ VGND VGND VPWR VPWR _03446_ sky130_fd_sc_hd__a31o_1
X_24319_ _09326_ net4391 _10328_ VGND VGND VPWR VPWR _10335_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28087_ _12443_ net3768 _12501_ VGND VGND VPWR VPWR _12508_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25299_ _10892_ VGND VGND VPWR VPWR _02696_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27038_ _11837_ _11899_ VGND VGND VPWR VPWR _11908_ sky130_fd_sc_hd__and2_1
X_15052_ _13358_ VGND VGND VPWR VPWR _13599_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_181_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_3172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput4 net4 VGND VGND VPWR VPWR Instr[11] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_112_3183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23354__991 clknet_1_0__leaf__10137_ VGND VGND VPWR VPWR net1117 sky130_fd_sc_hd__inv_2
X_19860_ datamem.data_ram\[0\]\[1\] _06990_ _06966_ datamem.data_ram\[3\]\[1\] VGND
+ VGND VPWR VPWR _07155_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_183_4884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18811_ _06094_ _06157_ _05706_ VGND VGND VPWR VPWR _06158_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_183_4895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19791_ datamem.data_ram\[54\]\[9\] _07085_ _06633_ datamem.data_ram\[51\]\[9\] VGND
+ VGND VPWR VPWR _07086_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_125_3500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28989_ _12696_ net2140 _12999_ VGND VGND VPWR VPWR _13004_ sky130_fd_sc_hd__mux2_1
X_18742_ _06025_ VGND VGND VPWR VPWR _06093_ sky130_fd_sc_hd__inv_2
X_15954_ net3883 _13187_ _14311_ VGND VGND VPWR VPWR _14314_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14905_ _13315_ _13455_ VGND VGND VPWR VPWR _13456_ sky130_fd_sc_hd__nor2_1
X_18673_ _05805_ _06024_ _06027_ _05702_ VGND VGND VPWR VPWR _06028_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_121_3408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30951_ clknet_leaf_263_clk _02686_ VGND VGND VPWR VPWR datamem.data_ram\[3\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_222_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_196_clk clknet_5_29__leaf_clk VGND VGND VPWR VPWR clknet_leaf_196_clk
+ sky130_fd_sc_hd__clkbuf_8
X_15885_ _14277_ VGND VGND VPWR VPWR _02082_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_208_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_86_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14836_ _13388_ VGND VGND VPWR VPWR _13389_ sky130_fd_sc_hd__buf_4
XFILLER_0_188_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17624_ _05084_ VGND VGND VPWR VPWR _01226_ sky130_fd_sc_hd__clkbuf_1
X_30882_ clknet_leaf_180_clk _02617_ VGND VGND VPWR VPWR datamem.data_ram\[42\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_187_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17555_ _13184_ net4315 _05046_ VGND VGND VPWR VPWR _05048_ sky130_fd_sc_hd__mux2_1
X_32621_ clknet_leaf_287_clk _04043_ VGND VGND VPWR VPWR datamem.data_ram\[20\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_14767_ _13305_ VGND VGND VPWR VPWR _13320_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_15_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23854__417 clknet_1_0__leaf__10219_ VGND VGND VPWR VPWR net543 sky130_fd_sc_hd__inv_2
XFILLER_0_128_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16506_ net2527 _14466_ _04489_ VGND VGND VPWR VPWR _04491_ sky130_fd_sc_hd__mux2_1
X_32552_ clknet_leaf_272_clk _03974_ VGND VGND VPWR VPWR datamem.data_ram\[23\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17486_ _05011_ VGND VGND VPWR VPWR _01299_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14698_ _13258_ VGND VGND VPWR VPWR _03179_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_15_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31503_ clknet_leaf_24_clk rvcpu.dp.lAuiPCE\[29\] VGND VGND VPWR VPWR rvcpu.dp.plem.lAuiPCM\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_119_3348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19225_ _06531_ rvcpu.dp.plde.ImmExtE\[26\] _06493_ VGND VGND VPWR VPWR _06532_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_119_3359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16437_ _04453_ VGND VGND VPWR VPWR _01822_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32483_ clknet_leaf_240_clk _03905_ VGND VGND VPWR VPWR datamem.data_ram\[25\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_211_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31434_ clknet_leaf_103_clk _03137_ VGND VGND VPWR VPWR datamem.data_ram\[14\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_19156_ _06464_ _06470_ VGND VGND VPWR VPWR _06471_ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16368_ net1872 _14466_ _14547_ VGND VGND VPWR VPWR _14549_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18107_ rvcpu.dp.plde.RD1E\[20\] _05292_ _05474_ VGND VGND VPWR VPWR _05475_ sky130_fd_sc_hd__o21a_2
XFILLER_0_5_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15319_ _13359_ _13410_ _13465_ _13855_ rvcpu.dp.pcreg.q\[9\] VGND VGND VPWR VPWR
+ _13856_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_41_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19087_ _06408_ _06410_ VGND VGND VPWR VPWR _06411_ sky130_fd_sc_hd__xnor2_2
X_31365_ clknet_leaf_24_clk _03068_ VGND VGND VPWR VPWR rvcpu.dp.plde.ImmExtE\[14\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_152_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_120_clk clknet_5_27__leaf_clk VGND VGND VPWR VPWR clknet_leaf_120_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_112_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16299_ _14512_ VGND VGND VPWR VPWR _01887_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18038_ rvcpu.dp.plde.RD1E\[11\] _05267_ _05271_ _13243_ _05407_ VGND VGND VPWR VPWR
+ _05408_ sky130_fd_sc_hd__a221oi_4
X_30316_ net662 _02051_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[5\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31296_ clknet_leaf_38_clk _02999_ VGND VGND VPWR VPWR rvcpu.dp.plde.PCPlus4E\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30247_ net601 _01982_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[6\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20000_ datamem.data_ram\[29\]\[2\] _06919_ _06953_ datamem.data_ram\[28\]\[2\] VGND
+ VGND VPWR VPWR _07294_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_226_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24178__19 clknet_1_0__leaf__10265_ VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__inv_2
X_30178_ clknet_leaf_205_clk _01913_ VGND VGND VPWR VPWR datamem.data_ram\[58\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_19989_ datamem.data_ram\[2\]\[2\] _06931_ _06920_ datamem.data_ram\[5\]\[2\] VGND
+ VGND VPWR VPWR _07283_ sky130_fd_sc_hd__a22o_1
XFILLER_0_226_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_179_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21951_ rvcpu.dp.rf.reg_file_arr\[28\]\[30\] rvcpu.dp.rf.reg_file_arr\[30\]\[30\]
+ rvcpu.dp.rf.reg_file_arr\[29\]\[30\] rvcpu.dp.rf.reg_file_arr\[31\]\[30\] _08533_
+ _08636_ VGND VGND VPWR VPWR _09183_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_2_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_187_clk clknet_5_22__leaf_clk VGND VGND VPWR VPWR clknet_leaf_187_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_206_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20902_ _07823_ datamem.data_ram\[11\]\[22\] _07835_ datamem.data_ram\[10\]\[22\]
+ _07845_ VGND VGND VPWR VPWR _08192_ sky130_fd_sc_hd__o221a_1
X_24670_ _10076_ _10532_ VGND VGND VPWR VPWR _10541_ sky130_fd_sc_hd__and2_1
X_21882_ rvcpu.dp.rf.reg_file_arr\[12\]\[26\] rvcpu.dp.rf.reg_file_arr\[13\]\[26\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[26\] rvcpu.dp.rf.reg_file_arr\[15\]\[26\] _08578_
+ _08684_ VGND VGND VPWR VPWR _09118_ sky130_fd_sc_hd__mux4_1
XFILLER_0_96_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20833_ _08082_ _08095_ _08122_ VGND VGND VPWR VPWR _08123_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_49_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32819_ clknet_leaf_212_clk _04241_ VGND VGND VPWR VPWR datamem.data_ram\[12\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_204_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26340_ _11501_ net1811 _11496_ _11505_ VGND VGND VPWR VPWR _03124_ sky130_fd_sc_hd__a31o_1
XFILLER_0_159_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_194_Right_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20764_ datamem.data_ram\[50\]\[6\] _07000_ _07133_ datamem.data_ram\[49\]\[6\] VGND
+ VGND VPWR VPWR _08054_ sky130_fd_sc_hd__a22o_1
X_26493__46 clknet_1_1__leaf__11601_ VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__inv_2
XFILLER_0_193_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22503_ rvcpu.dp.rf.reg_file_arr\[24\]\[10\] rvcpu.dp.rf.reg_file_arr\[25\]\[10\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[10\] rvcpu.dp.rf.reg_file_arr\[27\]\[10\] _09385_
+ _09637_ VGND VGND VPWR VPWR _09659_ sky130_fd_sc_hd__mux4_1
XFILLER_0_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24052__580 clknet_1_0__leaf__10246_ VGND VGND VPWR VPWR net706 sky130_fd_sc_hd__inv_2
X_26271_ net1807 _11467_ VGND VGND VPWR VPWR _11468_ sky130_fd_sc_hd__and2_1
XFILLER_0_162_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20695_ _07976_ _07980_ _07071_ _07985_ VGND VGND VPWR VPWR _07986_ sky130_fd_sc_hd__o211a_1
X_28010_ _12361_ net3665 net97 VGND VGND VPWR VPWR _12467_ sky130_fd_sc_hd__mux2_1
XFILLER_0_190_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25222_ _10850_ VGND VGND VPWR VPWR _02661_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22434_ _09389_ _09584_ _09589_ _09593_ VGND VGND VPWR VPWR _09594_ sky130_fd_sc_hd__and4_1
XFILLER_0_91_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25153_ _10764_ net2604 _10802_ VGND VGND VPWR VPWR _10809_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_111_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_111_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_66_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22365_ _09421_ VGND VGND VPWR VPWR _09528_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_33_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21316_ _08517_ VGND VGND VPWR VPWR _08578_ sky130_fd_sc_hd__clkbuf_8
X_29961_ net331 _01696_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[15\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25084_ _10773_ VGND VGND VPWR VPWR _02600_ sky130_fd_sc_hd__clkbuf_1
X_22296_ _09452_ VGND VGND VPWR VPWR _09461_ sky130_fd_sc_hd__buf_4
XFILLER_0_14_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21247_ rvcpu.dp.plfd.InstrD\[19\] VGND VGND VPWR VPWR _08509_ sky130_fd_sc_hd__inv_2
X_28912_ _12961_ VGND VGND VPWR VPWR _04240_ sky130_fd_sc_hd__clkbuf_1
X_24035_ clknet_1_1__leaf__10244_ VGND VGND VPWR VPWR _10245_ sky130_fd_sc_hd__buf_1
Xhold360 datamem.data_ram\[31\]\[2\] VGND VGND VPWR VPWR net1510 sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 datamem.data_ram\[54\]\[2\] VGND VGND VPWR VPWR net1521 sky130_fd_sc_hd__dlygate4sd3_1
X_29892_ net270 _01627_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[17\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold382 datamem.data_ram\[63\]\[2\] VGND VGND VPWR VPWR net1532 sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 datamem.data_ram\[19\]\[1\] VGND VGND VPWR VPWR net1543 sky130_fd_sc_hd__dlygate4sd3_1
X_21178_ _06580_ _08465_ VGND VGND VPWR VPWR _08467_ sky130_fd_sc_hd__or2_1
X_28843_ _12737_ net2408 net69 VGND VGND VPWR VPWR _12925_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_225_5891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20129_ datamem.data_ram\[10\]\[27\] _06804_ _07037_ datamem.data_ram\[13\]\[27\]
+ _07421_ VGND VGND VPWR VPWR _07422_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_196_5209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28774_ _12888_ VGND VGND VPWR VPWR _04175_ sky130_fd_sc_hd__clkbuf_1
X_25986_ _11157_ VGND VGND VPWR VPWR _11317_ sky130_fd_sc_hd__clkbuf_2
X_24094__603 clknet_1_0__leaf__10248_ VGND VGND VPWR VPWR net729 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_221_5788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_221_5799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27725_ _12301_ VGND VGND VPWR VPWR _03713_ sky130_fd_sc_hd__clkbuf_1
X_24937_ _10113_ _10630_ _10611_ VGND VGND VPWR VPWR _10687_ sky130_fd_sc_hd__a21oi_4
Xclkbuf_leaf_178_clk clknet_5_19__leaf_clk VGND VGND VPWR VPWR clknet_leaf_178_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold1060 rvcpu.dp.rf.reg_file_arr\[10\]\[8\] VGND VGND VPWR VPWR net2210 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1071 rvcpu.dp.rf.reg_file_arr\[23\]\[26\] VGND VGND VPWR VPWR net2221 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27656_ _12264_ VGND VGND VPWR VPWR _03681_ sky130_fd_sc_hd__clkbuf_1
Xhold1082 rvcpu.dp.rf.reg_file_arr\[9\]\[0\] VGND VGND VPWR VPWR net2232 sky130_fd_sc_hd__dlygate4sd3_1
X_15670_ _14150_ VGND VGND VPWR VPWR _02178_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_200 _09476_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24868_ _09226_ _10601_ _10611_ VGND VGND VPWR VPWR _10650_ sky130_fd_sc_hd__a21oi_1
Xhold1093 rvcpu.dp.rf.reg_file_arr\[18\]\[18\] VGND VGND VPWR VPWR net2243 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_211 _09635_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_213_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_222 _09953_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_212_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14621_ rvcpu.dp.plmw.ALUResultW\[25\] rvcpu.dp.plmw.ReadDataW\[25\] rvcpu.dp.plmw.PCPlus4W\[25\]
+ rvcpu.dp.plmw.lAuiPCW\[25\] _13192_ _13193_ VGND VGND VPWR VPWR _13200_ sky130_fd_sc_hd__mux4_2
X_26607_ _11651_ VGND VGND VPWR VPWR _03245_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_233 _10142_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_4205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_244 _11687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_213_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_155_4216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27587_ _12227_ VGND VGND VPWR VPWR _03649_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_213_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_155_4227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24799_ _10439_ net3258 _10612_ VGND VGND VPWR VPWR _10613_ sky130_fd_sc_hd__mux2_1
XANTENNA_255 _13200_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_266 _13225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_0__10207_ _10207_ VGND VGND VPWR VPWR clknet_0__10207_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_184_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29326_ clknet_leaf_141_clk _01061_ VGND VGND VPWR VPWR datamem.data_ram\[62\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_17340_ _04933_ VGND VGND VPWR VPWR _01375_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_277 _13244_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26538_ _11083_ _11610_ VGND VGND VPWR VPWR _11613_ sky130_fd_sc_hd__and2_1
Xclkbuf_1_1__f__10107_ clknet_0__10107_ VGND VGND VPWR VPWR clknet_1_1__leaf__10107_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_23_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_288 _13304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_299 _13891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_161_Right_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_484 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0__10138_ _10138_ VGND VGND VPWR VPWR clknet_0__10138_ sky130_fd_sc_hd__clkbuf_16
X_29257_ _09259_ net3614 _13141_ VGND VGND VPWR VPWR _13149_ sky130_fd_sc_hd__mux2_1
X_17271_ _04896_ VGND VGND VPWR VPWR _01407_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_181_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26469_ _11535_ rvcpu.ALUResultE\[28\] _11288_ VGND VGND VPWR VPWR _11591_ sky130_fd_sc_hd__a21o_1
XFILLER_0_138_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_181_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19010_ _05661_ _06115_ _06341_ _06343_ VGND VGND VPWR VPWR _06344_ sky130_fd_sc_hd__a211o_1
XFILLER_0_138_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16222_ net2247 _14466_ _14464_ VGND VGND VPWR VPWR _14467_ sky130_fd_sc_hd__mux2_1
X_28208_ _12462_ net3074 _12564_ VGND VGND VPWR VPWR _12572_ sky130_fd_sc_hd__mux2_1
X_29188_ _13111_ VGND VGND VPWR VPWR _04366_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_114_3223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_3234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload208 clknet_leaf_202_clk VGND VGND VPWR VPWR clkload208/Y sky130_fd_sc_hd__clkinvlp_2
X_28139_ _12535_ VGND VGND VPWR VPWR _03893_ sky130_fd_sc_hd__clkbuf_1
Xclkload219 clknet_leaf_175_clk VGND VGND VPWR VPWR clkload219/Y sky130_fd_sc_hd__clkinvlp_4
X_16153_ _14419_ VGND VGND VPWR VPWR _01948_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_102_clk clknet_5_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_102_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_144_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15104_ _13297_ _13560_ VGND VGND VPWR VPWR _13649_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_185_4924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31150_ clknet_leaf_70_clk rvcpu.ALUResultE\[9\] VGND VGND VPWR VPWR rvcpu.dp.plem.ALUResultM\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_185_4935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16084_ net2379 _13278_ _14348_ VGND VGND VPWR VPWR _14383_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_185_4946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24029__560 clknet_1_0__leaf__10243_ VGND VGND VPWR VPWR net686 sky130_fd_sc_hd__inv_2
XFILLER_0_146_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30101_ net463 _01836_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[11\]\[24\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_75_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15035_ _13324_ _13489_ _13381_ VGND VGND VPWR VPWR _13582_ sky130_fd_sc_hd__o21ba_1
X_19912_ datamem.data_ram\[44\]\[17\] _06621_ _07206_ _07081_ VGND VGND VPWR VPWR
+ _07207_ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31081_ clknet_leaf_107_clk _02816_ VGND VGND VPWR VPWR datamem.data_ram\[20\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30032_ net394 _01767_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[13\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19843_ _06973_ VGND VGND VPWR VPWR _07138_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_88_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19774_ _06713_ _07047_ _07058_ _07068_ _06797_ VGND VGND VPWR VPWR _07069_ sky130_fd_sc_hd__a32o_1
XFILLER_0_223_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_3953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16986_ _04745_ VGND VGND VPWR VPWR _01549_ sky130_fd_sc_hd__clkbuf_1
X_18725_ _05658_ _06004_ VGND VGND VPWR VPWR _06077_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_169_clk clknet_5_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_169_clk
+ sky130_fd_sc_hd__clkbuf_8
X_15937_ _14304_ VGND VGND VPWR VPWR _02057_ sky130_fd_sc_hd__clkbuf_1
X_31983_ clknet_leaf_119_clk _03405_ VGND VGND VPWR VPWR datamem.data_ram\[37\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_56 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18656_ _05427_ _05726_ _05974_ _05425_ _06011_ VGND VGND VPWR VPWR _06012_ sky130_fd_sc_hd__a221o_1
X_30934_ clknet_leaf_280_clk _02669_ VGND VGND VPWR VPWR datamem.data_ram\[40\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_15868_ _14266_ VGND VGND VPWR VPWR _02088_ sky130_fd_sc_hd__clkbuf_1
Xwire38 _06472_ VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_1
XFILLER_0_153_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14819_ _13371_ _13300_ VGND VGND VPWR VPWR _13372_ sky130_fd_sc_hd__nor2_2
XFILLER_0_149_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17607_ _13263_ net3579 _05068_ VGND VGND VPWR VPWR _05075_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30865_ clknet_leaf_261_clk _02600_ VGND VGND VPWR VPWR datamem.data_ram\[43\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_18587_ _05790_ _05941_ _05942_ _05945_ VGND VGND VPWR VPWR _05946_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_47_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15799_ _14229_ VGND VGND VPWR VPWR _02128_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32604_ clknet_leaf_244_clk _04026_ VGND VGND VPWR VPWR datamem.data_ram\[20\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17538_ _05038_ VGND VGND VPWR VPWR _01274_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_175_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30796_ clknet_leaf_172_clk _02531_ VGND VGND VPWR VPWR datamem.data_ram\[46\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_43_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17469_ _14183_ net4030 _04996_ VGND VGND VPWR VPWR _05002_ sky130_fd_sc_hd__mux2_1
X_32535_ clknet_leaf_184_clk _03957_ VGND VGND VPWR VPWR datamem.data_ram\[23\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_229_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_190_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19208_ _06501_ _06510_ _06508_ _06507_ VGND VGND VPWR VPWR _06517_ sky130_fd_sc_hd__a31o_1
X_20480_ datamem.data_ram\[52\]\[20\] _06618_ _07770_ _07771_ VGND VGND VPWR VPWR
+ _07772_ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32466_ clknet_leaf_81_clk _03888_ VGND VGND VPWR VPWR datamem.data_ram\[26\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_229_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31417_ clknet_leaf_53_clk _03120_ VGND VGND VPWR VPWR datamem.data_ram\[15\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_19139_ rvcpu.dp.plde.ImmExtE\[16\] rvcpu.dp.plde.PCE\[16\] VGND VGND VPWR VPWR _06456_
+ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_89_Left_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32397_ clknet_leaf_78_clk _03819_ VGND VGND VPWR VPWR datamem.data_ram\[29\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_22150_ _09279_ net3782 net62 VGND VGND VPWR VPWR _09345_ sky130_fd_sc_hd__mux2_1
X_31348_ clknet_leaf_22_clk _03051_ VGND VGND VPWR VPWR rvcpu.dp.plde.luiE sky130_fd_sc_hd__dfxtp_2
XFILLER_0_89_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21101_ datamem.data_ram\[9\]\[7\] _06944_ _06642_ _08389_ VGND VGND VPWR VPWR _08390_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_112_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22081_ _09294_ VGND VGND VPWR VPWR _09295_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31279_ clknet_leaf_125_clk _02982_ VGND VGND VPWR VPWR datamem.data_ram\[24\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__10127_ clknet_0__10127_ VGND VGND VPWR VPWR clknet_1_0__leaf__10127_
+ sky130_fd_sc_hd__clkbuf_16
X_21032_ _08318_ _08319_ _08320_ _07820_ _07866_ VGND VGND VPWR VPWR _08321_ sky130_fd_sc_hd__a221o_1
XFILLER_0_196_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_5_28__f_clk clknet_2_3_0_clk VGND VGND VPWR VPWR clknet_5_28__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_196_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25840_ rvcpu.dp.plfd.PCPlus4D\[24\] _11223_ _11142_ VGND VGND VPWR VPWR _11224_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_226_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25771_ _11149_ _11168_ _11169_ VGND VGND VPWR VPWR _11170_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_98_Left_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27510_ _12186_ VGND VGND VPWR VPWR _03613_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24722_ _10480_ net3042 _10561_ VGND VGND VPWR VPWR _10569_ sky130_fd_sc_hd__mux2_1
X_28490_ _12727_ net1591 _12723_ _12729_ VGND VGND VPWR VPWR _04050_ sky130_fd_sc_hd__a31o_1
X_21934_ _08686_ _09166_ _08806_ VGND VGND VPWR VPWR _09167_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_215_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27441_ _12146_ VGND VGND VPWR VPWR _03584_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24653_ _10530_ VGND VGND VPWR VPWR _10531_ sky130_fd_sc_hd__buf_2
XFILLER_0_136_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21865_ rvcpu.dp.rf.reg_file_arr\[8\]\[25\] rvcpu.dp.rf.reg_file_arr\[10\]\[25\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[25\] rvcpu.dp.rf.reg_file_arr\[11\]\[25\] _08635_
+ _08637_ VGND VGND VPWR VPWR _09102_ sky130_fd_sc_hd__mux4_1
XFILLER_0_78_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_985 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20816_ datamem.data_ram\[58\]\[30\] _06940_ _07832_ _08105_ VGND VGND VPWR VPWR
+ _08106_ sky130_fd_sc_hd__o211a_1
X_27372_ _12104_ VGND VGND VPWR VPWR _03557_ sky130_fd_sc_hd__clkbuf_1
X_24584_ _10388_ net3763 _10491_ VGND VGND VPWR VPWR _10493_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21796_ _08842_ _09036_ VGND VGND VPWR VPWR _09037_ sky130_fd_sc_hd__or2_1
X_29111_ _09278_ net2581 _13067_ VGND VGND VPWR VPWR _13071_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26323_ _07791_ _10932_ _11494_ VGND VGND VPWR VPWR _11495_ sky130_fd_sc_hd__or3_1
X_20747_ _06604_ _08029_ _08036_ _07858_ VGND VGND VPWR VPWR _08037_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_150_4102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_189_5024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_189_5035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29042_ _13018_ net1682 _13030_ _13034_ VGND VGND VPWR VPWR _04297_ sky130_fd_sc_hd__a31o_1
XFILLER_0_68_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26254_ net116 _11457_ _11439_ net4295 VGND VGND VPWR VPWR _03084_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_174_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23466_ clknet_1_1__leaf__10152_ VGND VGND VPWR VPWR _10158_ sky130_fd_sc_hd__buf_1
X_20678_ datamem.data_ram\[43\]\[5\] _07137_ _07125_ datamem.data_ram\[47\]\[5\] _07968_
+ VGND VGND VPWR VPWR _07969_ sky130_fd_sc_hd__a221o_1
XFILLER_0_162_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25205_ _10841_ VGND VGND VPWR VPWR _02653_ sky130_fd_sc_hd__clkbuf_1
X_22417_ _08595_ VGND VGND VPWR VPWR _09577_ sky130_fd_sc_hd__buf_4
XFILLER_0_61_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26185_ _11429_ VGND VGND VPWR VPWR _03045_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23397_ _10149_ VGND VGND VPWR VPWR _01537_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25136_ _10478_ net2470 _10793_ VGND VGND VPWR VPWR _10800_ sky130_fd_sc_hd__mux2_1
X_22348_ rvcpu.dp.plfd.InstrD\[22\] VGND VGND VPWR VPWR _09511_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_227_5942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_227_5953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_148_4042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25067_ _10763_ VGND VGND VPWR VPWR _02593_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_148_4053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29944_ net314 _01679_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[15\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_22279_ rvcpu.dp.rf.reg_file_arr\[16\]\[1\] rvcpu.dp.rf.reg_file_arr\[17\]\[1\] rvcpu.dp.rf.reg_file_arr\[18\]\[1\]
+ rvcpu.dp.rf.reg_file_arr\[19\]\[1\] _09416_ _09443_ VGND VGND VPWR VPWR _09444_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_218_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_223_5839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_4810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold190 datamem.data_ram\[44\]\[5\] VGND VGND VPWR VPWR net1340 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_180_4821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29875_ net253 _01610_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[17\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_24102__610 clknet_1_1__leaf__10258_ VGND VGND VPWR VPWR net736 sky130_fd_sc_hd__inv_2
XFILLER_0_229_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23582__204 clknet_1_0__leaf__10176_ VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__inv_2
XFILLER_0_40_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_218_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28826_ _12754_ net2892 _12914_ VGND VGND VPWR VPWR _12916_ sky130_fd_sc_hd__mux2_1
X_16840_ net2412 _14459_ _04659_ VGND VGND VPWR VPWR _04668_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_6_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16771_ _04631_ VGND VGND VPWR VPWR _01658_ sky130_fd_sc_hd__clkbuf_1
X_25969_ net4349 _11302_ _11300_ _11307_ VGND VGND VPWR VPWR _02951_ sky130_fd_sc_hd__o211a_1
X_28757_ _12690_ net3723 _12877_ VGND VGND VPWR VPWR _12879_ sky130_fd_sc_hd__mux2_1
XFILLER_0_219_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23662__261 clknet_1_0__leaf__10191_ VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_107_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18510_ _05675_ _05871_ VGND VGND VPWR VPWR _05872_ sky130_fd_sc_hd__nor2_1
X_15722_ _14185_ net3238 _14173_ VGND VGND VPWR VPWR _14186_ sky130_fd_sc_hd__mux2_1
X_27708_ _12292_ VGND VGND VPWR VPWR _03705_ sky130_fd_sc_hd__clkbuf_1
X_19490_ datamem.data_ram\[16\]\[16\] _06779_ _06783_ datamem.data_ram\[17\]\[16\]
+ _06785_ VGND VGND VPWR VPWR _06786_ sky130_fd_sc_hd__o221a_1
X_24059__586 clknet_1_0__leaf__10247_ VGND VGND VPWR VPWR net712 sky130_fd_sc_hd__inv_2
X_28688_ _12842_ VGND VGND VPWR VPWR _04135_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_178_4761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_185_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_178_4772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18441_ _05686_ _05801_ _05803_ _05669_ _05675_ VGND VGND VPWR VPWR _05804_ sky130_fd_sc_hd__a221o_1
X_15653_ _13194_ VGND VGND VPWR VPWR _14139_ sky130_fd_sc_hd__buf_4
X_27639_ _12132_ net2466 _12251_ VGND VGND VPWR VPWR _12255_ sky130_fd_sc_hd__mux2_1
XFILLER_0_186_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14604_ _13186_ VGND VGND VPWR VPWR _13187_ sky130_fd_sc_hd__buf_4
XFILLER_0_201_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18372_ _05275_ _05721_ _05724_ _05736_ VGND VGND VPWR VPWR _05737_ sky130_fd_sc_hd__a31o_1
X_22987__694 clknet_1_1__leaf__10083_ VGND VGND VPWR VPWR net820 sky130_fd_sc_hd__inv_2
X_30650_ clknet_leaf_189_clk _02385_ VGND VGND VPWR VPWR datamem.data_ram\[51\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15584_ _14099_ VGND VGND VPWR VPWR _02213_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_174_4669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17323_ rvcpu.dp.rf.reg_file_arr\[24\]\[11\] _13243_ _04924_ VGND VGND VPWR VPWR
+ _04925_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29309_ clknet_leaf_0_clk _01044_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD1E\[16\] sky130_fd_sc_hd__dfxtp_1
X_30581_ clknet_leaf_178_clk _02316_ VGND VGND VPWR VPWR datamem.data_ram\[53\]\[8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_139_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17254_ _14172_ net4320 _04887_ VGND VGND VPWR VPWR _04888_ sky130_fd_sc_hd__mux2_1
X_32320_ clknet_leaf_185_clk _03742_ VGND VGND VPWR VPWR datamem.data_ram\[31\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_3790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16205_ _13231_ VGND VGND VPWR VPWR _14455_ sky130_fd_sc_hd__buf_4
XFILLER_0_226_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32251_ clknet_leaf_167_clk _03673_ VGND VGND VPWR VPWR datamem.data_ram\[34\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17185_ _04828_ VGND VGND VPWR VPWR _04851_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_77_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_3676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31202_ clknet_leaf_30_clk _02905_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCPlus4D\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_133_3687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16136_ net2086 _13254_ _14407_ VGND VGND VPWR VPWR _14411_ sky130_fd_sc_hd__mux2_1
X_32182_ clknet_leaf_89_clk _03604_ VGND VGND VPWR VPWR datamem.data_ram\[37\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_133_3698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31133_ clknet_leaf_222_clk _02868_ VGND VGND VPWR VPWR datamem.data_ram\[4\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16067_ _14374_ VGND VGND VPWR VPWR _01989_ sky130_fd_sc_hd__clkbuf_1
Xhold3209 datamem.data_ram\[54\]\[17\] VGND VGND VPWR VPWR net4359 sky130_fd_sc_hd__dlygate4sd3_1
X_15018_ _13387_ _13565_ _13542_ VGND VGND VPWR VPWR _13566_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_52_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31064_ clknet_leaf_257_clk _02799_ VGND VGND VPWR VPWR datamem.data_ram\[8\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2508 datamem.data_ram\[5\]\[8\] VGND VGND VPWR VPWR net3658 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_36_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2519 datamem.data_ram\[41\]\[26\] VGND VGND VPWR VPWR net3669 sky130_fd_sc_hd__dlygate4sd3_1
X_30015_ net377 _01750_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[13\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_19826_ _05391_ _06586_ _07070_ _07119_ _07120_ VGND VGND VPWR VPWR _07121_ sky130_fd_sc_hd__o32a_1
Xhold1807 datamem.data_ram\[47\]\[22\] VGND VGND VPWR VPWR net2957 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1818 datamem.data_ram\[13\]\[17\] VGND VGND VPWR VPWR net2968 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1829 rvcpu.dp.rf.reg_file_arr\[14\]\[3\] VGND VGND VPWR VPWR net2979 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19757_ datamem.data_ram\[58\]\[25\] _07023_ _07048_ _07051_ VGND VGND VPWR VPWR
+ _07052_ sky130_fd_sc_hd__o211a_1
XFILLER_0_223_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16969_ _04736_ VGND VGND VPWR VPWR _01557_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_190_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18708_ _05775_ _05893_ VGND VGND VPWR VPWR _06061_ sky130_fd_sc_hd__nand2_1
X_31966_ clknet_leaf_120_clk _03388_ VGND VGND VPWR VPWR datamem.data_ram\[28\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_19688_ _06968_ _06975_ _06983_ _06716_ VGND VGND VPWR VPWR _06984_ sky130_fd_sc_hd__o211a_1
XFILLER_0_195_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18639_ _05980_ _05983_ _05992_ _05995_ VGND VGND VPWR VPWR _05996_ sky130_fd_sc_hd__or4b_1
X_30917_ clknet_leaf_221_clk _02652_ VGND VGND VPWR VPWR datamem.data_ram\[40\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31897_ _04437_ net120 VGND VGND VPWR VPWR datamem.rd_data_mem\[2\] sky130_fd_sc_hd__dlxtn_1
XFILLER_0_59_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21650_ _08672_ _08890_ _08894_ _08898_ VGND VGND VPWR VPWR _08899_ sky130_fd_sc_hd__and4_1
XFILLER_0_8_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30848_ clknet_leaf_223_clk _02583_ VGND VGND VPWR VPWR datamem.data_ram\[43\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20601_ _07889_ _07890_ _07891_ _07154_ VGND VGND VPWR VPWR _07892_ sky130_fd_sc_hd__a31o_1
X_21581_ _08511_ _08832_ VGND VGND VPWR VPWR _08833_ sky130_fd_sc_hd__nor2_1
X_30779_ clknet_leaf_192_clk _02514_ VGND VGND VPWR VPWR datamem.data_ram\[46\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20532_ _06605_ VGND VGND VPWR VPWR _07823_ sky130_fd_sc_hd__clkbuf_8
X_32518_ clknet_leaf_82_clk _03940_ VGND VGND VPWR VPWR datamem.data_ram\[24\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_201_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20463_ datamem.data_ram\[22\]\[20\] _07085_ _06646_ datamem.data_ram\[16\]\[20\]
+ _07754_ VGND VGND VPWR VPWR _07755_ sky130_fd_sc_hd__o221a_1
X_32449_ clknet_leaf_248_clk _03871_ VGND VGND VPWR VPWR datamem.data_ram\[27\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22202_ _09276_ net3910 _09371_ VGND VGND VPWR VPWR _09374_ sky130_fd_sc_hd__mux2_1
X_20394_ datamem.data_ram\[30\]\[28\] _06625_ _06684_ datamem.data_ram\[28\]\[28\]
+ VGND VGND VPWR VPWR _07686_ sky130_fd_sc_hd__o22a_1
XFILLER_0_207_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22133_ _09244_ net4079 _09332_ VGND VGND VPWR VPWR _09336_ sky130_fd_sc_hd__mux2_1
X_23531__158 clknet_1_1__leaf__10171_ VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__inv_2
X_27990_ _09278_ VGND VGND VPWR VPWR _12454_ sky130_fd_sc_hd__clkbuf_2
X_26941_ _11837_ _11842_ VGND VGND VPWR VPWR _11851_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22064_ _09281_ VGND VGND VPWR VPWR _09282_ sky130_fd_sc_hd__buf_2
XFILLER_0_227_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21015_ _07862_ _08303_ VGND VGND VPWR VPWR _08304_ sky130_fd_sc_hd__or2_1
X_26872_ _11795_ net1356 _11797_ _11806_ VGND VGND VPWR VPWR _03355_ sky130_fd_sc_hd__a31o_1
X_29660_ net1006 _01395_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[24\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_227_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25823_ _11208_ _11209_ VGND VGND VPWR VPWR _11210_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28611_ _12801_ VGND VGND VPWR VPWR _04099_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_226_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29591_ net945 _01326_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[26\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25754_ _11151_ VGND VGND VPWR VPWR _11157_ sky130_fd_sc_hd__buf_4
X_28542_ _12763_ VGND VGND VPWR VPWR _04068_ sky130_fd_sc_hd__clkbuf_1
X_22966_ clknet_1_0__leaf__10080_ VGND VGND VPWR VPWR _10082_ sky130_fd_sc_hd__buf_1
X_24705_ _10454_ net2083 _10552_ VGND VGND VPWR VPWR _10560_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28473_ _12458_ net3858 _12713_ VGND VGND VPWR VPWR _12719_ sky130_fd_sc_hd__mux2_1
X_21917_ _08626_ _09146_ _09148_ _09150_ _08808_ VGND VGND VPWR VPWR _09151_ sky130_fd_sc_hd__a221o_1
X_25685_ _11105_ net1672 _11111_ _11114_ VGND VGND VPWR VPWR _02860_ sky130_fd_sc_hd__a31o_1
XFILLER_0_168_946 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22897_ rvcpu.dp.rf.reg_file_arr\[0\]\[31\] rvcpu.dp.rf.reg_file_arr\[1\]\[31\] rvcpu.dp.rf.reg_file_arr\[2\]\[31\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[31\] _09477_ _09383_ VGND VGND VPWR VPWR _10032_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_139_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27424_ _12134_ net2372 _12126_ VGND VGND VPWR VPWR _12135_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24636_ _10385_ net3809 _10521_ VGND VGND VPWR VPWR _10522_ sky130_fd_sc_hd__mux2_1
X_21848_ _08835_ _09085_ VGND VGND VPWR VPWR _09086_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_216_5676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_216_5687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27355_ _09329_ VGND VGND VPWR VPWR _12095_ sky130_fd_sc_hd__buf_2
X_24567_ _10442_ net3522 _10482_ VGND VGND VPWR VPWR _10484_ sky130_fd_sc_hd__mux2_1
X_21779_ _08672_ _09012_ _09016_ _09020_ VGND VGND VPWR VPWR _09021_ sky130_fd_sc_hd__and4_1
XFILLER_0_93_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26306_ net1802 _11478_ VGND VGND VPWR VPWR _11486_ sky130_fd_sc_hd__and2_1
XFILLER_0_154_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23518_ _10167_ VGND VGND VPWR VPWR _01640_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27286_ _11968_ _12054_ VGND VGND VPWR VPWR _12056_ sky130_fd_sc_hd__and2_1
XFILLER_0_191_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24498_ _09351_ _10337_ _10366_ VGND VGND VPWR VPWR _10440_ sky130_fd_sc_hd__a21oi_4
X_23692__287 clknet_1_1__leaf__10195_ VGND VGND VPWR VPWR net413 sky130_fd_sc_hd__inv_2
XFILLER_0_68_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29025_ _13024_ VGND VGND VPWR VPWR _04290_ sky130_fd_sc_hd__clkbuf_1
X_26237_ _11379_ _03043_ _11454_ VGND VGND VPWR VPWR _03070_ sky130_fd_sc_hd__a21o_1
XFILLER_0_184_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26168_ _09478_ _11362_ VGND VGND VPWR VPWR _11421_ sky130_fd_sc_hd__and2_1
X_25119_ _10737_ net2095 _10784_ VGND VGND VPWR VPWR _10791_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26099_ _11384_ VGND VGND VPWR VPWR _03003_ sky130_fd_sc_hd__clkbuf_1
X_18990_ _05305_ _05562_ _05641_ _05655_ VGND VGND VPWR VPWR _06325_ sky130_fd_sc_hd__a31oi_1
XTAP_TAPCELL_ROW_167_4495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17941_ rvcpu.dp.plde.RD1E\[15\] _05267_ _05271_ _13231_ _05312_ VGND VGND VPWR VPWR
+ _05313_ sky130_fd_sc_hd__a221o_2
XFILLER_0_29_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29927_ net297 _01662_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[16\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_109_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_109_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_11__f_clk clknet_2_1_0_clk VGND VGND VPWR VPWR clknet_5_11__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_17872_ rvcpu.dp.plem.RdM\[3\] VGND VGND VPWR VPWR _05245_ sky130_fd_sc_hd__inv_2
X_29858_ net236 _01593_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[18\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19611_ _06680_ _06899_ _06901_ _06906_ VGND VGND VPWR VPWR _06907_ sky130_fd_sc_hd__a31o_1
XFILLER_0_40_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_219_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16823_ _04647_ VGND VGND VPWR VPWR _04659_ sky130_fd_sc_hd__buf_4
X_28809_ _12690_ net2669 _12905_ VGND VGND VPWR VPWR _12907_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_105_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29789_ net1135 _01524_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[20\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31820_ clknet_leaf_104_clk _03274_ VGND VGND VPWR VPWR datamem.data_ram\[9\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_19542_ datamem.data_ram\[24\]\[24\] _06837_ _06806_ datamem.data_ram\[28\]\[24\]
+ VGND VGND VPWR VPWR _06838_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_176_4709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16754_ _04622_ VGND VGND VPWR VPWR _01666_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_191_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_221_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15705_ _14174_ VGND VGND VPWR VPWR _02167_ sky130_fd_sc_hd__clkbuf_1
X_31751_ clknet_leaf_61_clk _03205_ VGND VGND VPWR VPWR datamem.data_ram\[45\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_19473_ _06732_ VGND VGND VPWR VPWR _06769_ sky130_fd_sc_hd__buf_8
X_16685_ _14149_ net3777 _04576_ VGND VGND VPWR VPWR _04586_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18424_ _05785_ _05787_ _05772_ VGND VGND VPWR VPWR _05788_ sky130_fd_sc_hd__a21o_1
X_30702_ clknet_leaf_217_clk _02437_ VGND VGND VPWR VPWR datamem.data_ram\[49\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15636_ _14126_ VGND VGND VPWR VPWR _02188_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_174_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31682_ clknet_5_1__leaf_clk net4316 VGND VGND VPWR VPWR rvcpu.dp.plmw.ALUResultW\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_139_3830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_3841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_415 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18355_ _05363_ _05375_ VGND VGND VPWR VPWR _05720_ sky130_fd_sc_hd__nand2_2
XFILLER_0_5_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30633_ clknet_leaf_219_clk _02368_ VGND VGND VPWR VPWR datamem.data_ram\[51\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_15567_ _13174_ rvcpu.dp.plmw.RdW\[3\] _13176_ VGND VGND VPWR VPWR _14089_ sky130_fd_sc_hd__or3b_2
XTAP_TAPCELL_ROW_29_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_3727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_3738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17306_ net4429 _13219_ _04913_ VGND VGND VPWR VPWR _04916_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30564_ clknet_leaf_199_clk _02299_ VGND VGND VPWR VPWR datamem.data_ram\[54\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_15498_ _13425_ _13847_ _13465_ _13513_ VGND VGND VPWR VPWR _14026_ sky130_fd_sc_hd__a211o_1
X_18286_ _05290_ _05647_ _05650_ VGND VGND VPWR VPWR _05651_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32303_ clknet_leaf_89_clk _03725_ VGND VGND VPWR VPWR datamem.data_ram\[32\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_25_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17237_ _14156_ net2579 _04876_ VGND VGND VPWR VPWR _04879_ sky130_fd_sc_hd__mux2_1
X_30495_ clknet_leaf_145_clk _02230_ VGND VGND VPWR VPWR datamem.data_ram\[57\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24109__616 clknet_1_0__leaf__10259_ VGND VGND VPWR VPWR net742 sky130_fd_sc_hd__inv_2
XFILLER_0_226_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold904 rvcpu.dp.rf.reg_file_arr\[5\]\[6\] VGND VGND VPWR VPWR net2054 sky130_fd_sc_hd__dlygate4sd3_1
X_17168_ _04842_ VGND VGND VPWR VPWR _01456_ sky130_fd_sc_hd__clkbuf_1
X_32234_ clknet_leaf_259_clk _03656_ VGND VGND VPWR VPWR datamem.data_ram\[35\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold915 rvcpu.dp.rf.reg_file_arr\[11\]\[28\] VGND VGND VPWR VPWR net2065 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold926 rvcpu.dp.rf.reg_file_arr\[8\]\[0\] VGND VGND VPWR VPWR net2076 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16119_ net2526 _13229_ _14396_ VGND VGND VPWR VPWR _14402_ sky130_fd_sc_hd__mux2_1
Xhold937 rvcpu.dp.rf.reg_file_arr\[3\]\[0\] VGND VGND VPWR VPWR net2087 sky130_fd_sc_hd__dlygate4sd3_1
X_32165_ clknet_leaf_242_clk _03587_ VGND VGND VPWR VPWR datamem.data_ram\[38\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold948 rvcpu.dp.rf.reg_file_arr\[30\]\[15\] VGND VGND VPWR VPWR net2098 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17099_ _14154_ net4233 _04804_ VGND VGND VPWR VPWR _04806_ sky130_fd_sc_hd__mux2_1
Xhold959 rvcpu.dp.rf.reg_file_arr\[11\]\[10\] VGND VGND VPWR VPWR net2109 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3006 datamem.data_ram\[23\]\[20\] VGND VGND VPWR VPWR net4156 sky130_fd_sc_hd__dlygate4sd3_1
X_31116_ clknet_leaf_61_clk _02851_ VGND VGND VPWR VPWR datamem.data_ram\[43\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3017 datamem.data_ram\[43\]\[21\] VGND VGND VPWR VPWR net4167 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3028 datamem.data_ram\[4\]\[19\] VGND VGND VPWR VPWR net4178 sky130_fd_sc_hd__dlygate4sd3_1
X_32096_ clknet_leaf_209_clk _03518_ VGND VGND VPWR VPWR datamem.data_ram\[8\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3039 datamem.data_ram\[15\]\[20\] VGND VGND VPWR VPWR net4189 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2305 rvcpu.dp.rf.reg_file_arr\[16\]\[10\] VGND VGND VPWR VPWR net3455 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2316 datamem.data_ram\[27\]\[28\] VGND VGND VPWR VPWR net3466 sky130_fd_sc_hd__dlygate4sd3_1
X_31047_ clknet_leaf_213_clk _02782_ VGND VGND VPWR VPWR datamem.data_ram\[9\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2327 datamem.data_ram\[25\]\[10\] VGND VGND VPWR VPWR net3477 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2338 datamem.data_ram\[35\]\[9\] VGND VGND VPWR VPWR net3488 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1604 datamem.data_ram\[45\]\[17\] VGND VGND VPWR VPWR net2754 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2349 datamem.data_ram\[22\]\[20\] VGND VGND VPWR VPWR net3499 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1615 datamem.data_ram\[17\]\[8\] VGND VGND VPWR VPWR net2765 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1626 datamem.data_ram\[15\]\[11\] VGND VGND VPWR VPWR net2776 sky130_fd_sc_hd__dlygate4sd3_1
X_19809_ datamem.data_ram\[5\]\[9\] _06724_ _06738_ datamem.data_ram\[3\]\[9\] _07103_
+ VGND VGND VPWR VPWR _07104_ sky130_fd_sc_hd__o221a_1
XFILLER_0_193_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1637 datamem.data_ram\[15\]\[23\] VGND VGND VPWR VPWR net2787 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1648 rvcpu.dp.rf.reg_file_arr\[27\]\[14\] VGND VGND VPWR VPWR net2798 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1659 datamem.data_ram\[33\]\[18\] VGND VGND VPWR VPWR net2809 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22820_ _09957_ _09958_ _09380_ VGND VGND VPWR VPWR _09959_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_212_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_224_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24155__658 clknet_1_0__leaf__10263_ VGND VGND VPWR VPWR net784 sky130_fd_sc_hd__inv_2
XFILLER_0_205_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_189_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22751_ rvcpu.dp.rf.reg_file_arr\[4\]\[23\] rvcpu.dp.rf.reg_file_arr\[5\]\[23\] rvcpu.dp.rf.reg_file_arr\[6\]\[23\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[23\] _09416_ _09716_ VGND VGND VPWR VPWR _09894_
+ sky130_fd_sc_hd__mux4_1
X_31949_ clknet_leaf_92_clk _03371_ VGND VGND VPWR VPWR datamem.data_ram\[32\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_91_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_91_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_149_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21702_ rvcpu.dp.rf.reg_file_arr\[4\]\[16\] rvcpu.dp.rf.reg_file_arr\[5\]\[16\] rvcpu.dp.rf.reg_file_arr\[6\]\[16\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[16\] _08839_ _08840_ VGND VGND VPWR VPWR _08948_
+ sky130_fd_sc_hd__mux4_1
X_25470_ _10055_ VGND VGND VPWR VPWR _10991_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22682_ _09481_ _09828_ VGND VGND VPWR VPWR _09829_ sky130_fd_sc_hd__and2_1
XFILLER_0_137_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24421_ _09278_ VGND VGND VPWR VPWR _10392_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21633_ rvcpu.dp.rf.reg_file_arr\[16\]\[13\] rvcpu.dp.rf.reg_file_arr\[17\]\[13\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[13\] rvcpu.dp.rf.reg_file_arr\[19\]\[13\] _08524_
+ _08800_ VGND VGND VPWR VPWR _08882_ sky130_fd_sc_hd__mux4_1
XFILLER_0_212_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_1326 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27140_ _10063_ VGND VGND VPWR VPWR _11972_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23302__944 clknet_1_1__leaf__10132_ VGND VGND VPWR VPWR net1070 sky130_fd_sc_hd__inv_2
XFILLER_0_75_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24352_ _10353_ VGND VGND VPWR VPWR _02288_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_192_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21564_ _08523_ VGND VGND VPWR VPWR _08817_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_211_5551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_211_5562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23303_ clknet_1_1__leaf__10130_ VGND VGND VPWR VPWR _10133_ sky130_fd_sc_hd__buf_1
X_27071_ _11919_ net1632 _11923_ _11928_ VGND VGND VPWR VPWR _03432_ sky130_fd_sc_hd__a31o_1
X_20515_ _06604_ _07803_ _07805_ _06916_ VGND VGND VPWR VPWR _07806_ sky130_fd_sc_hd__a31o_1
XFILLER_0_172_481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24283_ _10314_ VGND VGND VPWR VPWR _02258_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21495_ _08511_ _08750_ VGND VGND VPWR VPWR _08751_ sky130_fd_sc_hd__nor2_1
X_26022_ rvcpu.c.ad.funct7b5 _11329_ _11325_ _11336_ VGND VGND VPWR VPWR _02975_ sky130_fd_sc_hd__o211a_1
XFILLER_0_144_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20446_ datamem.data_ram\[5\]\[20\] _06702_ _06706_ datamem.data_ram\[7\]\[20\] VGND
+ VGND VPWR VPWR _07738_ sky130_fd_sc_hd__o22a_1
XFILLER_0_160_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20377_ datamem.data_ram\[58\]\[28\] _06802_ _06695_ datamem.data_ram\[56\]\[28\]
+ VGND VGND VPWR VPWR _07669_ sky130_fd_sc_hd__o22a_1
XFILLER_0_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22116_ rvcpu.dp.plem.WriteDataM\[6\] _08488_ _09293_ VGND VGND VPWR VPWR _09324_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_101_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_219_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27973_ _12442_ VGND VGND VPWR VPWR _03820_ sky130_fd_sc_hd__clkbuf_1
X_23728__320 clknet_1_1__leaf__10198_ VGND VGND VPWR VPWR net446 sky130_fd_sc_hd__inv_2
XFILLER_0_100_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29712_ net1058 _01447_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[22\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_26924_ _11840_ VGND VGND VPWR VPWR _11841_ sky130_fd_sc_hd__buf_2
X_22047_ _09227_ net112 VGND VGND VPWR VPWR _09269_ sky130_fd_sc_hd__nor2_8
XTAP_TAPCELL_ROW_162_4381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2850 datamem.data_ram\[33\]\[11\] VGND VGND VPWR VPWR net4000 sky130_fd_sc_hd__dlygate4sd3_1
X_29643_ net989 _01378_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[24\]\[6\] sky130_fd_sc_hd__dfxtp_1
Xhold2861 datamem.data_ram\[7\]\[14\] VGND VGND VPWR VPWR net4011 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_214_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26855_ _11725_ _11039_ VGND VGND VPWR VPWR _11796_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_162_4392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23430__82 clknet_1_1__leaf__10154_ VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__inv_2
Xhold2872 datamem.data_ram\[41\]\[27\] VGND VGND VPWR VPWR net4022 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_214_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2883 datamem.data_ram\[12\]\[10\] VGND VGND VPWR VPWR net4033 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2894 rvcpu.dp.rf.reg_file_arr\[14\]\[23\] VGND VGND VPWR VPWR net4044 sky130_fd_sc_hd__dlygate4sd3_1
X_25806_ net1650 _11181_ _11177_ _11196_ VGND VGND VPWR VPWR _02899_ sky130_fd_sc_hd__o211a_1
X_26786_ _11753_ net1618 _11748_ _11755_ VGND VGND VPWR VPWR _03320_ sky130_fd_sc_hd__a31o_1
XFILLER_0_199_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29574_ net928 _01309_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[26\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_833 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_218_5716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_218_5727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_218_5738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25737_ _11142_ VGND VGND VPWR VPWR _11143_ sky130_fd_sc_hd__clkbuf_4
X_28525_ _12279_ _10114_ _12668_ VGND VGND VPWR VPWR _12752_ sky130_fd_sc_hd__a21oi_4
X_22949_ _10075_ VGND VGND VPWR VPWR _10076_ sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_82_clk clknet_5_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_82_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16470_ net3166 _14430_ _04467_ VGND VGND VPWR VPWR _04472_ sky130_fd_sc_hd__mux2_1
X_25668_ _11085_ net2072 _11097_ _11102_ VGND VGND VPWR VPWR _02855_ sky130_fd_sc_hd__a31o_1
X_28456_ _12441_ net3294 _12704_ VGND VGND VPWR VPWR _12710_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_171_4606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15421_ _13298_ _13341_ _13336_ _13333_ VGND VGND VPWR VPWR _13953_ sky130_fd_sc_hd__o211a_1
XFILLER_0_210_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24619_ _10512_ VGND VGND VPWR VPWR _02396_ sky130_fd_sc_hd__clkbuf_1
X_27407_ _12123_ VGND VGND VPWR VPWR _03573_ sky130_fd_sc_hd__clkbuf_1
X_28387_ _12430_ net4087 _12669_ VGND VGND VPWR VPWR _12670_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25599_ _10418_ _11055_ VGND VGND VPWR VPWR _11063_ sky130_fd_sc_hd__and2_1
XFILLER_0_167_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23774__362 clknet_1_1__leaf__10202_ VGND VGND VPWR VPWR net488 sky130_fd_sc_hd__inv_2
XFILLER_0_182_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15352_ _13874_ _13875_ _13877_ _13887_ VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__o31a_1
X_18140_ rvcpu.dp.plde.RD1E\[16\] _05265_ _05269_ _13228_ _05505_ VGND VGND VPWR VPWR
+ _05506_ sky130_fd_sc_hd__a221o_4
X_27338_ _12083_ net3443 _12081_ VGND VGND VPWR VPWR _12084_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18071_ _05311_ _05318_ _05436_ _05438_ VGND VGND VPWR VPWR _05439_ sky130_fd_sc_hd__nand4_1
X_15283_ _13821_ VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_1
X_27269_ _10816_ net3715 _12043_ VGND VGND VPWR VPWR _12046_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_130_3613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17022_ net3045 _14436_ _04757_ VGND VGND VPWR VPWR _04765_ sky130_fd_sc_hd__mux2_1
X_29008_ _10066_ _13010_ VGND VGND VPWR VPWR _13015_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_130_3624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_169_4546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30280_ clknet_leaf_144_clk _02015_ VGND VGND VPWR VPWR datamem.data_ram\[58\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_169_4557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_91_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18973_ _05305_ _05641_ _05655_ _06308_ VGND VGND VPWR VPWR _06309_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_91_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17924_ rvcpu.dp.plde.ImmExtE\[29\] rvcpu.dp.SrcBFW_Mux.y\[29\] _05279_ VGND VGND
+ VPWR VPWR _05297_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_3564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_3575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32921_ clknet_leaf_262_clk _04343_ VGND VGND VPWR VPWR datamem.data_ram\[0\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_17855_ _05231_ VGND VGND VPWR VPWR rvcpu.dp.SrcBFW_Mux.y\[9\] sky130_fd_sc_hd__buf_1
XFILLER_0_227_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16806_ _04650_ VGND VGND VPWR VPWR _01634_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_205_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32852_ clknet_leaf_233_clk _04274_ VGND VGND VPWR VPWR datamem.data_ram\[11\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_17786_ net1581 _05178_ _05181_ _05182_ VGND VGND VPWR VPWR rvcpu.dp.SrcBFW_Mux.y\[1\]
+ sky130_fd_sc_hd__o22a_1
X_23480__127 clknet_1_0__leaf__10159_ VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_50_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14998_ _13287_ _13391_ VGND VGND VPWR VPWR _13546_ sky130_fd_sc_hd__nor2_4
XFILLER_0_205_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_220_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31803_ clknet_leaf_98_clk _03257_ VGND VGND VPWR VPWR datamem.data_ram\[46\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19525_ _06820_ VGND VGND VPWR VPWR _06821_ sky130_fd_sc_hd__buf_8
X_16737_ net2641 _14424_ _04612_ VGND VGND VPWR VPWR _04614_ sky130_fd_sc_hd__mux2_1
X_32783_ clknet_leaf_157_clk _04205_ VGND VGND VPWR VPWR datamem.data_ram\[14\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_73_clk clknet_5_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_73_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_163_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23560__184 clknet_1_1__leaf__10174_ VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__inv_2
X_19456_ _06751_ VGND VGND VPWR VPWR _06752_ sky130_fd_sc_hd__buf_8
X_31734_ net183 _03192_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[9\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16668_ _04577_ VGND VGND VPWR VPWR _01707_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18407_ rvcpu.dp.plde.RD1E\[0\] _05266_ _05270_ _13277_ _05393_ VGND VGND VPWR VPWR
+ _05771_ sky130_fd_sc_hd__a221o_2
XTAP_TAPCELL_ROW_27_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15619_ net3928 _13254_ _14114_ VGND VGND VPWR VPWR _14118_ sky130_fd_sc_hd__mux2_1
X_31665_ clknet_leaf_67_clk net1254 VGND VGND VPWR VPWR rvcpu.dp.plmw.ALUResultW\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_19387_ _06682_ VGND VGND VPWR VPWR _06683_ sky130_fd_sc_hd__buf_6
XFILLER_0_173_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16599_ _14127_ net2726 _04540_ VGND VGND VPWR VPWR _04541_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18338_ _05702_ VGND VGND VPWR VPWR _05703_ sky130_fd_sc_hd__buf_2
X_30616_ clknet_leaf_149_clk _02351_ VGND VGND VPWR VPWR datamem.data_ram\[52\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_31596_ clknet_leaf_51_clk net1182 VGND VGND VPWR VPWR rvcpu.dp.plmw.PCPlus4W\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30547_ clknet_leaf_139_clk _02282_ VGND VGND VPWR VPWR datamem.data_ram\[55\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_18269_ _05531_ _05633_ _05534_ VGND VGND VPWR VPWR _05634_ sky130_fd_sc_hd__or3_1
XFILLER_0_170_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20300_ datamem.data_ram\[7\]\[19\] _06761_ _07591_ _07592_ VGND VGND VPWR VPWR _07593_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_682 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21280_ _08541_ VGND VGND VPWR VPWR _08542_ sky130_fd_sc_hd__buf_4
Xhold701 datamem.data_ram\[62\]\[7\] VGND VGND VPWR VPWR net1851 sky130_fd_sc_hd__dlygate4sd3_1
X_30478_ net156 _02213_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[19\]\[25\] sky130_fd_sc_hd__dfxtp_1
Xhold712 rvcpu.dp.pcreg.q\[20\] VGND VGND VPWR VPWR net1862 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold723 datamem.data_ram\[41\]\[31\] VGND VGND VPWR VPWR net1873 sky130_fd_sc_hd__dlygate4sd3_1
X_20231_ datamem.data_ram\[7\]\[3\] _06925_ _06947_ datamem.data_ram\[1\]\[3\] VGND
+ VGND VPWR VPWR _07524_ sky130_fd_sc_hd__a22o_1
X_32217_ clknet_leaf_226_clk _03639_ VGND VGND VPWR VPWR datamem.data_ram\[35\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold734 rvcpu.dp.plfd.PCD\[5\] VGND VGND VPWR VPWR net1884 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_203_Left_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold745 datamem.data_ram\[35\]\[22\] VGND VGND VPWR VPWR net1895 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_57_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold756 rvcpu.dp.rf.reg_file_arr\[5\]\[3\] VGND VGND VPWR VPWR net1906 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold767 rvcpu.dp.rf.reg_file_arr\[10\]\[31\] VGND VGND VPWR VPWR net1917 sky130_fd_sc_hd__dlygate4sd3_1
Xhold778 datamem.data_ram\[35\]\[1\] VGND VGND VPWR VPWR net1928 sky130_fd_sc_hd__dlygate4sd3_1
X_20162_ datamem.data_ram\[16\]\[27\] _06695_ _06725_ datamem.data_ram\[23\]\[27\]
+ VGND VGND VPWR VPWR _07455_ sky130_fd_sc_hd__o22a_1
X_32148_ clknet_leaf_225_clk _03570_ VGND VGND VPWR VPWR datamem.data_ram\[38\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold789 rvcpu.dp.rf.reg_file_arr\[7\]\[20\] VGND VGND VPWR VPWR net1939 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2102 datamem.data_ram\[63\]\[18\] VGND VGND VPWR VPWR net3252 sky130_fd_sc_hd__dlygate4sd3_1
X_24970_ _10704_ VGND VGND VPWR VPWR _02555_ sky130_fd_sc_hd__clkbuf_1
X_20093_ datamem.data_ram\[59\]\[10\] _06828_ _07386_ _06851_ VGND VGND VPWR VPWR
+ _07387_ sky130_fd_sc_hd__o211a_1
Xhold2113 datamem.data_ram\[18\]\[30\] VGND VGND VPWR VPWR net3263 sky130_fd_sc_hd__dlygate4sd3_1
X_32079_ clknet_leaf_93_clk _03501_ VGND VGND VPWR VPWR datamem.data_ram\[33\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2124 rvcpu.dp.rf.reg_file_arr\[31\]\[7\] VGND VGND VPWR VPWR net3274 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2135 datamem.data_ram\[62\]\[28\] VGND VGND VPWR VPWR net3285 sky130_fd_sc_hd__dlygate4sd3_1
X_23944__498 clknet_1_1__leaf__10228_ VGND VGND VPWR VPWR net624 sky130_fd_sc_hd__inv_2
Xhold1401 rvcpu.dp.rf.reg_file_arr\[1\]\[19\] VGND VGND VPWR VPWR net2551 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2146 datamem.data_ram\[18\]\[26\] VGND VGND VPWR VPWR net3296 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2157 datamem.data_ram\[27\]\[12\] VGND VGND VPWR VPWR net3307 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1412 rvcpu.dp.rf.reg_file_arr\[30\]\[7\] VGND VGND VPWR VPWR net2562 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2168 datamem.data_ram\[40\]\[8\] VGND VGND VPWR VPWR net3318 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1423 datamem.data_ram\[23\]\[30\] VGND VGND VPWR VPWR net2573 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1434 datamem.data_ram\[58\]\[25\] VGND VGND VPWR VPWR net2584 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2179 datamem.data_ram\[24\]\[31\] VGND VGND VPWR VPWR net3329 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1445 datamem.data_ram\[41\]\[14\] VGND VGND VPWR VPWR net2595 sky130_fd_sc_hd__dlygate4sd3_1
X_26640_ _11083_ _11663_ VGND VGND VPWR VPWR _11667_ sky130_fd_sc_hd__and2_1
Xhold1456 rvcpu.dp.rf.reg_file_arr\[21\]\[12\] VGND VGND VPWR VPWR net2606 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_225_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_174_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1467 rvcpu.dp.rf.reg_file_arr\[2\]\[18\] VGND VGND VPWR VPWR net2617 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_212_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1478 rvcpu.dp.rf.reg_file_arr\[28\]\[22\] VGND VGND VPWR VPWR net2628 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_200_5285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1489 datamem.data_ram\[41\]\[10\] VGND VGND VPWR VPWR net2639 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__10240_ _10240_ VGND VGND VPWR VPWR clknet_0__10240_ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_200_5296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22803_ _09442_ _09938_ _09940_ _09942_ VGND VGND VPWR VPWR _09943_ sky130_fd_sc_hd__o2bb2a_1
X_26571_ _10727_ net3222 _11629_ VGND VGND VPWR VPWR _11631_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1__f__10140_ clknet_0__10140_ VGND VGND VPWR VPWR clknet_1_1__leaf__10140_
+ sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_212_Left_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20995_ _06594_ _08276_ _08283_ VGND VGND VPWR VPWR _08284_ sky130_fd_sc_hd__or3_1
XFILLER_0_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_64_clk clknet_5_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_64_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25522_ _10991_ net1381 _11009_ _11017_ VGND VGND VPWR VPWR _02794_ sky130_fd_sc_hd__a31o_1
Xclkbuf_0__10171_ _10171_ VGND VGND VPWR VPWR clknet_0__10171_ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_0_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28310_ _12628_ VGND VGND VPWR VPWR _03971_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_177_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29290_ _13166_ VGND VGND VPWR VPWR _04413_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_0_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22734_ _09636_ _09877_ VGND VGND VPWR VPWR _09878_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_0_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_213_5602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_192_5097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_213_5613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28241_ _12443_ net4345 _12583_ VGND VGND VPWR VPWR _12590_ sky130_fd_sc_hd__mux2_1
X_25453_ _10782_ _10981_ _10982_ net1307 VGND VGND VPWR VPWR _02760_ sky130_fd_sc_hd__a22o_1
X_23226__875 clknet_1_0__leaf__10125_ VGND VGND VPWR VPWR net1001 sky130_fd_sc_hd__inv_2
X_22665_ _09627_ _09810_ _09812_ _09795_ VGND VGND VPWR VPWR _09813_ sky130_fd_sc_hd__a211o_1
XFILLER_0_164_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24404_ _10381_ VGND VGND VPWR VPWR _02312_ sky130_fd_sc_hd__clkbuf_1
X_21616_ rvcpu.dp.rf.reg_file_arr\[20\]\[12\] rvcpu.dp.rf.reg_file_arr\[21\]\[12\]
+ rvcpu.dp.rf.reg_file_arr\[22\]\[12\] rvcpu.dp.rf.reg_file_arr\[23\]\[12\] _08516_
+ _08518_ VGND VGND VPWR VPWR _08866_ sky130_fd_sc_hd__mux4_1
X_28172_ _12369_ net2676 _12546_ VGND VGND VPWR VPWR _12553_ sky130_fd_sc_hd__mux2_1
X_25384_ _10418_ _10936_ VGND VGND VPWR VPWR _10944_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22596_ _09391_ _09746_ VGND VGND VPWR VPWR _09747_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27123_ _11956_ net1804 _11952_ _11960_ VGND VGND VPWR VPWR _03452_ sky130_fd_sc_hd__a31o_1
X_24335_ _09252_ net4308 _10338_ VGND VGND VPWR VPWR _10344_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21547_ _08526_ VGND VGND VPWR VPWR _08800_ sky130_fd_sc_hd__buf_4
X_23537__164 clknet_1_1__leaf__10171_ VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__inv_2
XFILLER_0_181_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27054_ _11904_ net1848 _11910_ _11917_ VGND VGND VPWR VPWR _03426_ sky130_fd_sc_hd__a31o_1
XFILLER_0_65_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24266_ _10305_ VGND VGND VPWR VPWR _02250_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_221_Left_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_209_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21478_ _08663_ _08732_ _08734_ _08652_ VGND VGND VPWR VPWR _08735_ sky130_fd_sc_hd__o211a_1
XFILLER_0_181_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26005_ net16 _11153_ _11325_ _11327_ VGND VGND VPWR VPWR _02967_ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20429_ datamem.data_ram\[11\]\[12\] _06632_ _06780_ datamem.data_ram\[9\]\[12\]
+ VGND VGND VPWR VPWR _07721_ sky130_fd_sc_hd__o22a_1
XFILLER_0_132_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_164_4421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_164_4432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_4443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27956_ _12178_ _12335_ _12356_ VGND VGND VPWR VPWR _12431_ sky130_fd_sc_hd__a21oi_4
X_23079_ _10101_ VGND VGND VPWR VPWR _01267_ sky130_fd_sc_hd__clkbuf_1
X_15970_ _14310_ VGND VGND VPWR VPWR _14322_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_160_4329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14921_ _13341_ _13336_ VGND VGND VPWR VPWR _13470_ sky130_fd_sc_hd__nor2_1
X_26907_ _10063_ VGND VGND VPWR VPWR _11829_ sky130_fd_sc_hd__clkbuf_4
X_27887_ _10209_ _10049_ _11898_ VGND VGND VPWR VPWR _12394_ sky130_fd_sc_hd__and3_2
Xhold50 rvcpu.dp.plde.PCPlus4E\[25\] VGND VGND VPWR VPWR net1200 sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 rvcpu.dp.plem.lAuiPCM\[6\] VGND VGND VPWR VPWR net1211 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2680 datamem.data_ram\[47\]\[18\] VGND VGND VPWR VPWR net3830 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 rvcpu.dp.plem.PCPlus4M\[0\] VGND VGND VPWR VPWR net1222 sky130_fd_sc_hd__dlygate4sd3_1
X_29626_ net980 _01361_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[25\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17640_ _05092_ VGND VGND VPWR VPWR _01218_ sky130_fd_sc_hd__clkbuf_1
X_26838_ _11676_ _11786_ VGND VGND VPWR VPWR _11787_ sky130_fd_sc_hd__and2_1
Xhold83 rvcpu.dp.plem.PCPlus4M\[15\] VGND VGND VPWR VPWR net1233 sky130_fd_sc_hd__dlygate4sd3_1
X_14852_ _13368_ _13396_ _13404_ VGND VGND VPWR VPWR _13405_ sky130_fd_sc_hd__o21ai_1
Xhold2691 datamem.data_ram\[49\]\[10\] VGND VGND VPWR VPWR net3841 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 rvcpu.dp.plem.lAuiPCM\[13\] VGND VGND VPWR VPWR net1244 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_202_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_3450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26499__52 clknet_1_0__leaf__11601_ VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__inv_2
XFILLER_0_216_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1990 datamem.data_ram\[31\]\[19\] VGND VGND VPWR VPWR net3140 sky130_fd_sc_hd__dlygate4sd3_1
X_14783_ rvcpu.dp.pcreg.q\[5\] rvcpu.dp.pcreg.q\[2\] VGND VGND VPWR VPWR _13336_ sky130_fd_sc_hd__nand2_8
X_29557_ net911 _01292_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[27\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_17571_ _13210_ net2628 _05046_ VGND VGND VPWR VPWR _05056_ sky130_fd_sc_hd__mux2_1
X_26769_ _11735_ net1683 _11737_ _11744_ VGND VGND VPWR VPWR _03314_ sky130_fd_sc_hd__a31o_1
XFILLER_0_202_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_63_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_55_clk clknet_5_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_55_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_63_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19310_ _06584_ rvcpu.dp.plem.ALUResultM\[3\] VGND VGND VPWR VPWR _06606_ sky130_fd_sc_hd__nand2_8
X_16522_ net1932 _14482_ _04489_ VGND VGND VPWR VPWR _04499_ sky130_fd_sc_hd__mux2_1
X_28508_ _12740_ VGND VGND VPWR VPWR _04057_ sky130_fd_sc_hd__clkbuf_1
X_29488_ net850 _01223_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[2\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23698__293 clknet_1_0__leaf__10195_ VGND VGND VPWR VPWR net419 sky130_fd_sc_hd__inv_2
XFILLER_0_168_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_195_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19241_ _06545_ rvcpu.dp.plde.ImmExtE\[28\] _06493_ VGND VGND VPWR VPWR _06546_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16453_ _04461_ VGND VGND VPWR VPWR _01814_ sky130_fd_sc_hd__clkbuf_1
X_28439_ _09325_ VGND VGND VPWR VPWR _12700_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_151_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15404_ _13402_ _13505_ _13737_ _13431_ VGND VGND VPWR VPWR _13936_ sky130_fd_sc_hd__a22o_1
X_19172_ _06485_ VGND VGND VPWR VPWR rvcpu.dp.lAuiPCE\[19\] sky130_fd_sc_hd__clkbuf_1
X_31450_ clknet_leaf_2_clk rvcpu.dp.SrcBFW_Mux.y\[8\] VGND VGND VPWR VPWR rvcpu.dp.plem.WriteDataM\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_16384_ net2162 _14482_ _14547_ VGND VGND VPWR VPWR _14557_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_22_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_307 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15335_ _13849_ _13861_ _13871_ VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__a21oi_1
XFILLER_0_137_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18123_ rvcpu.dp.plde.RD1E\[18\] _05292_ _05489_ VGND VGND VPWR VPWR _05490_ sky130_fd_sc_hd__o21a_2
XTAP_TAPCELL_ROW_22_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30401_ net739 _02136_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[31\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_186_1278 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31381_ clknet_leaf_21_clk _03084_ VGND VGND VPWR VPWR rvcpu.dp.plde.ImmExtE\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15266_ _13431_ _13589_ VGND VGND VPWR VPWR _13805_ sky130_fd_sc_hd__nand2_1
X_18054_ rvcpu.dp.plem.ALUResultM\[8\] _05422_ _05177_ VGND VGND VPWR VPWR _05423_
+ sky130_fd_sc_hd__mux2_1
X_30332_ net678 _02067_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[4\]\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_93_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_298 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_3 _01133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_1_0__f__10160_ clknet_0__10160_ VGND VGND VPWR VPWR clknet_1_0__leaf__10160_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_112_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17005_ _13174_ _13175_ _13176_ VGND VGND VPWR VPWR _04755_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_188_4999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30263_ net617 _01998_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[6\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_15197_ _13706_ _13459_ _13348_ _13737_ _13738_ VGND VGND VPWR VPWR _13739_ sky130_fd_sc_hd__a41o_1
XFILLER_0_151_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_663 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__10091_ clknet_0__10091_ VGND VGND VPWR VPWR clknet_1_0__leaf__10091_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_5_9__f_clk clknet_2_1_0_clk VGND VGND VPWR VPWR clknet_5_9__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_32002_ clknet_leaf_133_clk _03424_ VGND VGND VPWR VPWR datamem.data_ram\[52\]\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_21_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30194_ net548 _01929_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[8\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18956_ _05543_ _05547_ _06291_ VGND VGND VPWR VPWR _06293_ sky130_fd_sc_hd__or3_1
XFILLER_0_225_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23331__970 clknet_1_0__leaf__10135_ VGND VGND VPWR VPWR net1096 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_52_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17907_ rvcpu.dp.plde.ImmExtE\[31\] rvcpu.dp.SrcBFW_Mux.y\[31\] _05279_ VGND VGND
+ VPWR VPWR _05280_ sky130_fd_sc_hd__mux2_1
XFILLER_0_225_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18887_ _06055_ _06227_ _06228_ VGND VGND VPWR VPWR _06229_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_222_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32904_ clknet_leaf_208_clk _04326_ VGND VGND VPWR VPWR datamem.data_ram\[0\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_222_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_175_Right_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17838_ rvcpu.dp.plem.ALUResultM\[19\] _05219_ _05177_ VGND VGND VPWR VPWR _05220_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_206_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_179_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_179_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32835_ clknet_leaf_254_clk _04257_ VGND VGND VPWR VPWR datamem.data_ram\[12\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_222_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17769_ rvcpu.dp.plem.RdM\[1\] _05165_ rvcpu.dp.plde.Rs2E\[0\] _05162_ _05166_ VGND
+ VGND VPWR VPWR _05167_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_46_clk clknet_5_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_46_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_156_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19508_ _06803_ VGND VGND VPWR VPWR _06804_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_18_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32766_ clknet_leaf_283_clk _04188_ VGND VGND VPWR VPWR datamem.data_ram\[15\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_20780_ datamem.data_ram\[4\]\[30\] datamem.data_ram\[5\]\[30\] _07849_ VGND VGND
+ VPWR VPWR _08070_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_187_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19439_ datamem.data_ram\[37\]\[16\] _06724_ _06727_ _06734_ VGND VGND VPWR VPWR
+ _06735_ sky130_fd_sc_hd__o211a_1
X_31717_ net166 _03175_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[9\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32697_ clknet_leaf_244_clk _04119_ VGND VGND VPWR VPWR datamem.data_ram\[17\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22450_ rvcpu.dp.rf.reg_file_arr\[8\]\[7\] rvcpu.dp.rf.reg_file_arr\[10\]\[7\] rvcpu.dp.rf.reg_file_arr\[9\]\[7\]
+ rvcpu.dp.rf.reg_file_arr\[11\]\[7\] _09608_ _09532_ VGND VGND VPWR VPWR _09609_
+ sky130_fd_sc_hd__mux4_1
X_31648_ clknet_leaf_25_clk net1155 VGND VGND VPWR VPWR rvcpu.dp.plmw.lAuiPCW\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21401_ _08627_ _08656_ _08658_ _08660_ VGND VGND VPWR VPWR _08661_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22381_ rvcpu.dp.rf.reg_file_arr\[16\]\[4\] rvcpu.dp.rf.reg_file_arr\[17\]\[4\] rvcpu.dp.rf.reg_file_arr\[18\]\[4\]
+ rvcpu.dp.rf.reg_file_arr\[19\]\[4\] _09406_ _09395_ VGND VGND VPWR VPWR _09543_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_72_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31579_ clknet_leaf_75_clk datamem.rd_data_mem\[29\] VGND VGND VPWR VPWR rvcpu.dp.plmw.ReadDataW\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21332_ rvcpu.dp.plfd.InstrD\[23\] _08582_ rvcpu.dp.plde.RdE\[4\] _08589_ _08593_
+ VGND VGND VPWR VPWR _08594_ sky130_fd_sc_hd__o221a_1
XFILLER_0_115_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold520 datamem.data_ram\[18\]\[0\] VGND VGND VPWR VPWR net1670 sky130_fd_sc_hd__dlygate4sd3_1
X_21263_ _08524_ VGND VGND VPWR VPWR _08525_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_206_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold531 datamem.data_ram\[13\]\[0\] VGND VGND VPWR VPWR net1681 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold542 rvcpu.dp.plfd.PCD\[22\] VGND VGND VPWR VPWR net1692 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold553 datamem.data_ram\[10\]\[5\] VGND VGND VPWR VPWR net1703 sky130_fd_sc_hd__dlygate4sd3_1
X_20214_ _06590_ _07506_ VGND VGND VPWR VPWR _07507_ sky130_fd_sc_hd__nor2_1
XFILLER_0_229_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold564 datamem.data_ram\[16\]\[3\] VGND VGND VPWR VPWR net1714 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold575 datamem.data_ram\[27\]\[0\] VGND VGND VPWR VPWR net1725 sky130_fd_sc_hd__dlygate4sd3_1
X_21194_ _07277_ net37 _07461_ _06915_ VGND VGND VPWR VPWR _08478_ sky130_fd_sc_hd__o22ai_1
Xhold586 rvcpu.dp.plfd.PCPlus4D\[12\] VGND VGND VPWR VPWR net1736 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold597 datamem.data_ram\[9\]\[3\] VGND VGND VPWR VPWR net1747 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_206_5450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1047 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27810_ _12145_ net3564 net78 VGND VGND VPWR VPWR _12348_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20145_ datamem.data_ram\[61\]\[27\] _06815_ _06781_ datamem.data_ram\[57\]\[27\]
+ VGND VGND VPWR VPWR _07438_ sky130_fd_sc_hd__o22a_1
X_28790_ _12734_ net3344 net70 VGND VGND VPWR VPWR _12897_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_202_5336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_202_5347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24953_ _10695_ VGND VGND VPWR VPWR _02547_ sky130_fd_sc_hd__clkbuf_1
X_27741_ _12130_ net3814 _12307_ VGND VGND VPWR VPWR _12310_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_198_5240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20076_ datamem.data_ram\[45\]\[10\] _07037_ _06837_ datamem.data_ram\[40\]\[10\]
+ _07369_ VGND VGND VPWR VPWR _07370_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_198_5251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1220 rvcpu.dp.rf.reg_file_arr\[27\]\[8\] VGND VGND VPWR VPWR net2370 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1231 rvcpu.dp.rf.reg_file_arr\[17\]\[14\] VGND VGND VPWR VPWR net2381 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1242 rvcpu.dp.rf.reg_file_arr\[1\]\[3\] VGND VGND VPWR VPWR net2392 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_142_Right_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1253 rvcpu.dp.rf.reg_file_arr\[10\]\[29\] VGND VGND VPWR VPWR net2403 sky130_fd_sc_hd__dlygate4sd3_1
X_27672_ _12085_ net4085 net51 VGND VGND VPWR VPWR _12273_ sky130_fd_sc_hd__mux2_1
X_24884_ _10658_ VGND VGND VPWR VPWR _02515_ sky130_fd_sc_hd__clkbuf_1
Xhold1264 datamem.data_ram\[6\]\[8\] VGND VGND VPWR VPWR net2414 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1275 rvcpu.dp.rf.reg_file_arr\[20\]\[10\] VGND VGND VPWR VPWR net2425 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_213_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_194_5148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29411_ clknet_leaf_290_clk _01146_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD2E\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_212_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_194_5159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26623_ _09231_ _11659_ VGND VGND VPWR VPWR _11660_ sky130_fd_sc_hd__nor2_2
Xhold1286 datamem.data_ram\[3\]\[8\] VGND VGND VPWR VPWR net2436 sky130_fd_sc_hd__dlygate4sd3_1
X_23835_ _09314_ net2577 _10210_ VGND VGND VPWR VPWR _10214_ sky130_fd_sc_hd__mux2_1
Xhold1297 rvcpu.dp.rf.reg_file_arr\[27\]\[11\] VGND VGND VPWR VPWR net2447 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_404 _06632_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_415 _06716_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_37_clk clknet_5_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_37_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_426 _06783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0__10223_ _10223_ VGND VGND VPWR VPWR clknet_0__10223_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_212_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26554_ _10814_ net3089 _11620_ VGND VGND VPWR VPWR _11622_ sky130_fd_sc_hd__mux2_1
X_29342_ clknet_leaf_206_clk _01077_ VGND VGND VPWR VPWR datamem.data_ram\[61\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_437 _06933_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23766_ clknet_1_1__leaf__10192_ VGND VGND VPWR VPWR _10202_ sky130_fd_sc_hd__buf_1
XANTENNA_448 _07860_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_200_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20978_ _07819_ _08265_ _08266_ _06641_ VGND VGND VPWR VPWR _08267_ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_459 _08634_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22717_ _09415_ _09859_ _09861_ _09489_ VGND VGND VPWR VPWR _09862_ sky130_fd_sc_hd__o211a_1
Xclkbuf_0__10154_ _10154_ VGND VGND VPWR VPWR clknet_0__10154_ sky130_fd_sc_hd__clkbuf_16
X_25505_ _11007_ VGND VGND VPWR VPWR _02787_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29273_ _13157_ VGND VGND VPWR VPWR _04405_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_193_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_109_Left_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25436_ _10974_ VGND VGND VPWR VPWR _02751_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__10085_ _10085_ VGND VGND VPWR VPWR clknet_0__10085_ sky130_fd_sc_hd__clkbuf_16
X_28224_ _12369_ net4159 net45 VGND VGND VPWR VPWR _12581_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_705 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22648_ _09705_ _09786_ _09791_ _09796_ VGND VGND VPWR VPWR _09797_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_153_4166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_211_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_153_4177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25367_ _07019_ _10932_ _10044_ VGND VGND VPWR VPWR _10933_ sky130_fd_sc_hd__or3_1
XFILLER_0_24_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_703 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28155_ _12460_ net4358 net73 VGND VGND VPWR VPWR _12544_ sky130_fd_sc_hd__mux2_1
X_22579_ rvcpu.dp.rf.reg_file_arr\[24\]\[14\] rvcpu.dp.rf.reg_file_arr\[25\]\[14\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[14\] rvcpu.dp.rf.reg_file_arr\[27\]\[14\] _09484_
+ _09431_ VGND VGND VPWR VPWR _09731_ sky130_fd_sc_hd__mux4_1
X_15120_ _13320_ VGND VGND VPWR VPWR _13665_ sky130_fd_sc_hd__clkbuf_4
X_27106_ _11837_ _11941_ VGND VGND VPWR VPWR _11950_ sky130_fd_sc_hd__and2_1
X_24318_ _10334_ VGND VGND VPWR VPWR _02273_ sky130_fd_sc_hd__clkbuf_1
X_28086_ _12507_ VGND VGND VPWR VPWR _03868_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25298_ _10760_ net3717 _10887_ VGND VGND VPWR VPWR _10892_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15051_ _13297_ _13526_ VGND VGND VPWR VPWR _13598_ sky130_fd_sc_hd__nand2_2
X_27037_ _11904_ net1574 _11897_ _11907_ VGND VGND VPWR VPWR _03419_ sky130_fd_sc_hd__a31o_1
XFILLER_0_161_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24249_ _09291_ net3773 _10288_ VGND VGND VPWR VPWR _10296_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23812__395 clknet_1_1__leaf__10207_ VGND VGND VPWR VPWR net521 sky130_fd_sc_hd__inv_2
XFILLER_0_160_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_3173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput5 net5 VGND VGND VPWR VPWR Instr[12] sky130_fd_sc_hd__buf_2
XFILLER_0_121_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_112_3184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_222_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_118_Left_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18810_ _06156_ VGND VGND VPWR VPWR _06157_ sky130_fd_sc_hd__inv_2
XFILLER_0_208_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_183_4885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19790_ _06743_ VGND VGND VPWR VPWR _07085_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_183_4896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28988_ _13003_ VGND VGND VPWR VPWR _04274_ sky130_fd_sc_hd__clkbuf_1
X_23053__753 clknet_1_1__leaf__10090_ VGND VGND VPWR VPWR net879 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_125_3501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18741_ _06085_ _06089_ _05654_ VGND VGND VPWR VPWR _06092_ sky130_fd_sc_hd__a21oi_1
X_27939_ _12355_ net3015 _12421_ VGND VGND VPWR VPWR _12422_ sky130_fd_sc_hd__mux2_1
X_15953_ _14313_ VGND VGND VPWR VPWR _02050_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_223_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14904_ _13317_ _13454_ VGND VGND VPWR VPWR _13455_ sky130_fd_sc_hd__nand2_1
X_18672_ _05798_ _06026_ _05696_ VGND VGND VPWR VPWR _06027_ sky130_fd_sc_hd__mux2_1
X_30950_ clknet_leaf_272_clk _02685_ VGND VGND VPWR VPWR datamem.data_ram\[3\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_121_3409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15884_ net2643 _13184_ _14275_ VGND VGND VPWR VPWR _14277_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23168__840 clknet_1_0__leaf__10110_ VGND VGND VPWR VPWR net966 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_86_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29609_ net963 _01344_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[25\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_17623_ net3027 _13183_ _05082_ VGND VGND VPWR VPWR _05084_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_86_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14835_ rvcpu.dp.pcreg.q\[3\] _13280_ VGND VGND VPWR VPWR _13388_ sky130_fd_sc_hd__or2_1
XFILLER_0_215_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_142_3892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30881_ clknet_leaf_264_clk _02616_ VGND VGND VPWR VPWR datamem.data_ram\[42\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_28_clk clknet_5_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_28_clk sky130_fd_sc_hd__clkbuf_8
X_32620_ clknet_leaf_253_clk _04042_ VGND VGND VPWR VPWR datamem.data_ram\[20\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17554_ _05047_ VGND VGND VPWR VPWR _01259_ sky130_fd_sc_hd__clkbuf_1
X_14766_ _13318_ VGND VGND VPWR VPWR _13319_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_175_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_127_Left_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16505_ _04490_ VGND VGND VPWR VPWR _01791_ sky130_fd_sc_hd__clkbuf_1
X_32551_ clknet_leaf_274_clk _03973_ VGND VGND VPWR VPWR datamem.data_ram\[23\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17485_ _13173_ net3696 _05010_ VGND VGND VPWR VPWR _05011_ sky130_fd_sc_hd__mux2_1
X_14697_ net2031 _13257_ _13245_ VGND VGND VPWR VPWR _13258_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19224_ _06529_ _06530_ VGND VGND VPWR VPWR _06531_ sky130_fd_sc_hd__xor2_1
X_31502_ clknet_leaf_23_clk rvcpu.dp.lAuiPCE\[28\] VGND VGND VPWR VPWR rvcpu.dp.plem.lAuiPCM\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_3349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16436_ net2109 _14466_ _04451_ VGND VGND VPWR VPWR _04453_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32482_ clknet_leaf_239_clk _03904_ VGND VGND VPWR VPWR datamem.data_ram\[25\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_45_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23969__505 clknet_1_0__leaf__10238_ VGND VGND VPWR VPWR net631 sky130_fd_sc_hd__inv_2
X_31433_ clknet_leaf_54_clk _03136_ VGND VGND VPWR VPWR datamem.data_ram\[14\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_19155_ _06463_ rvcpu.dp.plde.PCE\[16\] rvcpu.dp.plde.ImmExtE\[16\] VGND VGND VPWR
+ VPWR _06470_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_186_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16367_ _14548_ VGND VGND VPWR VPWR _01855_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18106_ rvcpu.dp.plem.ALUResultM\[20\] _05339_ _05340_ _13216_ VGND VGND VPWR VPWR
+ _05474_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_41_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15318_ _13366_ _13301_ _13426_ VGND VGND VPWR VPWR _13855_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_41_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19086_ _06400_ _06403_ _06409_ VGND VGND VPWR VPWR _06410_ sky130_fd_sc_hd__a21oi_1
X_31364_ clknet_leaf_24_clk _03067_ VGND VGND VPWR VPWR rvcpu.dp.plde.ImmExtE\[13\]
+ sky130_fd_sc_hd__dfxtp_2
X_16298_ net4326 _14463_ _14511_ VGND VGND VPWR VPWR _14512_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18037_ rvcpu.dp.plem.ALUResultM\[11\] _05272_ VGND VGND VPWR VPWR _05407_ sky130_fd_sc_hd__and2_1
X_30315_ net661 _02050_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[5\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_15249_ _13501_ _13566_ _13659_ _13787_ _13788_ VGND VGND VPWR VPWR _13789_ sky130_fd_sc_hd__o311a_1
XFILLER_0_169_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_495 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31295_ clknet_leaf_16_clk _02998_ VGND VGND VPWR VPWR rvcpu.dp.plde.RegWriteE sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_136_Left_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_99_Right_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30246_ net600 _01981_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[6\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30177_ clknet_leaf_205_clk _01912_ VGND VGND VPWR VPWR datamem.data_ram\[58\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_19988_ datamem.data_ram\[8\]\[2\] _06990_ _07278_ _07281_ VGND VGND VPWR VPWR _07282_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_226_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23486__133 clknet_1_0__leaf__10159_ VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__inv_2
XFILLER_0_10_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18939_ _05240_ _06264_ _06265_ _06277_ VGND VGND VPWR VPWR rvcpu.ALUResultE\[25\]
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_201_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21950_ _08673_ _09181_ VGND VGND VPWR VPWR _09182_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_206_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20901_ datamem.data_ram\[13\]\[22\] _07837_ _08190_ _07863_ VGND VGND VPWR VPWR
+ _08191_ sky130_fd_sc_hd__a211o_1
XFILLER_0_179_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21881_ _08510_ _09116_ VGND VGND VPWR VPWR _09117_ sky130_fd_sc_hd__nor2_1
XFILLER_0_171_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_19_clk clknet_5_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_19_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_145_Left_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20832_ _08108_ _08121_ _06604_ VGND VGND VPWR VPWR _08122_ sky130_fd_sc_hd__o21a_1
X_32818_ clknet_leaf_212_clk _04240_ VGND VGND VPWR VPWR datamem.data_ram\[12\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20763_ _07131_ _08045_ _08052_ _06596_ VGND VGND VPWR VPWR _08053_ sky130_fd_sc_hd__o211a_1
XFILLER_0_119_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32749_ clknet_leaf_233_clk _04171_ VGND VGND VPWR VPWR datamem.data_ram\[15\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_22502_ _09452_ _09657_ VGND VGND VPWR VPWR _09658_ sky130_fd_sc_hd__nor2_1
X_26270_ _11413_ VGND VGND VPWR VPWR _11467_ sky130_fd_sc_hd__buf_2
XFILLER_0_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20694_ datamem.data_ram\[62\]\[5\] _07159_ _07981_ _07984_ VGND VGND VPWR VPWR _07985_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_190_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25221_ _10754_ net3726 _10848_ VGND VGND VPWR VPWR _10850_ sky130_fd_sc_hd__mux2_1
X_22433_ _09429_ _09590_ _09592_ _09438_ VGND VGND VPWR VPWR _09593_ sky130_fd_sc_hd__a211o_1
XFILLER_0_73_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25152_ _10808_ VGND VGND VPWR VPWR _02633_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22364_ rvcpu.dp.rf.reg_file_arr\[0\]\[3\] rvcpu.dp.rf.reg_file_arr\[1\]\[3\] rvcpu.dp.rf.reg_file_arr\[2\]\[3\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[3\] _09417_ _09419_ VGND VGND VPWR VPWR _09527_ sky130_fd_sc_hd__mux4_1
XFILLER_0_143_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_154_Left_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23338__976 clknet_1_0__leaf__10136_ VGND VGND VPWR VPWR net1102 sky130_fd_sc_hd__inv_2
X_21315_ _08565_ _08571_ _08574_ _08576_ VGND VGND VPWR VPWR _08577_ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29960_ net330 _01695_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[15\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_25083_ _10733_ net3287 net89 VGND VGND VPWR VPWR _10773_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22295_ _09441_ _09459_ VGND VGND VPWR VPWR _09460_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_211_Right_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28911_ _12690_ net3465 _12959_ VGND VGND VPWR VPWR _12961_ sky130_fd_sc_hd__mux2_1
X_24034_ clknet_1_1__leaf__10078_ VGND VGND VPWR VPWR _10244_ sky130_fd_sc_hd__buf_1
Xhold350 datamem.data_ram\[3\]\[5\] VGND VGND VPWR VPWR net1500 sky130_fd_sc_hd__dlygate4sd3_1
X_21246_ _08491_ _08495_ _08508_ VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__nor3_1
XFILLER_0_229_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold361 datamem.data_ram\[13\]\[5\] VGND VGND VPWR VPWR net1511 sky130_fd_sc_hd__dlygate4sd3_1
X_29891_ net269 _01626_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[17\]\[22\] sky130_fd_sc_hd__dfxtp_1
Xhold372 datamem.data_ram\[15\]\[7\] VGND VGND VPWR VPWR net1522 sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 datamem.data_ram\[22\]\[0\] VGND VGND VPWR VPWR net1533 sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 datamem.data_ram\[1\]\[6\] VGND VGND VPWR VPWR net1544 sky130_fd_sc_hd__dlygate4sd3_1
X_28842_ _12924_ VGND VGND VPWR VPWR _04207_ sky130_fd_sc_hd__clkbuf_1
X_21177_ _08354_ _08465_ _06588_ VGND VGND VPWR VPWR _08466_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_225_5892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20128_ datamem.data_ram\[11\]\[27\] _06828_ _06656_ datamem.data_ram\[9\]\[27\]
+ VGND VGND VPWR VPWR _07421_ sky130_fd_sc_hd__o22a_1
X_28773_ _12751_ net2443 _12887_ VGND VGND VPWR VPWR _12888_ sky130_fd_sc_hd__mux2_1
XFILLER_0_176_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25985_ rvcpu.dp.plfd.InstrD\[13\] _11315_ _11312_ _11316_ VGND VGND VPWR VPWR _02958_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_221_5789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27724_ _12085_ net3018 net49 VGND VGND VPWR VPWR _12301_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20059_ _06600_ _07350_ _07352_ _06592_ VGND VGND VPWR VPWR _07353_ sky130_fd_sc_hd__a31o_1
X_24936_ _10686_ VGND VGND VPWR VPWR _02539_ sky130_fd_sc_hd__clkbuf_1
Xhold1050 rvcpu.dp.rf.reg_file_arr\[21\]\[18\] VGND VGND VPWR VPWR net2200 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_198_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_163_Left_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1061 rvcpu.dp.rf.reg_file_arr\[7\]\[23\] VGND VGND VPWR VPWR net2211 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1072 rvcpu.dp.rf.reg_file_arr\[20\]\[18\] VGND VGND VPWR VPWR net2222 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_159_4320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1083 datamem.data_ram\[30\]\[20\] VGND VGND VPWR VPWR net2233 sky130_fd_sc_hd__dlygate4sd3_1
X_27655_ _12147_ net2951 net79 VGND VGND VPWR VPWR _12264_ sky130_fd_sc_hd__mux2_1
X_24867_ _10649_ VGND VGND VPWR VPWR _02507_ sky130_fd_sc_hd__clkbuf_1
Xhold1094 rvcpu.dp.rf.reg_file_arr\[17\]\[24\] VGND VGND VPWR VPWR net2244 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_201 _09479_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_212 _09636_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_201_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_223 _10041_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26606_ _10811_ net3545 _11650_ VGND VGND VPWR VPWR _11651_ sky130_fd_sc_hd__mux2_1
X_14620_ _13199_ VGND VGND VPWR VPWR _03198_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_234 _10209_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_212_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_245 _11965_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_4206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27586_ _12130_ net2151 _12224_ VGND VGND VPWR VPWR _12227_ sky130_fd_sc_hd__mux2_1
X_24798_ _10297_ _10337_ _10611_ VGND VGND VPWR VPWR _10612_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_169_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_4217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0__10206_ _10206_ VGND VGND VPWR VPWR clknet_0__10206_ sky130_fd_sc_hd__clkbuf_16
XANTENNA_256 _13200_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29325_ clknet_leaf_144_clk _01060_ VGND VGND VPWR VPWR datamem.data_ram\[62\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_267 _13225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_1_1__f__10106_ clknet_0__10106_ VGND VGND VPWR VPWR clknet_1_1__leaf__10106_
+ sky130_fd_sc_hd__clkbuf_16
X_26537_ _11517_ net1580 _11608_ _11612_ VGND VGND VPWR VPWR _03214_ sky130_fd_sc_hd__a31o_1
XFILLER_0_28_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_278 _13248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_289 _13309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_184_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0__10137_ _10137_ VGND VGND VPWR VPWR clknet_0__10137_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_95_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29256_ _13148_ VGND VGND VPWR VPWR _04397_ sky130_fd_sc_hd__clkbuf_1
X_17270_ _14189_ net2664 _04887_ VGND VGND VPWR VPWR _04896_ sky130_fd_sc_hd__mux2_1
X_26468_ net1929 _11573_ _11590_ _11570_ VGND VGND VPWR VPWR _03167_ sky130_fd_sc_hd__o211a_1
XFILLER_0_3_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16221_ _13247_ VGND VGND VPWR VPWR _14466_ sky130_fd_sc_hd__buf_4
X_28207_ _12571_ VGND VGND VPWR VPWR _03925_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_180_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25419_ _10965_ VGND VGND VPWR VPWR _02743_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26399_ _11143_ VGND VGND VPWR VPWR _11542_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_180_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29187_ _09259_ net2324 _13103_ VGND VGND VPWR VPWR _13111_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16152_ net1919 _13278_ _14384_ VGND VGND VPWR VPWR _14419_ sky130_fd_sc_hd__mux2_1
Xclkload209 clknet_leaf_203_clk VGND VGND VPWR VPWR clkload209/Y sky130_fd_sc_hd__clkinv_1
XFILLER_0_180_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28138_ _12443_ net2926 _12528_ VGND VGND VPWR VPWR _12535_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15103_ _13488_ _13492_ VGND VGND VPWR VPWR _13648_ sky130_fd_sc_hd__nor2_1
XFILLER_0_180_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_185_4925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16083_ _14382_ VGND VGND VPWR VPWR _01981_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_185_4936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28069_ _12498_ VGND VGND VPWR VPWR _03860_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_185_4947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15034_ _13483_ VGND VGND VPWR VPWR _13581_ sky130_fd_sc_hd__clkbuf_4
X_19911_ datamem.data_ram\[40\]\[17\] _06648_ _06707_ datamem.data_ram\[47\]\[17\]
+ _07205_ VGND VGND VPWR VPWR _07206_ sky130_fd_sc_hd__o221a_1
X_30100_ net462 _01835_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[11\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_31080_ clknet_leaf_100_clk _02815_ VGND VGND VPWR VPWR datamem.data_ram\[20\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_75_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30031_ net393 _01766_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[13\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_19842_ _06943_ VGND VGND VPWR VPWR _07137_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_88_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19773_ _06681_ _07060_ _07062_ _07067_ VGND VGND VPWR VPWR _07068_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_88_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16985_ net2164 _14468_ _04742_ VGND VGND VPWR VPWR _04745_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_144_3943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_3954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18724_ _06071_ _06074_ _06075_ VGND VGND VPWR VPWR _06076_ sky130_fd_sc_hd__or3b_1
X_15936_ net2568 _13263_ _14297_ VGND VGND VPWR VPWR _14304_ sky130_fd_sc_hd__mux2_1
XFILLER_0_189_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31982_ clknet_leaf_147_clk _03404_ VGND VGND VPWR VPWR datamem.data_ram\[53\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18655_ _05421_ _05424_ _05729_ VGND VGND VPWR VPWR _06011_ sky130_fd_sc_hd__o21a_1
XFILLER_0_64_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30933_ clknet_leaf_264_clk _02668_ VGND VGND VPWR VPWR datamem.data_ram\[40\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15867_ net2155 _13266_ _14258_ VGND VGND VPWR VPWR _14266_ sky130_fd_sc_hd__mux2_1
XFILLER_0_203_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17606_ _05074_ VGND VGND VPWR VPWR _01234_ sky130_fd_sc_hd__clkbuf_1
X_14818_ _13286_ _13288_ VGND VGND VPWR VPWR _13371_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18586_ _05588_ _05726_ _05879_ _05944_ VGND VGND VPWR VPWR _05945_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_47_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30864_ clknet_leaf_260_clk _02599_ VGND VGND VPWR VPWR datamem.data_ram\[43\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_15798_ _14187_ net2621 _14221_ VGND VGND VPWR VPWR _14229_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32603_ clknet_leaf_239_clk _04025_ VGND VGND VPWR VPWR datamem.data_ram\[20\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_24036__565 clknet_1_0__leaf__10245_ VGND VGND VPWR VPWR net691 sky130_fd_sc_hd__inv_2
X_17537_ _13260_ net2622 _05032_ VGND VGND VPWR VPWR _05038_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14749_ _13298_ _13301_ VGND VGND VPWR VPWR _13302_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30795_ clknet_leaf_172_clk _02530_ VGND VGND VPWR VPWR datamem.data_ram\[46\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32534_ clknet_leaf_240_clk _03956_ VGND VGND VPWR VPWR datamem.data_ram\[23\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17468_ _05001_ VGND VGND VPWR VPWR _01307_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22964__673 clknet_1_1__leaf__10081_ VGND VGND VPWR VPWR net799 sky130_fd_sc_hd__inv_2
X_19207_ _06514_ _06515_ VGND VGND VPWR VPWR _06516_ sky130_fd_sc_hd__and2_1
XFILLER_0_156_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16419_ net1893 _14449_ _14572_ VGND VGND VPWR VPWR _14576_ sky130_fd_sc_hd__mux2_1
X_32465_ clknet_leaf_77_clk _03887_ VGND VGND VPWR VPWR datamem.data_ram\[26\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17399_ _14181_ net2834 _04960_ VGND VGND VPWR VPWR _04965_ sky130_fd_sc_hd__mux2_1
X_31416_ clknet_leaf_104_clk _03119_ VGND VGND VPWR VPWR datamem.data_ram\[15\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_19138_ rvcpu.dp.plde.ImmExtE\[16\] rvcpu.dp.plde.PCE\[16\] VGND VGND VPWR VPWR _06455_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_171_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_229_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32396_ clknet_leaf_80_clk _03818_ VGND VGND VPWR VPWR datamem.data_ram\[29\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19069_ rvcpu.dp.plde.ImmExtE\[7\] rvcpu.dp.plde.PCE\[7\] VGND VGND VPWR VPWR _06395_
+ sky130_fd_sc_hd__or2_1
X_31347_ clknet_leaf_19_clk _03050_ VGND VGND VPWR VPWR rvcpu.dp.plde.ALUControlE\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_8_clk clknet_5_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_14_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21100_ datamem.data_ram\[8\]\[7\] _06652_ VGND VGND VPWR VPWR _08389_ sky130_fd_sc_hd__or2_1
X_22080_ rvcpu.dp.plem.MemWriteM _06911_ _09216_ VGND VGND VPWR VPWR _09294_ sky130_fd_sc_hd__and3_1
X_31278_ clknet_leaf_125_clk _02981_ VGND VGND VPWR VPWR datamem.data_ram\[24\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__10126_ clknet_0__10126_ VGND VGND VPWR VPWR clknet_1_0__leaf__10126_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_100_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21031_ datamem.data_ram\[18\]\[31\] datamem.data_ram\[19\]\[31\] _07824_ VGND VGND
+ VPWR VPWR _08320_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30229_ net583 _01964_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[7\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_226_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25770_ _13539_ _08598_ _11165_ VGND VGND VPWR VPWR _11169_ sky130_fd_sc_hd__and3_1
XFILLER_0_97_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21933_ rvcpu.dp.rf.reg_file_arr\[24\]\[29\] rvcpu.dp.rf.reg_file_arr\[25\]\[29\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[29\] rvcpu.dp.rf.reg_file_arr\[27\]\[29\] _08536_
+ _08693_ VGND VGND VPWR VPWR _09166_ sky130_fd_sc_hd__mux4_1
X_24721_ _10568_ VGND VGND VPWR VPWR _02442_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24652_ _07182_ _10042_ _10044_ VGND VGND VPWR VPWR _10530_ sky130_fd_sc_hd__or3_1
XFILLER_0_145_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27440_ _12145_ net2719 _12143_ VGND VGND VPWR VPWR _12146_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21864_ rvcpu.dp.rf.reg_file_arr\[12\]\[25\] rvcpu.dp.rf.reg_file_arr\[13\]\[25\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[25\] rvcpu.dp.rf.reg_file_arr\[15\]\[25\] _08578_
+ _08684_ VGND VGND VPWR VPWR _09101_ sky130_fd_sc_hd__mux4_1
XFILLER_0_49_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20815_ datamem.data_ram\[62\]\[30\] _07859_ _07862_ datamem.data_ram\[60\]\[30\]
+ _08104_ VGND VGND VPWR VPWR _08105_ sky130_fd_sc_hd__o221a_1
X_27371_ _12093_ net3169 _12097_ VGND VGND VPWR VPWR _12104_ sky130_fd_sc_hd__mux2_1
X_24583_ _10492_ VGND VGND VPWR VPWR _02380_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_997 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21795_ rvcpu.dp.rf.reg_file_arr\[0\]\[21\] rvcpu.dp.rf.reg_file_arr\[1\]\[21\] rvcpu.dp.rf.reg_file_arr\[2\]\[21\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[21\] _08566_ _08554_ VGND VGND VPWR VPWR _09036_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_182_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29110_ _13070_ VGND VGND VPWR VPWR _04329_ sky130_fd_sc_hd__clkbuf_1
X_26322_ _10043_ VGND VGND VPWR VPWR _11494_ sky130_fd_sc_hd__buf_2
X_20746_ _08030_ _08035_ VGND VGND VPWR VPWR _08036_ sky130_fd_sc_hd__or2_1
XFILLER_0_175_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_150_4103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_189_5025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29041_ _10060_ _13031_ VGND VGND VPWR VPWR _13034_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_189_5036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26253_ net116 _11457_ _11459_ net1300 VGND VGND VPWR VPWR _03083_ sky130_fd_sc_hd__a2bb2o_1
X_20677_ datamem.data_ram\[42\]\[5\] _06989_ _06921_ datamem.data_ram\[45\]\[5\] VGND
+ VGND VPWR VPWR _07968_ sky130_fd_sc_hd__a22o_1
XFILLER_0_190_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25204_ _10814_ net2912 net56 VGND VGND VPWR VPWR _10841_ sky130_fd_sc_hd__mux2_1
X_22416_ _09511_ _09575_ VGND VGND VPWR VPWR _09576_ sky130_fd_sc_hd__or2_1
X_26184_ _08513_ _11413_ VGND VGND VPWR VPWR _11429_ sky130_fd_sc_hd__and2_1
X_23396_ _09322_ net2812 _10143_ VGND VGND VPWR VPWR _10149_ sky130_fd_sc_hd__mux2_1
X_25135_ _10799_ VGND VGND VPWR VPWR _02625_ sky130_fd_sc_hd__clkbuf_1
X_22347_ _09411_ VGND VGND VPWR VPWR _09510_ sky130_fd_sc_hd__buf_2
XFILLER_0_131_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_227_5932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23437__88 clknet_1_1__leaf__10155_ VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_227_5943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23271__916 clknet_1_0__leaf__10129_ VGND VGND VPWR VPWR net1042 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_227_5954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25066_ _10762_ net4167 _10752_ VGND VGND VPWR VPWR _10763_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29943_ net313 _01678_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[15\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_148_4043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22278_ _09381_ VGND VGND VPWR VPWR _09443_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_103_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_148_4054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23883__444 clknet_1_1__leaf__10221_ VGND VGND VPWR VPWR net570 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_180_4811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold180 datamem.data_ram\[44\]\[6\] VGND VGND VPWR VPWR net1330 sky130_fd_sc_hd__dlygate4sd3_1
X_21229_ datamem.data_ram\[52\]\[6\] datamem.data_ram\[53\]\[6\] datamem.data_ram\[52\]\[30\]
+ datamem.data_ram\[52\]\[22\] VGND VGND VPWR VPWR _08492_ sky130_fd_sc_hd__or4_2
Xhold191 datamem.data_ram\[42\]\[5\] VGND VGND VPWR VPWR net1341 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_180_4822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29874_ net252 _01609_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[17\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_229_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28825_ _12915_ VGND VGND VPWR VPWR _04199_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_6_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_171_Left_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_219_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_189_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16770_ net2717 _14457_ _04623_ VGND VGND VPWR VPWR _04631_ sky130_fd_sc_hd__mux2_1
X_28756_ _12878_ VGND VGND VPWR VPWR _04167_ sky130_fd_sc_hd__clkbuf_1
X_25968_ net30 _11289_ VGND VGND VPWR VPWR _11307_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_107_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15721_ _13262_ VGND VGND VPWR VPWR _14185_ sky130_fd_sc_hd__buf_4
X_27707_ _12147_ net4179 _12289_ VGND VGND VPWR VPWR _12292_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24919_ _10677_ VGND VGND VPWR VPWR _02531_ sky130_fd_sc_hd__clkbuf_1
X_28687_ _12734_ net2765 net42 VGND VGND VPWR VPWR _12842_ sky130_fd_sc_hd__mux2_1
X_25899_ _13706_ _11256_ _11258_ _11267_ VGND VGND VPWR VPWR _02921_ sky130_fd_sc_hd__o211a_1
XFILLER_0_217_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_178_4762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18440_ _05373_ _05663_ _05802_ VGND VGND VPWR VPWR _05803_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_17_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_4773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27638_ _12254_ VGND VGND VPWR VPWR _03673_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_17_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15652_ _14138_ VGND VGND VPWR VPWR _02184_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14603_ rvcpu.dp.plmw.ALUResultW\[29\] rvcpu.dp.plmw.ReadDataW\[29\] rvcpu.dp.plmw.PCPlus4W\[29\]
+ rvcpu.dp.plmw.lAuiPCW\[29\] _13168_ _13170_ VGND VGND VPWR VPWR _13186_ sky130_fd_sc_hd__mux4_2
X_18371_ _05283_ _05728_ _05730_ _05281_ _05735_ VGND VGND VPWR VPWR _05736_ sky130_fd_sc_hd__a221o_1
X_15583_ net3408 _13201_ _14092_ VGND VGND VPWR VPWR _14099_ sky130_fd_sc_hd__mux2_1
X_27569_ _12085_ net3012 net82 VGND VGND VPWR VPWR _12218_ sky130_fd_sc_hd__mux2_1
XFILLER_0_185_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17322_ _04901_ VGND VGND VPWR VPWR _04924_ sky130_fd_sc_hd__clkbuf_4
X_29308_ clknet_leaf_0_clk _01043_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD1E\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_945 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30580_ clknet_leaf_178_clk _02315_ VGND VGND VPWR VPWR datamem.data_ram\[54\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_180_Left_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_682 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17253_ _04864_ VGND VGND VPWR VPWR _04887_ sky130_fd_sc_hd__clkbuf_4
X_29239_ _13139_ VGND VGND VPWR VPWR _04389_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_3780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_3791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16204_ _14454_ VGND VGND VPWR VPWR _01932_ sky130_fd_sc_hd__clkbuf_1
X_32250_ clknet_leaf_87_clk _03672_ VGND VGND VPWR VPWR datamem.data_ram\[34\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17184_ _04850_ VGND VGND VPWR VPWR _01448_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31201_ clknet_leaf_28_clk _02904_ VGND VGND VPWR VPWR rvcpu.dp.plfd.PCPlus4D\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_133_3677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_133_3688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16135_ _14410_ VGND VGND VPWR VPWR _01957_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_133_3699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32181_ clknet_leaf_166_clk _03603_ VGND VGND VPWR VPWR datamem.data_ram\[37\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31132_ clknet_leaf_125_clk _02867_ VGND VGND VPWR VPWR datamem.data_ram\[25\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_224_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16066_ net2261 _13251_ _14371_ VGND VGND VPWR VPWR _14374_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15017_ _13397_ _13390_ VGND VGND VPWR VPWR _13565_ sky130_fd_sc_hd__nand2_2
X_23133__809 clknet_1_1__leaf__10106_ VGND VGND VPWR VPWR net935 sky130_fd_sc_hd__inv_2
XFILLER_0_110_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31063_ clknet_leaf_255_clk _02798_ VGND VGND VPWR VPWR datamem.data_ram\[8\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2509 rvcpu.dp.rf.reg_file_arr\[26\]\[5\] VGND VGND VPWR VPWR net3659 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_36_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19825_ rvcpu.dp.plem.ALUResultM\[1\] _06588_ VGND VGND VPWR VPWR _07120_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_36_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30014_ net376 _01749_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[13\]\[1\] sky130_fd_sc_hd__dfxtp_1
Xhold1808 datamem.data_ram\[0\]\[28\] VGND VGND VPWR VPWR net2958 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1819 rvcpu.dp.rf.reg_file_arr\[20\]\[29\] VGND VGND VPWR VPWR net2969 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19756_ datamem.data_ram\[62\]\[25\] _06719_ _06810_ _07050_ VGND VGND VPWR VPWR
+ _07051_ sky130_fd_sc_hd__o211a_1
X_16968_ net2296 _14451_ _04731_ VGND VGND VPWR VPWR _04736_ sky130_fd_sc_hd__mux2_1
X_18707_ _05697_ _05749_ _05906_ _05889_ VGND VGND VPWR VPWR _06060_ sky130_fd_sc_hd__a31o_1
X_15919_ net3590 _13238_ _14286_ VGND VGND VPWR VPWR _14295_ sky130_fd_sc_hd__mux2_1
X_19687_ datamem.data_ram\[60\]\[0\] _06977_ _06979_ _06982_ VGND VGND VPWR VPWR _06983_
+ sky130_fd_sc_hd__a211o_1
X_31965_ clknet_leaf_120_clk _03387_ VGND VGND VPWR VPWR datamem.data_ram\[28\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_16899_ _04699_ VGND VGND VPWR VPWR _01590_ sky130_fd_sc_hd__clkbuf_1
X_18638_ _05993_ _05654_ _05994_ VGND VGND VPWR VPWR _05995_ sky130_fd_sc_hd__or3_1
X_30916_ clknet_leaf_281_clk _02651_ VGND VGND VPWR VPWR datamem.data_ram\[41\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31896_ _04426_ net120 VGND VGND VPWR VPWR datamem.rd_data_mem\[1\] sky130_fd_sc_hd__dlxtn_1
XFILLER_0_188_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_77 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18569_ _05912_ _05913_ _05924_ _05928_ VGND VGND VPWR VPWR _05929_ sky130_fd_sc_hd__o211a_1
X_30847_ clknet_leaf_203_clk _02582_ VGND VGND VPWR VPWR datamem.data_ram\[43\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20600_ datamem.data_ram\[6\]\[13\] _06682_ _06671_ datamem.data_ram\[7\]\[13\] VGND
+ VGND VPWR VPWR _07891_ sky130_fd_sc_hd__o22a_1
XFILLER_0_129_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21580_ _08627_ _08827_ _08829_ _08831_ VGND VGND VPWR VPWR _08832_ sky130_fd_sc_hd__o2bb2a_1
X_30778_ clknet_leaf_221_clk _02513_ VGND VGND VPWR VPWR datamem.data_ram\[46\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32517_ clknet_leaf_78_clk _03939_ VGND VGND VPWR VPWR datamem.data_ram\[24\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20531_ _07821_ VGND VGND VPWR VPWR _07822_ sky130_fd_sc_hd__buf_8
XFILLER_0_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20462_ datamem.data_ram\[21\]\[20\] _06661_ _06704_ datamem.data_ram\[23\]\[20\]
+ VGND VGND VPWR VPWR _07754_ sky130_fd_sc_hd__o22a_1
X_32448_ clknet_leaf_4_clk _03870_ VGND VGND VPWR VPWR datamem.data_ram\[27\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_330 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22201_ _09373_ VGND VGND VPWR VPWR _01117_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_160_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32379_ clknet_leaf_164_clk _03801_ VGND VGND VPWR VPWR datamem.data_ram\[2\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_20393_ datamem.data_ram\[31\]\[28\] _06725_ _06655_ datamem.data_ram\[25\]\[28\]
+ _07684_ VGND VGND VPWR VPWR _07685_ sky130_fd_sc_hd__o221a_1
XFILLER_0_43_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22132_ _09335_ VGND VGND VPWR VPWR _01086_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_203_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26940_ _11849_ net1542 _11841_ _11850_ VGND VGND VPWR VPWR _03379_ sky130_fd_sc_hd__a31o_1
X_22063_ rvcpu.dp.plem.WriteDataM\[4\] _09264_ _09265_ rvcpu.dp.plem.WriteDataM\[12\]
+ VGND VGND VPWR VPWR _09281_ sky130_fd_sc_hd__a22o_4
XFILLER_0_11_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__10109_ clknet_0__10109_ VGND VGND VPWR VPWR clknet_1_0__leaf__10109_
+ sky130_fd_sc_hd__clkbuf_16
X_21014_ datamem.data_ram\[60\]\[31\] datamem.data_ram\[61\]\[31\] _07912_ VGND VGND
+ VPWR VPWR _08303_ sky130_fd_sc_hd__mux2_1
XFILLER_0_227_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26871_ _11689_ _11798_ VGND VGND VPWR VPWR _11806_ sky130_fd_sc_hd__and2_1
XFILLER_0_226_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_250_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_250_clk
+ sky130_fd_sc_hd__clkbuf_8
X_28610_ _12696_ net3313 _12796_ VGND VGND VPWR VPWR _12801_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25822_ rvcpu.dp.pcreg.q\[20\] _11200_ rvcpu.dp.pcreg.q\[21\] VGND VGND VPWR VPWR
+ _11209_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_227_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29590_ net944 _01325_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[26\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_28541_ _12762_ net3154 _12752_ VGND VGND VPWR VPWR _12763_ sky130_fd_sc_hd__mux2_1
XFILLER_0_214_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25753_ _11153_ _11154_ _11156_ _11147_ VGND VGND VPWR VPWR _02886_ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_195_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24704_ _10559_ VGND VGND VPWR VPWR _02434_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28472_ _12718_ VGND VGND VPWR VPWR _04043_ sky130_fd_sc_hd__clkbuf_1
X_21916_ _08531_ _09149_ _08806_ VGND VGND VPWR VPWR _09150_ sky130_fd_sc_hd__o21a_1
X_25684_ _11078_ _11113_ VGND VGND VPWR VPWR _11114_ sky130_fd_sc_hd__and2_1
X_22896_ _09510_ _10024_ _10026_ _10030_ _08589_ VGND VGND VPWR VPWR _10031_ sky130_fd_sc_hd__a311o_1
XFILLER_0_168_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27423_ _09247_ VGND VGND VPWR VPWR _12134_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_139_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24635_ _10520_ _10347_ _10501_ VGND VGND VPWR VPWR _10521_ sky130_fd_sc_hd__a21oi_4
X_21847_ rvcpu.dp.rf.reg_file_arr\[8\]\[24\] rvcpu.dp.rf.reg_file_arr\[10\]\[24\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[24\] rvcpu.dp.rf.reg_file_arr\[11\]\[24\] _08635_
+ _08561_ VGND VGND VPWR VPWR _09085_ sky130_fd_sc_hd__mux4_1
X_24132__637 clknet_1_1__leaf__10261_ VGND VGND VPWR VPWR net763 sky130_fd_sc_hd__inv_2
XFILLER_0_66_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_468 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_216_5677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_216_5688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24566_ _10483_ VGND VGND VPWR VPWR _02372_ sky130_fd_sc_hd__clkbuf_1
X_27354_ _12094_ VGND VGND VPWR VPWR _03549_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_182_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21778_ _08817_ _09017_ _09019_ _08700_ VGND VGND VPWR VPWR _09020_ sky130_fd_sc_hd__a211o_1
XFILLER_0_33_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26305_ _11485_ VGND VGND VPWR VPWR _03109_ sky130_fd_sc_hd__clkbuf_1
X_20729_ datamem.data_ram\[28\]\[6\] datamem.data_ram\[29\]\[6\] _07829_ VGND VGND
+ VPWR VPWR _08019_ sky130_fd_sc_hd__mux2_1
X_23517_ _09248_ net4158 _10162_ VGND VGND VPWR VPWR _10167_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27285_ _12036_ net1454 _12053_ _12055_ VGND VGND VPWR VPWR _03519_ sky130_fd_sc_hd__a31o_1
X_24497_ _09223_ VGND VGND VPWR VPWR _10439_ sky130_fd_sc_hd__buf_2
XFILLER_0_80_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29024_ _12741_ net3961 net66 VGND VGND VPWR VPWR _13024_ sky130_fd_sc_hd__mux2_1
X_26236_ _11379_ _03042_ _11454_ VGND VGND VPWR VPWR _03069_ sky130_fd_sc_hd__a21o_1
XFILLER_0_110_1286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26167_ _11420_ VGND VGND VPWR VPWR _03036_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25118_ _10790_ VGND VGND VPWR VPWR _02617_ sky130_fd_sc_hd__clkbuf_1
X_26098_ net1623 _11372_ VGND VGND VPWR VPWR _11384_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_72_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25049_ _09223_ VGND VGND VPWR VPWR _10751_ sky130_fd_sc_hd__buf_2
X_17940_ rvcpu.dp.plem.ALUResultM\[15\] _05272_ VGND VGND VPWR VPWR _05312_ sky130_fd_sc_hd__and2_1
X_29926_ net296 _01661_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[16\]\[17\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_167_4496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_109_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17871_ _05241_ rvcpu.dp.plem.RdM\[0\] _05242_ rvcpu.dp.plde.Rs1E\[3\] _05243_ VGND
+ VGND VPWR VPWR _05244_ sky130_fd_sc_hd__o221a_1
X_29857_ net235 _01592_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[18\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19610_ _06810_ _06903_ _06905_ VGND VGND VPWR VPWR _06906_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_241_clk clknet_5_17__leaf_clk VGND VGND VPWR VPWR clknet_leaf_241_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_205_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28808_ _12906_ VGND VGND VPWR VPWR _04191_ sky130_fd_sc_hd__clkbuf_1
X_16822_ _04658_ VGND VGND VPWR VPWR _01626_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_206_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_105_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29788_ net1134 _01523_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[20\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_31_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19541_ _06807_ VGND VGND VPWR VPWR _06837_ sky130_fd_sc_hd__buf_6
XFILLER_0_45_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28739_ _12869_ VGND VGND VPWR VPWR _04159_ sky130_fd_sc_hd__clkbuf_1
X_16753_ net3882 _14440_ _04612_ VGND VGND VPWR VPWR _04622_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_219_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_220_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15704_ _14172_ net2933 _14173_ VGND VGND VPWR VPWR _14174_ sky130_fd_sc_hd__mux2_1
X_31750_ clknet_leaf_58_clk _03204_ VGND VGND VPWR VPWR datamem.data_ram\[45\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_19472_ _06722_ VGND VGND VPWR VPWR _06768_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_88_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16684_ _04585_ VGND VGND VPWR VPWR _01699_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_216_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_213_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18423_ _00003_ _05786_ _05395_ VGND VGND VPWR VPWR _05787_ sky130_fd_sc_hd__a21o_1
X_30701_ clknet_leaf_217_clk _02436_ VGND VGND VPWR VPWR datamem.data_ram\[49\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15635_ net2949 _13278_ _14091_ VGND VGND VPWR VPWR _14126_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31681_ clknet_leaf_13_clk net1265 VGND VGND VPWR VPWR rvcpu.dp.plmw.ALUResultW\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_139_3820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_186_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_139_3831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_139_3842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18354_ _05380_ _05668_ _05662_ VGND VGND VPWR VPWR _05719_ sky130_fd_sc_hd__or3_2
XFILLER_0_29_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30632_ clknet_leaf_220_clk _02367_ VGND VGND VPWR VPWR datamem.data_ram\[51\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_15566_ _14088_ VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_29_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17305_ _04915_ VGND VGND VPWR VPWR _01392_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_185_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_3728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_185_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18285_ _05283_ _05649_ VGND VGND VPWR VPWR _05650_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_3739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30563_ clknet_leaf_195_clk _02298_ VGND VGND VPWR VPWR datamem.data_ram\[54\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_15497_ _13517_ _13337_ _13853_ VGND VGND VPWR VPWR _14025_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32302_ clknet_leaf_88_clk _03724_ VGND VGND VPWR VPWR datamem.data_ram\[32\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17236_ _04878_ VGND VGND VPWR VPWR _01424_ sky130_fd_sc_hd__clkbuf_1
X_23751__341 clknet_1_1__leaf__10200_ VGND VGND VPWR VPWR net467 sky130_fd_sc_hd__inv_2
X_30494_ clknet_leaf_141_clk _02229_ VGND VGND VPWR VPWR datamem.data_ram\[57\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_32233_ clknet_leaf_242_clk _03655_ VGND VGND VPWR VPWR datamem.data_ram\[35\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17167_ _14154_ net4133 _04840_ VGND VGND VPWR VPWR _04842_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold905 rvcpu.dp.rf.reg_file_arr\[3\]\[20\] VGND VGND VPWR VPWR net2055 sky130_fd_sc_hd__dlygate4sd3_1
Xhold916 rvcpu.dp.rf.reg_file_arr\[19\]\[21\] VGND VGND VPWR VPWR net2066 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_49_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold927 rvcpu.dp.rf.reg_file_arr\[17\]\[20\] VGND VGND VPWR VPWR net2077 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16118_ _14401_ VGND VGND VPWR VPWR _01965_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold938 rvcpu.dp.rf.reg_file_arr\[11\]\[5\] VGND VGND VPWR VPWR net2088 sky130_fd_sc_hd__dlygate4sd3_1
X_32164_ clknet_leaf_256_clk _03586_ VGND VGND VPWR VPWR datamem.data_ram\[38\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_17098_ _04805_ VGND VGND VPWR VPWR _01489_ sky130_fd_sc_hd__clkbuf_1
Xhold949 rvcpu.dp.rf.reg_file_arr\[12\]\[5\] VGND VGND VPWR VPWR net2099 sky130_fd_sc_hd__dlygate4sd3_1
X_23416__69 clknet_1_0__leaf__10153_ VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__inv_2
X_31115_ clknet_leaf_61_clk _02850_ VGND VGND VPWR VPWR datamem.data_ram\[43\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3007 datamem.data_ram\[56\]\[17\] VGND VGND VPWR VPWR net4157 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3018 datamem.data_ram\[40\]\[16\] VGND VGND VPWR VPWR net4168 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16049_ net3168 _13226_ _14360_ VGND VGND VPWR VPWR _14365_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3029 datamem.data_ram\[33\]\[10\] VGND VGND VPWR VPWR net4179 sky130_fd_sc_hd__dlygate4sd3_1
X_32095_ clknet_leaf_209_clk _03517_ VGND VGND VPWR VPWR datamem.data_ram\[8\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2306 datamem.data_ram\[54\]\[25\] VGND VGND VPWR VPWR net3456 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31046_ clknet_leaf_212_clk _02781_ VGND VGND VPWR VPWR datamem.data_ram\[9\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2317 rvcpu.dp.rf.reg_file_arr\[26\]\[21\] VGND VGND VPWR VPWR net3467 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2328 datamem.data_ram\[20\]\[22\] VGND VGND VPWR VPWR net3478 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2339 rvcpu.dp.rf.reg_file_arr\[7\]\[31\] VGND VGND VPWR VPWR net3489 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1605 rvcpu.dp.rf.reg_file_arr\[22\]\[7\] VGND VGND VPWR VPWR net2755 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_232_clk clknet_5_20__leaf_clk VGND VGND VPWR VPWR clknet_leaf_232_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold1616 rvcpu.dp.rf.reg_file_arr\[18\]\[12\] VGND VGND VPWR VPWR net2766 sky130_fd_sc_hd__dlygate4sd3_1
X_19808_ datamem.data_ram\[4\]\[9\] _06766_ _06699_ datamem.data_ram\[1\]\[9\] VGND
+ VGND VPWR VPWR _07103_ sky130_fd_sc_hd__o22a_1
Xhold1627 datamem.data_ram\[28\]\[18\] VGND VGND VPWR VPWR net2777 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1638 datamem.data_ram\[38\]\[19\] VGND VGND VPWR VPWR net2788 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1649 rvcpu.dp.rf.reg_file_arr\[8\]\[2\] VGND VGND VPWR VPWR net2799 sky130_fd_sc_hd__dlygate4sd3_1
X_19739_ datamem.data_ram\[6\]\[25\] _07028_ _07029_ _07033_ VGND VGND VPWR VPWR _07034_
+ sky130_fd_sc_hd__o211a_1
X_22750_ rvcpu.dp.rf.reg_file_arr\[0\]\[23\] rvcpu.dp.rf.reg_file_arr\[1\]\[23\] rvcpu.dp.rf.reg_file_arr\[2\]\[23\]
+ rvcpu.dp.rf.reg_file_arr\[3\]\[23\] _09714_ _09383_ VGND VGND VPWR VPWR _09893_
+ sky130_fd_sc_hd__mux4_1
X_31948_ clknet_leaf_117_clk _03370_ VGND VGND VPWR VPWR datamem.data_ram\[32\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_223_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21701_ _08663_ _08944_ _08946_ _08558_ VGND VGND VPWR VPWR _08947_ sky130_fd_sc_hd__o211a_1
X_22681_ rvcpu.dp.rf.reg_file_arr\[12\]\[19\] rvcpu.dp.rf.reg_file_arr\[13\]\[19\]
+ rvcpu.dp.rf.reg_file_arr\[14\]\[19\] rvcpu.dp.rf.reg_file_arr\[15\]\[19\] _09462_
+ _09721_ VGND VGND VPWR VPWR _09828_ sky130_fd_sc_hd__mux4_1
X_31879_ clknet_leaf_124_clk _03333_ VGND VGND VPWR VPWR datamem.data_ram\[57\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24420_ _10391_ VGND VGND VPWR VPWR _02318_ sky130_fd_sc_hd__clkbuf_1
X_21632_ _08881_ VGND VGND VPWR VPWR _01040_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_192_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24351_ _09282_ net2594 _10348_ VGND VGND VPWR VPWR _10353_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_1338 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21563_ _08682_ _08812_ _08815_ VGND VGND VPWR VPWR _08816_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_211_5552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27070_ _11829_ _11924_ VGND VGND VPWR VPWR _11928_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_211_5563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20514_ datamem.data_ram\[58\]\[21\] _06613_ _07791_ datamem.data_ram\[63\]\[21\]
+ _07804_ VGND VGND VPWR VPWR _07805_ sky130_fd_sc_hd__o221a_1
XFILLER_0_118_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24282_ _09256_ net3199 _10307_ VGND VGND VPWR VPWR _10314_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21494_ _08627_ _08744_ _08746_ _08749_ VGND VGND VPWR VPWR _08750_ sky130_fd_sc_hd__o2bb2a_1
X_23949__503 clknet_1_1__leaf__10228_ VGND VGND VPWR VPWR net629 sky130_fd_sc_hd__inv_2
X_23001__706 clknet_1_1__leaf__10085_ VGND VGND VPWR VPWR net832 sky130_fd_sc_hd__inv_2
XFILLER_0_172_493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26021_ net25 _11152_ VGND VGND VPWR VPWR _11336_ sky130_fd_sc_hd__or2_1
X_20445_ _07714_ _07736_ VGND VGND VPWR VPWR _07737_ sky130_fd_sc_hd__nor2_4
XFILLER_0_160_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20376_ _06714_ _07662_ _07667_ VGND VGND VPWR VPWR _07668_ sky130_fd_sc_hd__or3_2
XFILLER_0_63_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_189_Right_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22115_ _09323_ VGND VGND VPWR VPWR _01081_ sky130_fd_sc_hd__clkbuf_1
X_27972_ _12441_ net2302 _12431_ VGND VGND VPWR VPWR _12442_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23095_ clknet_1_0__leaf__10087_ VGND VGND VPWR VPWR _10103_ sky130_fd_sc_hd__buf_1
X_29711_ net1057 _01446_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[22\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26923_ _07791_ _10402_ _11839_ VGND VGND VPWR VPWR _11840_ sky130_fd_sc_hd__or3_1
X_22046_ _09264_ _09265_ VGND VGND VPWR VPWR _09268_ sky130_fd_sc_hd__nor2_8
XFILLER_0_227_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_223_clk clknet_5_21__leaf_clk VGND VGND VPWR VPWR clknet_leaf_223_clk
+ sky130_fd_sc_hd__clkbuf_8
X_29642_ net988 _01377_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[24\]\[5\] sky130_fd_sc_hd__dfxtp_1
Xhold2840 datamem.data_ram\[5\]\[15\] VGND VGND VPWR VPWR net3990 sky130_fd_sc_hd__dlygate4sd3_1
X_26854_ _11752_ VGND VGND VPWR VPWR _11795_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_162_4382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2851 datamem.data_ram\[23\]\[23\] VGND VGND VPWR VPWR net4001 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_162_4393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2862 datamem.data_ram\[49\]\[27\] VGND VGND VPWR VPWR net4012 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2873 datamem.data_ram\[10\]\[28\] VGND VGND VPWR VPWR net4023 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2884 rvcpu.dp.rf.reg_file_arr\[26\]\[30\] VGND VGND VPWR VPWR net4034 sky130_fd_sc_hd__dlygate4sd3_1
X_25805_ _11194_ _11195_ _11157_ VGND VGND VPWR VPWR _11196_ sky130_fd_sc_hd__a21o_1
XFILLER_0_138_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2895 datamem.data_ram\[46\]\[23\] VGND VGND VPWR VPWR net4045 sky130_fd_sc_hd__dlygate4sd3_1
X_29573_ net927 _01308_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[26\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_23921__477 clknet_1_1__leaf__10226_ VGND VGND VPWR VPWR net603 sky130_fd_sc_hd__inv_2
X_26785_ _11684_ _11749_ VGND VGND VPWR VPWR _11755_ sky130_fd_sc_hd__and2_1
XFILLER_0_216_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_218_5717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28524_ _09223_ VGND VGND VPWR VPWR _12751_ sky130_fd_sc_hd__buf_2
XFILLER_0_138_1175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_218_5728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25736_ _08598_ VGND VGND VPWR VPWR _11142_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_218_5739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22948_ rvcpu.dp.plem.WriteDataM\[7\] VGND VGND VPWR VPWR _10075_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23620__238 clknet_1_1__leaf__10180_ VGND VGND VPWR VPWR net364 sky130_fd_sc_hd__inv_2
XFILLER_0_70_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28455_ _12709_ VGND VGND VPWR VPWR _04035_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_65_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25667_ _11086_ _11098_ VGND VGND VPWR VPWR _11102_ sky130_fd_sc_hd__and2_1
XFILLER_0_35_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22879_ rvcpu.dp.rf.reg_file_arr\[4\]\[30\] rvcpu.dp.rf.reg_file_arr\[5\]\[30\] rvcpu.dp.rf.reg_file_arr\[6\]\[30\]
+ rvcpu.dp.rf.reg_file_arr\[7\]\[30\] _09416_ _09418_ VGND VGND VPWR VPWR _10015_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_171_4607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15420_ _13504_ _13949_ _13951_ _13319_ _13539_ VGND VGND VPWR VPWR _13952_ sky130_fd_sc_hd__a221o_1
X_27406_ _12093_ net2125 _12116_ VGND VGND VPWR VPWR _12123_ sky130_fd_sc_hd__mux2_1
X_24618_ _10439_ net3853 _10511_ VGND VGND VPWR VPWR _10512_ sky130_fd_sc_hd__mux2_1
X_28386_ _12178_ _12612_ _12668_ VGND VGND VPWR VPWR _12669_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_109_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25598_ _11057_ net1428 _11053_ _11062_ VGND VGND VPWR VPWR _02825_ sky130_fd_sc_hd__a31o_1
XFILLER_0_167_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15351_ _13608_ _13690_ _13878_ _13886_ VGND VGND VPWR VPWR _13887_ sky130_fd_sc_hd__a211o_1
XFILLER_0_26_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27337_ _09305_ VGND VGND VPWR VPWR _12083_ sky130_fd_sc_hd__buf_2
XFILLER_0_164_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24549_ _09313_ VGND VGND VPWR VPWR _10472_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_80_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23277__922 clknet_1_1__leaf__10129_ VGND VGND VPWR VPWR net1048 sky130_fd_sc_hd__inv_2
X_18070_ _05437_ _05323_ VGND VGND VPWR VPWR _05438_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_108_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15282_ _13638_ _13815_ _13820_ VGND VGND VPWR VPWR _13821_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_163_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27268_ _12045_ VGND VGND VPWR VPWR _03512_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29007_ _12995_ net1663 _13009_ _13014_ VGND VGND VPWR VPWR _04282_ sky130_fd_sc_hd__a31o_1
X_17021_ _04764_ VGND VGND VPWR VPWR _01525_ sky130_fd_sc_hd__clkbuf_1
X_26219_ _11447_ VGND VGND VPWR VPWR _03061_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_3614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_130_3625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27199_ _12005_ net1418 _12007_ _12009_ VGND VGND VPWR VPWR _03479_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_169_4547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_169_4558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_156_Right_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18972_ _05630_ _05631_ _05640_ _05305_ VGND VGND VPWR VPWR _06308_ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_91_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17923_ rvcpu.dp.plde.RD1E\[29\] _05292_ _05295_ VGND VGND VPWR VPWR _05296_ sky130_fd_sc_hd__o21a_1
XFILLER_0_147_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29909_ net279 _01644_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[16\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_128_3565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_214_clk clknet_5_20__leaf_clk VGND VGND VPWR VPWR clknet_leaf_214_clk
+ sky130_fd_sc_hd__clkbuf_8
X_32920_ clknet_leaf_152_clk _04342_ VGND VGND VPWR VPWR datamem.data_ram\[0\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_23781__367 clknet_1_0__leaf__10204_ VGND VGND VPWR VPWR net493 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_128_3576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17854_ rvcpu.dp.plem.ALUResultM\[9\] _05230_ _05176_ VGND VGND VPWR VPWR _05231_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_206_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16805_ net2236 _14424_ _04648_ VGND VGND VPWR VPWR _04650_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24000__534 clknet_1_0__leaf__10240_ VGND VGND VPWR VPWR net660 sky130_fd_sc_hd__inv_2
X_32851_ clknet_leaf_213_clk _04273_ VGND VGND VPWR VPWR datamem.data_ram\[11\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_17785_ _13274_ _05154_ _05161_ net114 VGND VGND VPWR VPWR _05182_ sky130_fd_sc_hd__a31o_1
XFILLER_0_227_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14997_ _13303_ _13322_ VGND VGND VPWR VPWR _13545_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_221_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_50_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31802_ clknet_leaf_59_clk _03256_ VGND VGND VPWR VPWR datamem.data_ram\[46\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_19524_ _06644_ VGND VGND VPWR VPWR _06820_ sky130_fd_sc_hd__buf_6
X_16736_ _04613_ VGND VGND VPWR VPWR _01675_ sky130_fd_sc_hd__clkbuf_1
X_32782_ clknet_leaf_91_clk _04204_ VGND VGND VPWR VPWR datamem.data_ram\[14\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_186_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19455_ _06750_ VGND VGND VPWR VPWR _06751_ sky130_fd_sc_hd__buf_8
X_31733_ net182 _03191_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[9\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16667_ _14127_ net4273 _04576_ VGND VGND VPWR VPWR _04577_ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23595__215 clknet_1_0__leaf__10178_ VGND VGND VPWR VPWR net341 sky130_fd_sc_hd__inv_2
XFILLER_0_186_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18406_ _05376_ _05382_ _05769_ VGND VGND VPWR VPWR _05770_ sky130_fd_sc_hd__mux2_1
X_15618_ _14117_ VGND VGND VPWR VPWR _02197_ sky130_fd_sc_hd__clkbuf_1
X_31664_ clknet_leaf_71_clk net1266 VGND VGND VPWR VPWR rvcpu.dp.plmw.ALUResultW\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_19386_ _06627_ VGND VGND VPWR VPWR _06682_ sky130_fd_sc_hd__buf_8
XFILLER_0_9_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16598_ _04539_ VGND VGND VPWR VPWR _04540_ sky130_fd_sc_hd__buf_4
XFILLER_0_57_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18337_ _05590_ _05660_ VGND VGND VPWR VPWR _05702_ sky130_fd_sc_hd__nor2_4
X_30615_ clknet_leaf_147_clk _02350_ VGND VGND VPWR VPWR datamem.data_ram\[52\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15549_ _13762_ _13878_ _14073_ _13572_ VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__o22a_1
X_23675__272 clknet_1_1__leaf__10193_ VGND VGND VPWR VPWR net398 sky130_fd_sc_hd__inv_2
XFILLER_0_5_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31595_ clknet_leaf_48_clk net1243 VGND VGND VPWR VPWR rvcpu.dp.plmw.PCPlus4W\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30546_ clknet_leaf_139_clk _02281_ VGND VGND VPWR VPWR datamem.data_ram\[55\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18268_ rvcpu.dp.plde.RD1E\[24\] _05291_ _05532_ VGND VGND VPWR VPWR _05633_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_114_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17219_ _04869_ VGND VGND VPWR VPWR _01432_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18199_ _05291_ VGND VGND VPWR VPWR _05564_ sky130_fd_sc_hd__clkbuf_4
X_30477_ net155 _02212_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[19\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_694 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold702 rvcpu.dp.plfd.PCD\[10\] VGND VGND VPWR VPWR net1852 sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 rvcpu.dp.plfd.PCD\[0\] VGND VGND VPWR VPWR net1863 sky130_fd_sc_hd__dlygate4sd3_1
X_20230_ datamem.data_ram\[3\]\[3\] _06961_ _06955_ datamem.data_ram\[4\]\[3\] VGND
+ VGND VPWR VPWR _07523_ sky130_fd_sc_hd__a22o_1
XFILLER_0_163_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32216_ clknet_leaf_276_clk _03638_ VGND VGND VPWR VPWR datamem.data_ram\[36\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold724 rvcpu.dp.rf.reg_file_arr\[18\]\[8\] VGND VGND VPWR VPWR net1874 sky130_fd_sc_hd__dlygate4sd3_1
Xhold735 datamem.data_ram\[51\]\[5\] VGND VGND VPWR VPWR net1885 sky130_fd_sc_hd__dlygate4sd3_1
Xhold746 rvcpu.dp.rf.reg_file_arr\[11\]\[23\] VGND VGND VPWR VPWR net1896 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_57_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold757 rvcpu.dp.rf.reg_file_arr\[6\]\[26\] VGND VGND VPWR VPWR net1907 sky130_fd_sc_hd__dlygate4sd3_1
X_20161_ datamem.data_ram\[18\]\[27\] _06728_ _06768_ datamem.data_ram\[21\]\[27\]
+ VGND VGND VPWR VPWR _07454_ sky130_fd_sc_hd__o22a_1
Xhold768 rvcpu.dp.rf.reg_file_arr\[19\]\[1\] VGND VGND VPWR VPWR net1918 sky130_fd_sc_hd__dlygate4sd3_1
X_32147_ clknet_leaf_210_clk _03569_ VGND VGND VPWR VPWR datamem.data_ram\[38\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold779 rvcpu.dp.pcreg.q\[27\] VGND VGND VPWR VPWR net1929 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_123_Right_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2103 datamem.data_ram\[12\]\[17\] VGND VGND VPWR VPWR net3253 sky130_fd_sc_hd__dlygate4sd3_1
X_32078_ clknet_leaf_93_clk _03500_ VGND VGND VPWR VPWR datamem.data_ram\[33\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2114 rvcpu.dp.rf.reg_file_arr\[8\]\[5\] VGND VGND VPWR VPWR net3264 sky130_fd_sc_hd__dlygate4sd3_1
X_20092_ datamem.data_ram\[56\]\[10\] _06811_ _06685_ datamem.data_ram\[60\]\[10\]
+ _07385_ VGND VGND VPWR VPWR _07386_ sky130_fd_sc_hd__o221a_1
XFILLER_0_225_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2125 datamem.data_ram\[54\]\[11\] VGND VGND VPWR VPWR net3275 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2136 datamem.data_ram\[27\]\[19\] VGND VGND VPWR VPWR net3286 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_205_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_205_clk
+ sky130_fd_sc_hd__clkbuf_8
X_31029_ clknet_leaf_102_clk _02764_ VGND VGND VPWR VPWR datamem.data_ram\[12\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2147 datamem.data_ram\[51\]\[23\] VGND VGND VPWR VPWR net3297 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1402 rvcpu.dp.rf.reg_file_arr\[2\]\[2\] VGND VGND VPWR VPWR net2552 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2158 datamem.data_ram\[12\]\[13\] VGND VGND VPWR VPWR net3308 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1413 datamem.data_ram\[35\]\[14\] VGND VGND VPWR VPWR net2563 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1424 rvcpu.dp.rf.reg_file_arr\[26\]\[29\] VGND VGND VPWR VPWR net2574 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2169 rvcpu.dp.rf.reg_file_arr\[23\]\[5\] VGND VGND VPWR VPWR net3319 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1435 datamem.data_ram\[62\]\[9\] VGND VGND VPWR VPWR net2585 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1446 datamem.data_ram\[20\]\[29\] VGND VGND VPWR VPWR net2596 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1457 datamem.data_ram\[11\]\[8\] VGND VGND VPWR VPWR net2607 sky130_fd_sc_hd__dlygate4sd3_1
X_23851_ clknet_1_1__leaf__10203_ VGND VGND VPWR VPWR _10219_ sky130_fd_sc_hd__buf_1
Xhold1468 rvcpu.dp.rf.reg_file_arr\[12\]\[25\] VGND VGND VPWR VPWR net2618 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_224_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1479 datamem.data_ram\[6\]\[14\] VGND VGND VPWR VPWR net2629 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_212_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_200_5286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23111__789 clknet_1_0__leaf__10104_ VGND VGND VPWR VPWR net915 sky130_fd_sc_hd__inv_2
X_22802_ _09422_ _09941_ _09472_ VGND VGND VPWR VPWR _09942_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_200_5297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26570_ _11630_ VGND VGND VPWR VPWR _03229_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_196_5190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20994_ _06917_ _08277_ _08282_ _06675_ VGND VGND VPWR VPWR _08283_ sky130_fd_sc_hd__o211a_1
XFILLER_0_196_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25521_ _10418_ _11010_ VGND VGND VPWR VPWR _11017_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22733_ rvcpu.dp.rf.reg_file_arr\[8\]\[22\] rvcpu.dp.rf.reg_file_arr\[10\]\[22\]
+ rvcpu.dp.rf.reg_file_arr\[9\]\[22\] rvcpu.dp.rf.reg_file_arr\[11\]\[22\] _09418_
+ _09453_ VGND VGND VPWR VPWR _09877_ sky130_fd_sc_hd__mux4_1
XFILLER_0_211_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23758__347 clknet_1_0__leaf__10201_ VGND VGND VPWR VPWR net473 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_220_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_213_5603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_192_5098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28240_ _12589_ VGND VGND VPWR VPWR _03940_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_213_5614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25452_ _10064_ _10981_ _10982_ net1347 VGND VGND VPWR VPWR _02759_ sky130_fd_sc_hd__a22o_1
XFILLER_0_192_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22664_ _09481_ _09811_ VGND VGND VPWR VPWR _09812_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21615_ rvcpu.dp.rf.reg_file_arr\[16\]\[12\] rvcpu.dp.rf.reg_file_arr\[17\]\[12\]
+ rvcpu.dp.rf.reg_file_arr\[18\]\[12\] rvcpu.dp.rf.reg_file_arr\[19\]\[12\] _08516_
+ _08518_ VGND VGND VPWR VPWR _08865_ sky130_fd_sc_hd__mux4_1
XFILLER_0_34_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24403_ _09282_ net3981 _10376_ VGND VGND VPWR VPWR _10381_ sky130_fd_sc_hd__mux2_1
X_28171_ _12552_ VGND VGND VPWR VPWR _03908_ sky130_fd_sc_hd__clkbuf_1
X_25383_ _10938_ net1511 _10934_ _10943_ VGND VGND VPWR VPWR _02729_ sky130_fd_sc_hd__a31o_1
X_22595_ rvcpu.dp.rf.reg_file_arr\[24\]\[15\] rvcpu.dp.rf.reg_file_arr\[25\]\[15\]
+ rvcpu.dp.rf.reg_file_arr\[26\]\[15\] rvcpu.dp.rf.reg_file_arr\[27\]\[15\] _09393_
+ _09465_ VGND VGND VPWR VPWR _09746_ sky130_fd_sc_hd__mux4_1
XFILLER_0_180_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27122_ _11833_ _11953_ VGND VGND VPWR VPWR _11960_ sky130_fd_sc_hd__and2_1
XFILLER_0_180_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24334_ _10343_ VGND VGND VPWR VPWR _02280_ sky130_fd_sc_hd__clkbuf_1
X_21546_ rvcpu.dp.plfd.InstrD\[15\] VGND VGND VPWR VPWR _08799_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_106_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_209_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_181_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27053_ _11833_ _11911_ VGND VGND VPWR VPWR _11917_ sky130_fd_sc_hd__and2_1
X_24265_ _09326_ net2241 _10298_ VGND VGND VPWR VPWR _10305_ sky130_fd_sc_hd__mux2_1
X_21477_ _08542_ _08733_ VGND VGND VPWR VPWR _08734_ sky130_fd_sc_hd__or2_1
XFILLER_0_205_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26004_ _09476_ _11153_ VGND VGND VPWR VPWR _11327_ sky130_fd_sc_hd__nand2_1
X_20428_ datamem.data_ram\[13\]\[12\] _06663_ _06647_ datamem.data_ram\[8\]\[12\]
+ VGND VGND VPWR VPWR _07720_ sky130_fd_sc_hd__o22a_1
XFILLER_0_132_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_164_4422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20359_ datamem.data_ram\[13\]\[28\] _06724_ _06742_ _07650_ VGND VGND VPWR VPWR
+ _07651_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_164_4433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27955_ _09223_ VGND VGND VPWR VPWR _12430_ sky130_fd_sc_hd__clkbuf_2
X_23078_ _09291_ net3990 _10093_ VGND VGND VPWR VPWR _10101_ sky130_fd_sc_hd__mux2_1
XFILLER_0_179_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26906_ _11813_ net1391 _11821_ _11828_ VGND VGND VPWR VPWR _03367_ sky130_fd_sc_hd__a31o_1
X_14920_ rvcpu.dp.pcreg.q\[9\] _13368_ VGND VGND VPWR VPWR _13469_ sky130_fd_sc_hd__nand2_4
X_22029_ _09253_ VGND VGND VPWR VPWR _01065_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_175_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27886_ _12392_ VGND VGND VPWR VPWR _12393_ sky130_fd_sc_hd__buf_2
Xhold40 rvcpu.dp.plem.lAuiPCM\[26\] VGND VGND VPWR VPWR net1190 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold51 rvcpu.dp.plde.PCPlus4E\[22\] VGND VGND VPWR VPWR net1201 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_199_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold62 rvcpu.dp.plem.PCPlus4M\[31\] VGND VGND VPWR VPWR net1212 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2670 datamem.data_ram\[23\]\[28\] VGND VGND VPWR VPWR net3820 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_67_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29625_ net979 _01360_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[25\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_26837_ _09351_ _10921_ _10922_ VGND VGND VPWR VPWR _11786_ sky130_fd_sc_hd__and3_1
X_14851_ _13398_ _13357_ _13403_ rvcpu.dp.pcreg.q\[9\] VGND VGND VPWR VPWR _13404_
+ sky130_fd_sc_hd__o31a_1
Xhold73 rvcpu.dp.plem.PCPlus4M\[27\] VGND VGND VPWR VPWR net1223 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2681 datamem.data_ram\[3\]\[29\] VGND VGND VPWR VPWR net3831 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_67_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2692 datamem.data_ram\[56\]\[14\] VGND VGND VPWR VPWR net3842 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 rvcpu.dp.plem.PCPlus4M\[9\] VGND VGND VPWR VPWR net1234 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_123_3440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold95 rvcpu.dp.plem.PCPlus4M\[8\] VGND VGND VPWR VPWR net1245 sky130_fd_sc_hd__dlygate4sd3_1
X_24138__643 clknet_1_0__leaf__10261_ VGND VGND VPWR VPWR net769 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_123_3451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23544__169 clknet_1_1__leaf__10173_ VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__inv_2
Xhold1980 datamem.data_ram\[9\]\[15\] VGND VGND VPWR VPWR net3130 sky130_fd_sc_hd__dlygate4sd3_1
X_17570_ _05055_ VGND VGND VPWR VPWR _01251_ sky130_fd_sc_hd__clkbuf_1
X_29556_ net910 _01291_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[27\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_26768_ _11687_ _11738_ VGND VGND VPWR VPWR _11744_ sky130_fd_sc_hd__and2_1
X_14782_ _13334_ VGND VGND VPWR VPWR _13335_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_187_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1991 datamem.data_ram\[33\]\[28\] VGND VGND VPWR VPWR net3141 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_63_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16521_ _04498_ VGND VGND VPWR VPWR _01783_ sky130_fd_sc_hd__clkbuf_1
X_28507_ _12739_ net3897 net43 VGND VGND VPWR VPWR _12740_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_63_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23086__766 clknet_1_1__leaf__10102_ VGND VGND VPWR VPWR net892 sky130_fd_sc_hd__inv_2
X_25719_ _10113_ _11123_ _10998_ VGND VGND VPWR VPWR _11133_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_196_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29487_ net849 _01222_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[2\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_26699_ _10741_ _11123_ _10998_ VGND VGND VPWR VPWR _11704_ sky130_fd_sc_hd__a21oi_4
X_19240_ _06542_ _06544_ VGND VGND VPWR VPWR _06545_ sky130_fd_sc_hd__xnor2_1
X_23817__400 clknet_1_1__leaf__10207_ VGND VGND VPWR VPWR net526 sky130_fd_sc_hd__inv_2
X_28438_ _12699_ VGND VGND VPWR VPWR _04028_ sky130_fd_sc_hd__clkbuf_1
X_16452_ net2462 _14482_ _04451_ VGND VGND VPWR VPWR _04461_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__10199_ clknet_0__10199_ VGND VGND VPWR VPWR clknet_1_1__leaf__10199_
+ sky130_fd_sc_hd__clkbuf_16
X_15403_ _13483_ _13416_ _13741_ _13921_ _13934_ VGND VGND VPWR VPWR _13935_ sky130_fd_sc_hd__o311a_1
XFILLER_0_13_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19171_ _06484_ rvcpu.dp.plde.ImmExtE\[19\] _06419_ VGND VGND VPWR VPWR _06485_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28369_ _12355_ net2880 _12659_ VGND VGND VPWR VPWR _12660_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16383_ _14556_ VGND VGND VPWR VPWR _01847_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_225_Right_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18122_ rvcpu.dp.plem.ALUResultM\[18\] _05339_ _05340_ _13222_ VGND VGND VPWR VPWR
+ _05489_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_22_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30400_ net738 _02135_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[31\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_15334_ _13410_ _13416_ _13590_ _13863_ _13870_ VGND VGND VPWR VPWR _13871_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_22_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31380_ clknet_leaf_22_clk _03083_ VGND VGND VPWR VPWR rvcpu.dp.plde.ImmExtE\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_206_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18053_ _13253_ rvcpu.dp.plde.RD2E\[8\] _05195_ VGND VGND VPWR VPWR _05422_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_117_3299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30331_ net677 _02066_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[4\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_15265_ _13784_ _13790_ _13804_ VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_10_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_4 _02993_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17004_ _04754_ VGND VGND VPWR VPWR _01540_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_227_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30262_ net616 _01997_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[6\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_15196_ _13301_ _13488_ _13550_ _13646_ VGND VGND VPWR VPWR _13738_ sky130_fd_sc_hd__o31a_1
Xclkbuf_1_0__f__10090_ clknet_0__10090_ VGND VGND VPWR VPWR clknet_1_0__leaf__10090_
+ sky130_fd_sc_hd__clkbuf_16
X_32001_ clknet_leaf_133_clk _03423_ VGND VGND VPWR VPWR datamem.data_ram\[52\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_675 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30193_ net547 _01928_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[8\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18955_ _05547_ _06291_ _05543_ VGND VGND VPWR VPWR _06292_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_52_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_52_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17906_ _05278_ VGND VGND VPWR VPWR _05279_ sky130_fd_sc_hd__clkbuf_4
X_18886_ _05624_ _06212_ _05467_ VGND VGND VPWR VPWR _06228_ sky130_fd_sc_hd__a21o_1
XFILLER_0_158_1337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17837_ _13219_ rvcpu.dp.plde.RD2E\[19\] _05195_ VGND VGND VPWR VPWR _05219_ sky130_fd_sc_hd__mux2_1
X_32903_ clknet_leaf_208_clk _04325_ VGND VGND VPWR VPWR datamem.data_ram\[0\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_179_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23030__732 clknet_1_1__leaf__10088_ VGND VGND VPWR VPWR net858 sky130_fd_sc_hd__inv_2
X_32834_ clknet_leaf_285_clk _04256_ VGND VGND VPWR VPWR datamem.data_ram\[12\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_222_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17768_ rvcpu.dp.plem.RdM\[2\] rvcpu.dp.plde.Rs2E\[2\] VGND VGND VPWR VPWR _05166_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_178_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_530 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16719_ _14183_ net2600 _04598_ VGND VGND VPWR VPWR _04604_ sky130_fd_sc_hd__mux2_1
X_19507_ _06802_ VGND VGND VPWR VPWR _06803_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_187_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32765_ clknet_leaf_286_clk _04187_ VGND VGND VPWR VPWR datamem.data_ram\[15\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17699_ _13198_ net2634 _05118_ VGND VGND VPWR VPWR _05124_ sky130_fd_sc_hd__mux2_1
XFILLER_0_190_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19438_ datamem.data_ram\[34\]\[16\] _06728_ _06731_ datamem.data_ram\[35\]\[16\]
+ _06733_ VGND VGND VPWR VPWR _06734_ sky130_fd_sc_hd__o221a_1
XFILLER_0_14_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31716_ net165 _03174_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[9\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32696_ clknet_leaf_283_clk _04118_ VGND VGND VPWR VPWR datamem.data_ram\[18\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31647_ clknet_leaf_25_clk net1216 VGND VGND VPWR VPWR rvcpu.dp.plmw.lAuiPCW\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_19369_ _06664_ VGND VGND VPWR VPWR _06665_ sky130_fd_sc_hd__buf_4
XFILLER_0_18_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21400_ _08515_ _08659_ _08513_ VGND VGND VPWR VPWR _08660_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_210_1280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22380_ _09451_ _09541_ _09404_ VGND VGND VPWR VPWR _09542_ sky130_fd_sc_hd__o21a_1
X_31578_ clknet_leaf_75_clk datamem.rd_data_mem\[28\] VGND VGND VPWR VPWR rvcpu.dp.plmw.ReadDataW\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_21331_ _08592_ rvcpu.dp.plde.RdE\[0\] VGND VGND VPWR VPWR _08593_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_30529_ clknet_leaf_268_clk _02264_ VGND VGND VPWR VPWR datamem.data_ram\[56\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold510 rvcpu.dp.plfd.PCPlus4D\[3\] VGND VGND VPWR VPWR net1660 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21262_ rvcpu.dp.plfd.InstrD\[15\] VGND VGND VPWR VPWR _08524_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_13_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold521 rvcpu.dp.plfd.PCPlus4D\[16\] VGND VGND VPWR VPWR net1671 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_229_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold532 datamem.data_ram\[10\]\[2\] VGND VGND VPWR VPWR net1682 sky130_fd_sc_hd__dlygate4sd3_1
Xhold543 datamem.data_ram\[51\]\[4\] VGND VGND VPWR VPWR net1693 sky130_fd_sc_hd__dlygate4sd3_1
X_20213_ _05391_ _06586_ _07461_ net37 _07120_ VGND VGND VPWR VPWR _07506_ sky130_fd_sc_hd__o32a_1
XFILLER_0_130_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold554 datamem.data_ram\[26\]\[2\] VGND VGND VPWR VPWR net1704 sky130_fd_sc_hd__dlygate4sd3_1
Xhold565 datamem.data_ram\[11\]\[5\] VGND VGND VPWR VPWR net1715 sky130_fd_sc_hd__dlygate4sd3_1
X_21193_ _08477_ VGND VGND VPWR VPWR _04416_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_229_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold576 datamem.data_ram\[31\]\[7\] VGND VGND VPWR VPWR net1726 sky130_fd_sc_hd__dlygate4sd3_1
Xhold587 datamem.data_ram\[23\]\[3\] VGND VGND VPWR VPWR net1737 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_206_5440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold598 datamem.data_ram\[61\]\[0\] VGND VGND VPWR VPWR net1748 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_206_5451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20144_ _06714_ _07431_ _07436_ VGND VGND VPWR VPWR _07437_ sky130_fd_sc_hd__or3_2
XFILLER_0_229_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_218_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27740_ _12309_ VGND VGND VPWR VPWR _03720_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_202_5337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24952_ _10454_ net2292 _10687_ VGND VGND VPWR VPWR _10695_ sky130_fd_sc_hd__mux2_1
X_20075_ datamem.data_ram\[46\]\[10\] _06718_ _06656_ datamem.data_ram\[41\]\[10\]
+ VGND VGND VPWR VPWR _07369_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_202_5348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_198_5241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1210 datamem.data_ram\[16\]\[16\] VGND VGND VPWR VPWR net2360 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_198_5252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1221 rvcpu.dp.rf.reg_file_arr\[11\]\[7\] VGND VGND VPWR VPWR net2371 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1232 datamem.data_ram\[43\]\[27\] VGND VGND VPWR VPWR net2382 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1243 datamem.data_ram\[41\]\[23\] VGND VGND VPWR VPWR net2393 sky130_fd_sc_hd__dlygate4sd3_1
X_27671_ _12272_ VGND VGND VPWR VPWR _03688_ sky130_fd_sc_hd__clkbuf_1
X_23463__112 clknet_1_1__leaf__10157_ VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__inv_2
X_24883_ _10480_ net1951 net92 VGND VGND VPWR VPWR _10658_ sky130_fd_sc_hd__mux2_1
Xhold1254 rvcpu.dp.rf.reg_file_arr\[18\]\[0\] VGND VGND VPWR VPWR net2404 sky130_fd_sc_hd__dlygate4sd3_1
X_29410_ clknet_leaf_290_clk _01145_ VGND VGND VPWR VPWR rvcpu.dp.plde.RD2E\[21\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1265 rvcpu.dp.rf.reg_file_arr\[19\]\[12\] VGND VGND VPWR VPWR net2415 sky130_fd_sc_hd__dlygate4sd3_1
X_26622_ _10600_ _10947_ VGND VGND VPWR VPWR _11659_ sky130_fd_sc_hd__nor2_4
Xhold1276 datamem.data_ram\[39\]\[11\] VGND VGND VPWR VPWR net2426 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_194_5149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23834_ _10213_ VGND VGND VPWR VPWR _01910_ sky130_fd_sc_hd__clkbuf_1
Xhold1287 datamem.data_ram\[63\]\[24\] VGND VGND VPWR VPWR net2437 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1298 datamem.data_ram\[7\]\[15\] VGND VGND VPWR VPWR net2448 sky130_fd_sc_hd__dlygate4sd3_1
X_23992__526 clknet_1_1__leaf__10240_ VGND VGND VPWR VPWR net652 sky130_fd_sc_hd__inv_2
XANTENNA_405 _06643_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0__10222_ _10222_ VGND VGND VPWR VPWR clknet_0__10222_ sky130_fd_sc_hd__clkbuf_16
XANTENNA_416 _06732_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_427 _06790_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29341_ clknet_leaf_205_clk _01076_ VGND VGND VPWR VPWR datamem.data_ram\[61\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_438 _06934_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26553_ _11621_ VGND VGND VPWR VPWR _03221_ sky130_fd_sc_hd__clkbuf_1
X_20977_ net122 datamem.data_ram\[47\]\[15\] _06639_ datamem.data_ram\[46\]\[15\]
+ _07838_ VGND VGND VPWR VPWR _08266_ sky130_fd_sc_hd__a221o_1
XANTENNA_449 _07860_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_0__10153_ _10153_ VGND VGND VPWR VPWR clknet_0__10153_ sky130_fd_sc_hd__clkbuf_16
X_25504_ _10826_ net2907 _10999_ VGND VGND VPWR VPWR _11007_ sky130_fd_sc_hd__mux2_1
X_22716_ _09636_ _09860_ VGND VGND VPWR VPWR _09861_ sky130_fd_sc_hd__or2_1
X_29272_ _09287_ net4014 _13150_ VGND VGND VPWR VPWR _13157_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_157_4270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28223_ _12580_ VGND VGND VPWR VPWR _03932_ sky130_fd_sc_hd__clkbuf_1
X_23007__712 clknet_1_0__leaf__10085_ VGND VGND VPWR VPWR net838 sky130_fd_sc_hd__inv_2
X_25435_ _10758_ net4004 _10970_ VGND VGND VPWR VPWR _10974_ sky130_fd_sc_hd__mux2_1
Xclkbuf_0__10084_ _10084_ VGND VGND VPWR VPWR clknet_0__10084_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_211_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_153_4156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22647_ _09627_ _09792_ _09794_ _09795_ VGND VGND VPWR VPWR _09796_ sky130_fd_sc_hd__a211o_1
XFILLER_0_153_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_153_4167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_4178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28154_ _12543_ VGND VGND VPWR VPWR _03900_ sky130_fd_sc_hd__clkbuf_1
X_25366_ _08151_ VGND VGND VPWR VPWR _10932_ sky130_fd_sc_hd__clkbuf_8
X_22578_ _09495_ _09729_ VGND VGND VPWR VPWR _09730_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27105_ _11938_ net1772 _11940_ _11949_ VGND VGND VPWR VPWR _03445_ sky130_fd_sc_hd__a31o_1
XFILLER_0_35_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24317_ _09322_ net3092 _10328_ VGND VGND VPWR VPWR _10334_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28085_ _12441_ net3798 _12501_ VGND VGND VPWR VPWR _12507_ sky130_fd_sc_hd__mux2_1
X_21529_ rvcpu.dp.rf.reg_file_arr\[24\]\[8\] rvcpu.dp.rf.reg_file_arr\[25\]\[8\] rvcpu.dp.rf.reg_file_arr\[26\]\[8\]
+ rvcpu.dp.rf.reg_file_arr\[27\]\[8\] _08517_ _08519_ VGND VGND VPWR VPWR _08783_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_90_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25297_ _10891_ VGND VGND VPWR VPWR _02695_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27036_ _11835_ _11899_ VGND VGND VPWR VPWR _11907_ sky130_fd_sc_hd__and2_1
X_15050_ _13333_ _13370_ VGND VGND VPWR VPWR _13597_ sky130_fd_sc_hd__nand2_1
X_24248_ _10295_ VGND VGND VPWR VPWR _02242_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_112_3174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput6 net6 VGND VGND VPWR VPWR Instr[13] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_112_3185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput30 net30 VGND VGND VPWR VPWR Instr[6] sky130_fd_sc_hd__buf_2
XFILLER_0_102_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23315__955 clknet_1_1__leaf__10134_ VGND VGND VPWR VPWR net1081 sky130_fd_sc_hd__inv_2
XFILLER_0_82_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_183_4886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28987_ _12694_ net2975 _12999_ VGND VGND VPWR VPWR _13003_ sky130_fd_sc_hd__mux2_1
X_23927__483 clknet_1_0__leaf__10226_ VGND VGND VPWR VPWR net609 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_183_4897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18740_ _05436_ _05438_ _06069_ VGND VGND VPWR VPWR _06091_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_125_3502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27938_ _12178_ _12325_ _12356_ VGND VGND VPWR VPWR _12421_ sky130_fd_sc_hd__a21oi_4
X_15952_ net4145 _13184_ _14311_ VGND VGND VPWR VPWR _14313_ sky130_fd_sc_hd__mux2_1
XFILLER_0_207_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold3190 rvcpu.dp.rf.reg_file_arr\[29\]\[31\] VGND VGND VPWR VPWR net4340 sky130_fd_sc_hd__dlygate4sd3_1
X_14903_ _13287_ _13390_ VGND VGND VPWR VPWR _13454_ sky130_fd_sc_hd__nor2_1
X_23626__244 clknet_1_1__leaf__10180_ VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__inv_2
X_18671_ _05939_ _06025_ _05705_ VGND VGND VPWR VPWR _06026_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27869_ _12383_ VGND VGND VPWR VPWR _03775_ sky130_fd_sc_hd__clkbuf_1
X_15883_ _14276_ VGND VGND VPWR VPWR _02083_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_216_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17622_ _05083_ VGND VGND VPWR VPWR _01227_ sky130_fd_sc_hd__clkbuf_1
X_14834_ _13287_ VGND VGND VPWR VPWR _13387_ sky130_fd_sc_hd__clkbuf_4
X_29608_ net962 _01343_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[25\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_4_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30880_ clknet_leaf_262_clk _02615_ VGND VGND VPWR VPWR datamem.data_ram\[42\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_86_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_142_3893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29539_ net893 _01274_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[27\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_17553_ _13173_ net4125 _05046_ VGND VGND VPWR VPWR _05047_ sky130_fd_sc_hd__mux2_1
X_14765_ rvcpu.dp.pcreg.q\[8\] _13313_ VGND VGND VPWR VPWR _13318_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23209__860 clknet_1_1__leaf__10112_ VGND VGND VPWR VPWR net986 sky130_fd_sc_hd__inv_2
X_16504_ net2685 _14463_ _04489_ VGND VGND VPWR VPWR _04490_ sky130_fd_sc_hd__mux2_1
X_32550_ clknet_leaf_271_clk _03972_ VGND VGND VPWR VPWR datamem.data_ram\[23\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17484_ _05009_ VGND VGND VPWR VPWR _05010_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_224_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14696_ _13256_ VGND VGND VPWR VPWR _13257_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_168_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23361__997 clknet_1_1__leaf__10138_ VGND VGND VPWR VPWR net1123 sky130_fd_sc_hd__inv_2
XFILLER_0_86_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19223_ _06521_ _06522_ _06523_ VGND VGND VPWR VPWR _06530_ sky130_fd_sc_hd__a21boi_2
X_31501_ clknet_leaf_25_clk rvcpu.dp.lAuiPCE\[27\] VGND VGND VPWR VPWR rvcpu.dp.plem.lAuiPCM\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16435_ _04452_ VGND VGND VPWR VPWR _01823_ sky130_fd_sc_hd__clkbuf_1
X_32481_ clknet_leaf_231_clk _03903_ VGND VGND VPWR VPWR datamem.data_ram\[25\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_15_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31432_ clknet_leaf_103_clk _03135_ VGND VGND VPWR VPWR datamem.data_ram\[14\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_19154_ _06469_ VGND VGND VPWR VPWR rvcpu.dp.lAuiPCE\[17\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16366_ net3747 _14463_ _14547_ VGND VGND VPWR VPWR _14548_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18105_ _05471_ _05472_ VGND VGND VPWR VPWR _05473_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_41_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15317_ _13398_ _13672_ _13853_ VGND VGND VPWR VPWR _13854_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_124_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19085_ rvcpu.dp.plde.ImmExtE\[8\] rvcpu.dp.plde.PCE\[8\] VGND VGND VPWR VPWR _06409_
+ sky130_fd_sc_hd__and2_1
X_31363_ clknet_leaf_24_clk _03066_ VGND VGND VPWR VPWR rvcpu.dp.plde.ImmExtE\[12\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_41_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16297_ _14488_ VGND VGND VPWR VPWR _14511_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18036_ _05346_ _05405_ _05344_ VGND VGND VPWR VPWR _05406_ sky130_fd_sc_hd__a21o_1
X_30314_ net660 _02049_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[5\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_15248_ _13343_ _13321_ _13401_ _13354_ VGND VGND VPWR VPWR _13788_ sky130_fd_sc_hd__or4_1
XFILLER_0_160_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31294_ clknet_leaf_18_clk _02997_ VGND VGND VPWR VPWR rvcpu.dp.plde.BranchE sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30245_ net599 _01980_ VGND VGND VPWR VPWR rvcpu.dp.rf.reg_file_arr\[6\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_15179_ _13401_ _13323_ _13721_ _13492_ _13321_ VGND VGND VPWR VPWR _13722_ sky130_fd_sc_hd__o32a_1
X_23787__373 clknet_1_1__leaf__10204_ VGND VGND VPWR VPWR net499 sky130_fd_sc_hd__inv_2
XFILLER_0_10_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30176_ clknet_leaf_204_clk _01911_ VGND VGND VPWR VPWR datamem.data_ram\[58\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_19987_ datamem.data_ram\[12\]\[2\] _06954_ _07280_ _06679_ VGND VGND VPWR VPWR _07281_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_201_1268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18938_ _05634_ _06055_ _06267_ _06268_ _06276_ VGND VGND VPWR VPWR _06277_ sky130_fd_sc_hd__a41o_1
.ends

