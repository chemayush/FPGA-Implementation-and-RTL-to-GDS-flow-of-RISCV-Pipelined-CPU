VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO pl_riscv_cpu
  CLASS BLOCK ;
  FOREIGN pl_riscv_cpu ;
  ORIGIN 0.000 0.000 ;
  SIZE 638.325 BY 649.045 ;
  PIN Instr[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 4.000 469.840 ;
    END
  END Instr[0]
  PIN Instr[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.040 4.000 561.640 ;
    END
  END Instr[10]
  PIN Instr[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END Instr[11]
  PIN Instr[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 489.640 4.000 490.240 ;
    END
  END Instr[12]
  PIN Instr[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.840 4.000 500.440 ;
    END
  END Instr[13]
  PIN Instr[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.840 4.000 534.440 ;
    END
  END Instr[14]
  PIN Instr[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.040 4.000 527.640 ;
    END
  END Instr[15]
  PIN Instr[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 574.640 4.000 575.240 ;
    END
  END Instr[16]
  PIN Instr[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 4.000 493.640 ;
    END
  END Instr[17]
  PIN Instr[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 564.440 4.000 565.040 ;
    END
  END Instr[18]
  PIN Instr[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 479.440 4.000 480.040 ;
    END
  END Instr[19]
  PIN Instr[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END Instr[1]
  PIN Instr[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.240 4.000 571.840 ;
    END
  END Instr[20]
  PIN Instr[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 591.640 4.000 592.240 ;
    END
  END Instr[21]
  PIN Instr[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 557.640 4.000 558.240 ;
    END
  END Instr[22]
  PIN Instr[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 4.000 599.040 ;
    END
  END Instr[23]
  PIN Instr[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.840 4.000 517.440 ;
    END
  END Instr[24]
  PIN Instr[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 4.000 551.440 ;
    END
  END Instr[25]
  PIN Instr[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 540.640 4.000 541.240 ;
    END
  END Instr[26]
  PIN Instr[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.240 4.000 520.840 ;
    END
  END Instr[27]
  PIN Instr[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.040 4.000 476.640 ;
    END
  END Instr[28]
  PIN Instr[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 506.640 4.000 507.240 ;
    END
  END Instr[29]
  PIN Instr[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 472.640 4.000 473.240 ;
    END
  END Instr[2]
  PIN Instr[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.040 4.000 510.640 ;
    END
  END Instr[30]
  PIN Instr[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 513.440 4.000 514.040 ;
    END
  END Instr[31]
  PIN Instr[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.240 4.000 486.840 ;
    END
  END Instr[3]
  PIN Instr[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 547.440 4.000 548.040 ;
    END
  END Instr[4]
  PIN Instr[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END Instr[5]
  PIN Instr[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 530.440 4.000 531.040 ;
    END
  END Instr[6]
  PIN Instr[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.040 4.000 544.640 ;
    END
  END Instr[7]
  PIN Instr[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END Instr[8]
  PIN Instr[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END Instr[9]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 10.640 333.140 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 10.640 486.740 636.720 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 632.740 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 632.740 184.810 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 336.390 632.740 337.990 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 489.570 632.740 491.170 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 636.720 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 632.740 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 632.740 181.510 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 333.090 632.740 334.690 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 486.270 632.740 487.870 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 634.325 71.440 638.325 72.040 ;
    END
  END clk
  PIN correct
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 634.325 340.040 638.325 340.640 ;
    END
  END correct
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 328.530 645.045 328.810 649.045 ;
    END
  END reset
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 632.690 636.565 ;
      LAYER li1 ;
        RECT 5.520 10.795 632.500 636.565 ;
      LAYER met1 ;
        RECT 2.370 10.640 634.270 637.120 ;
      LAYER met2 ;
        RECT 2.390 644.765 328.250 645.730 ;
        RECT 329.090 644.765 634.250 645.730 ;
        RECT 2.390 10.695 634.250 644.765 ;
      LAYER met3 ;
        RECT 2.110 599.440 634.325 636.645 ;
        RECT 4.400 598.040 634.325 599.440 ;
        RECT 2.110 592.640 634.325 598.040 ;
        RECT 4.400 591.240 634.325 592.640 ;
        RECT 2.110 575.640 634.325 591.240 ;
        RECT 4.400 574.240 634.325 575.640 ;
        RECT 2.110 572.240 634.325 574.240 ;
        RECT 4.400 570.840 634.325 572.240 ;
        RECT 2.110 565.440 634.325 570.840 ;
        RECT 4.400 564.040 634.325 565.440 ;
        RECT 2.110 562.040 634.325 564.040 ;
        RECT 4.400 560.640 634.325 562.040 ;
        RECT 2.110 558.640 634.325 560.640 ;
        RECT 4.400 557.240 634.325 558.640 ;
        RECT 2.110 551.840 634.325 557.240 ;
        RECT 4.400 550.440 634.325 551.840 ;
        RECT 2.110 548.440 634.325 550.440 ;
        RECT 4.400 547.040 634.325 548.440 ;
        RECT 2.110 545.040 634.325 547.040 ;
        RECT 4.400 543.640 634.325 545.040 ;
        RECT 2.110 541.640 634.325 543.640 ;
        RECT 4.400 540.240 634.325 541.640 ;
        RECT 2.110 538.240 634.325 540.240 ;
        RECT 4.400 536.840 634.325 538.240 ;
        RECT 2.110 534.840 634.325 536.840 ;
        RECT 4.400 533.440 634.325 534.840 ;
        RECT 2.110 531.440 634.325 533.440 ;
        RECT 4.400 530.040 634.325 531.440 ;
        RECT 2.110 528.040 634.325 530.040 ;
        RECT 4.400 526.640 634.325 528.040 ;
        RECT 2.110 524.640 634.325 526.640 ;
        RECT 4.400 523.240 634.325 524.640 ;
        RECT 2.110 521.240 634.325 523.240 ;
        RECT 4.400 519.840 634.325 521.240 ;
        RECT 2.110 517.840 634.325 519.840 ;
        RECT 4.400 516.440 634.325 517.840 ;
        RECT 2.110 514.440 634.325 516.440 ;
        RECT 4.400 513.040 634.325 514.440 ;
        RECT 2.110 511.040 634.325 513.040 ;
        RECT 4.400 509.640 634.325 511.040 ;
        RECT 2.110 507.640 634.325 509.640 ;
        RECT 4.400 506.240 634.325 507.640 ;
        RECT 2.110 504.240 634.325 506.240 ;
        RECT 4.400 502.840 634.325 504.240 ;
        RECT 2.110 500.840 634.325 502.840 ;
        RECT 4.400 499.440 634.325 500.840 ;
        RECT 2.110 497.440 634.325 499.440 ;
        RECT 4.400 496.040 634.325 497.440 ;
        RECT 2.110 494.040 634.325 496.040 ;
        RECT 4.400 492.640 634.325 494.040 ;
        RECT 2.110 490.640 634.325 492.640 ;
        RECT 4.400 489.240 634.325 490.640 ;
        RECT 2.110 487.240 634.325 489.240 ;
        RECT 4.400 485.840 634.325 487.240 ;
        RECT 2.110 483.840 634.325 485.840 ;
        RECT 4.400 482.440 634.325 483.840 ;
        RECT 2.110 480.440 634.325 482.440 ;
        RECT 4.400 479.040 634.325 480.440 ;
        RECT 2.110 477.040 634.325 479.040 ;
        RECT 4.400 475.640 634.325 477.040 ;
        RECT 2.110 473.640 634.325 475.640 ;
        RECT 4.400 472.240 634.325 473.640 ;
        RECT 2.110 470.240 634.325 472.240 ;
        RECT 4.400 468.840 634.325 470.240 ;
        RECT 2.110 341.040 634.325 468.840 ;
        RECT 2.110 339.640 633.925 341.040 ;
        RECT 2.110 72.440 634.325 339.640 ;
        RECT 2.110 71.040 633.925 72.440 ;
        RECT 2.110 10.715 634.325 71.040 ;
      LAYER met4 ;
        RECT 1.710 19.895 20.640 635.625 ;
        RECT 23.040 19.895 23.940 635.625 ;
        RECT 26.340 19.895 174.240 635.625 ;
        RECT 176.640 19.895 177.540 635.625 ;
        RECT 179.940 19.895 327.840 635.625 ;
        RECT 330.240 19.895 331.140 635.625 ;
        RECT 333.540 19.895 481.440 635.625 ;
        RECT 483.840 19.895 484.740 635.625 ;
        RECT 487.140 19.895 626.225 635.625 ;
      LAYER met5 ;
        RECT 1.500 492.770 613.060 624.700 ;
        RECT 1.500 484.670 3.680 492.770 ;
        RECT 1.500 339.590 613.060 484.670 ;
        RECT 1.500 331.490 3.680 339.590 ;
        RECT 1.500 186.410 613.060 331.490 ;
        RECT 1.500 178.310 3.680 186.410 ;
        RECT 1.500 99.500 613.060 178.310 ;
  END
END pl_riscv_cpu
END LIBRARY

