module pl_riscv_cpu (clk,
    correct,
    reset,
    Instr);
 input clk;
 output correct;
 input reset;
 output [31:0] Instr;

 wire _00000_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire _14291_;
 wire _14292_;
 wire _14293_;
 wire _14294_;
 wire _14295_;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14300_;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire _14308_;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire _14321_;
 wire _14322_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14333_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14340_;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14355_;
 wire _14356_;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire _14365_;
 wire _14366_;
 wire _14367_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire _14374_;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire _14378_;
 wire _14379_;
 wire _14380_;
 wire _14381_;
 wire _14382_;
 wire _14383_;
 wire _14384_;
 wire _14385_;
 wire _14386_;
 wire _14387_;
 wire _14388_;
 wire _14389_;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire _14393_;
 wire _14394_;
 wire _14395_;
 wire _14396_;
 wire _14397_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14402_;
 wire _14403_;
 wire _14404_;
 wire _14405_;
 wire _14406_;
 wire _14407_;
 wire _14408_;
 wire _14409_;
 wire _14410_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire _14415_;
 wire _14416_;
 wire _14417_;
 wire _14418_;
 wire _14419_;
 wire _14420_;
 wire _14421_;
 wire _14422_;
 wire _14423_;
 wire _14424_;
 wire _14425_;
 wire _14426_;
 wire _14427_;
 wire _14428_;
 wire _14429_;
 wire _14430_;
 wire _14431_;
 wire _14432_;
 wire _14433_;
 wire _14434_;
 wire _14435_;
 wire _14436_;
 wire _14437_;
 wire _14438_;
 wire _14439_;
 wire _14440_;
 wire _14441_;
 wire _14442_;
 wire _14443_;
 wire _14444_;
 wire _14445_;
 wire _14446_;
 wire _14447_;
 wire _14448_;
 wire _14449_;
 wire _14450_;
 wire _14451_;
 wire _14452_;
 wire _14453_;
 wire _14454_;
 wire _14455_;
 wire _14456_;
 wire _14457_;
 wire _14458_;
 wire _14459_;
 wire _14460_;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire _14464_;
 wire _14465_;
 wire _14466_;
 wire _14467_;
 wire _14468_;
 wire _14469_;
 wire _14470_;
 wire _14471_;
 wire _14472_;
 wire _14473_;
 wire _14474_;
 wire _14475_;
 wire _14476_;
 wire _14477_;
 wire _14478_;
 wire _14479_;
 wire _14480_;
 wire _14481_;
 wire _14482_;
 wire _14483_;
 wire _14484_;
 wire _14485_;
 wire _14486_;
 wire _14487_;
 wire _14488_;
 wire _14489_;
 wire _14490_;
 wire _14491_;
 wire _14492_;
 wire _14493_;
 wire _14494_;
 wire _14495_;
 wire _14496_;
 wire _14497_;
 wire _14498_;
 wire _14499_;
 wire _14500_;
 wire _14501_;
 wire _14502_;
 wire _14503_;
 wire _14504_;
 wire _14505_;
 wire _14506_;
 wire _14507_;
 wire _14508_;
 wire _14509_;
 wire _14510_;
 wire _14511_;
 wire _14512_;
 wire _14513_;
 wire _14514_;
 wire _14515_;
 wire _14516_;
 wire _14517_;
 wire _14518_;
 wire _14519_;
 wire _14520_;
 wire _14521_;
 wire _14522_;
 wire _14523_;
 wire _14524_;
 wire _14525_;
 wire _14526_;
 wire _14527_;
 wire _14528_;
 wire _14529_;
 wire _14530_;
 wire _14531_;
 wire _14532_;
 wire _14533_;
 wire _14534_;
 wire _14535_;
 wire _14536_;
 wire _14537_;
 wire _14538_;
 wire _14539_;
 wire _14540_;
 wire _14541_;
 wire _14542_;
 wire _14543_;
 wire _14544_;
 wire _14545_;
 wire _14546_;
 wire _14547_;
 wire _14548_;
 wire _14549_;
 wire _14550_;
 wire _14551_;
 wire _14552_;
 wire _14553_;
 wire _14554_;
 wire _14555_;
 wire _14556_;
 wire _14557_;
 wire _14558_;
 wire _14559_;
 wire _14560_;
 wire _14561_;
 wire _14562_;
 wire _14563_;
 wire _14564_;
 wire _14565_;
 wire _14566_;
 wire _14567_;
 wire _14568_;
 wire _14569_;
 wire _14570_;
 wire _14571_;
 wire _14572_;
 wire _14573_;
 wire _14574_;
 wire _14575_;
 wire _14576_;
 wire _14577_;
 wire _14578_;
 wire _14579_;
 wire _14580_;
 wire _14581_;
 wire _14582_;
 wire \datamem.data_ram[0][0] ;
 wire \datamem.data_ram[0][10] ;
 wire \datamem.data_ram[0][11] ;
 wire \datamem.data_ram[0][12] ;
 wire \datamem.data_ram[0][13] ;
 wire \datamem.data_ram[0][14] ;
 wire \datamem.data_ram[0][15] ;
 wire \datamem.data_ram[0][16] ;
 wire \datamem.data_ram[0][17] ;
 wire \datamem.data_ram[0][18] ;
 wire \datamem.data_ram[0][19] ;
 wire \datamem.data_ram[0][1] ;
 wire \datamem.data_ram[0][20] ;
 wire \datamem.data_ram[0][21] ;
 wire \datamem.data_ram[0][22] ;
 wire \datamem.data_ram[0][23] ;
 wire \datamem.data_ram[0][24] ;
 wire \datamem.data_ram[0][25] ;
 wire \datamem.data_ram[0][26] ;
 wire \datamem.data_ram[0][27] ;
 wire \datamem.data_ram[0][28] ;
 wire \datamem.data_ram[0][29] ;
 wire \datamem.data_ram[0][2] ;
 wire \datamem.data_ram[0][30] ;
 wire \datamem.data_ram[0][31] ;
 wire \datamem.data_ram[0][3] ;
 wire \datamem.data_ram[0][4] ;
 wire \datamem.data_ram[0][5] ;
 wire \datamem.data_ram[0][6] ;
 wire \datamem.data_ram[0][7] ;
 wire \datamem.data_ram[0][8] ;
 wire \datamem.data_ram[0][9] ;
 wire \datamem.data_ram[10][0] ;
 wire \datamem.data_ram[10][10] ;
 wire \datamem.data_ram[10][11] ;
 wire \datamem.data_ram[10][12] ;
 wire \datamem.data_ram[10][13] ;
 wire \datamem.data_ram[10][14] ;
 wire \datamem.data_ram[10][15] ;
 wire \datamem.data_ram[10][16] ;
 wire \datamem.data_ram[10][17] ;
 wire \datamem.data_ram[10][18] ;
 wire \datamem.data_ram[10][19] ;
 wire \datamem.data_ram[10][1] ;
 wire \datamem.data_ram[10][20] ;
 wire \datamem.data_ram[10][21] ;
 wire \datamem.data_ram[10][22] ;
 wire \datamem.data_ram[10][23] ;
 wire \datamem.data_ram[10][24] ;
 wire \datamem.data_ram[10][25] ;
 wire \datamem.data_ram[10][26] ;
 wire \datamem.data_ram[10][27] ;
 wire \datamem.data_ram[10][28] ;
 wire \datamem.data_ram[10][29] ;
 wire \datamem.data_ram[10][2] ;
 wire \datamem.data_ram[10][30] ;
 wire \datamem.data_ram[10][31] ;
 wire \datamem.data_ram[10][3] ;
 wire \datamem.data_ram[10][4] ;
 wire \datamem.data_ram[10][5] ;
 wire \datamem.data_ram[10][6] ;
 wire \datamem.data_ram[10][7] ;
 wire \datamem.data_ram[10][8] ;
 wire \datamem.data_ram[10][9] ;
 wire \datamem.data_ram[11][0] ;
 wire \datamem.data_ram[11][10] ;
 wire \datamem.data_ram[11][11] ;
 wire \datamem.data_ram[11][12] ;
 wire \datamem.data_ram[11][13] ;
 wire \datamem.data_ram[11][14] ;
 wire \datamem.data_ram[11][15] ;
 wire \datamem.data_ram[11][16] ;
 wire \datamem.data_ram[11][17] ;
 wire \datamem.data_ram[11][18] ;
 wire \datamem.data_ram[11][19] ;
 wire \datamem.data_ram[11][1] ;
 wire \datamem.data_ram[11][20] ;
 wire \datamem.data_ram[11][21] ;
 wire \datamem.data_ram[11][22] ;
 wire \datamem.data_ram[11][23] ;
 wire \datamem.data_ram[11][24] ;
 wire \datamem.data_ram[11][25] ;
 wire \datamem.data_ram[11][26] ;
 wire \datamem.data_ram[11][27] ;
 wire \datamem.data_ram[11][28] ;
 wire \datamem.data_ram[11][29] ;
 wire \datamem.data_ram[11][2] ;
 wire \datamem.data_ram[11][30] ;
 wire \datamem.data_ram[11][31] ;
 wire \datamem.data_ram[11][3] ;
 wire \datamem.data_ram[11][4] ;
 wire \datamem.data_ram[11][5] ;
 wire \datamem.data_ram[11][6] ;
 wire \datamem.data_ram[11][7] ;
 wire \datamem.data_ram[11][8] ;
 wire \datamem.data_ram[11][9] ;
 wire \datamem.data_ram[12][0] ;
 wire \datamem.data_ram[12][10] ;
 wire \datamem.data_ram[12][11] ;
 wire \datamem.data_ram[12][12] ;
 wire \datamem.data_ram[12][13] ;
 wire \datamem.data_ram[12][14] ;
 wire \datamem.data_ram[12][15] ;
 wire \datamem.data_ram[12][16] ;
 wire \datamem.data_ram[12][17] ;
 wire \datamem.data_ram[12][18] ;
 wire \datamem.data_ram[12][19] ;
 wire \datamem.data_ram[12][1] ;
 wire \datamem.data_ram[12][20] ;
 wire \datamem.data_ram[12][21] ;
 wire \datamem.data_ram[12][22] ;
 wire \datamem.data_ram[12][23] ;
 wire \datamem.data_ram[12][24] ;
 wire \datamem.data_ram[12][25] ;
 wire \datamem.data_ram[12][26] ;
 wire \datamem.data_ram[12][27] ;
 wire \datamem.data_ram[12][28] ;
 wire \datamem.data_ram[12][29] ;
 wire \datamem.data_ram[12][2] ;
 wire \datamem.data_ram[12][30] ;
 wire \datamem.data_ram[12][31] ;
 wire \datamem.data_ram[12][3] ;
 wire \datamem.data_ram[12][4] ;
 wire \datamem.data_ram[12][5] ;
 wire \datamem.data_ram[12][6] ;
 wire \datamem.data_ram[12][7] ;
 wire \datamem.data_ram[12][8] ;
 wire \datamem.data_ram[12][9] ;
 wire \datamem.data_ram[13][0] ;
 wire \datamem.data_ram[13][10] ;
 wire \datamem.data_ram[13][11] ;
 wire \datamem.data_ram[13][12] ;
 wire \datamem.data_ram[13][13] ;
 wire \datamem.data_ram[13][14] ;
 wire \datamem.data_ram[13][15] ;
 wire \datamem.data_ram[13][16] ;
 wire \datamem.data_ram[13][17] ;
 wire \datamem.data_ram[13][18] ;
 wire \datamem.data_ram[13][19] ;
 wire \datamem.data_ram[13][1] ;
 wire \datamem.data_ram[13][20] ;
 wire \datamem.data_ram[13][21] ;
 wire \datamem.data_ram[13][22] ;
 wire \datamem.data_ram[13][23] ;
 wire \datamem.data_ram[13][24] ;
 wire \datamem.data_ram[13][25] ;
 wire \datamem.data_ram[13][26] ;
 wire \datamem.data_ram[13][27] ;
 wire \datamem.data_ram[13][28] ;
 wire \datamem.data_ram[13][29] ;
 wire \datamem.data_ram[13][2] ;
 wire \datamem.data_ram[13][30] ;
 wire \datamem.data_ram[13][31] ;
 wire \datamem.data_ram[13][3] ;
 wire \datamem.data_ram[13][4] ;
 wire \datamem.data_ram[13][5] ;
 wire \datamem.data_ram[13][6] ;
 wire \datamem.data_ram[13][7] ;
 wire \datamem.data_ram[13][8] ;
 wire \datamem.data_ram[13][9] ;
 wire \datamem.data_ram[14][0] ;
 wire \datamem.data_ram[14][10] ;
 wire \datamem.data_ram[14][11] ;
 wire \datamem.data_ram[14][12] ;
 wire \datamem.data_ram[14][13] ;
 wire \datamem.data_ram[14][14] ;
 wire \datamem.data_ram[14][15] ;
 wire \datamem.data_ram[14][16] ;
 wire \datamem.data_ram[14][17] ;
 wire \datamem.data_ram[14][18] ;
 wire \datamem.data_ram[14][19] ;
 wire \datamem.data_ram[14][1] ;
 wire \datamem.data_ram[14][20] ;
 wire \datamem.data_ram[14][21] ;
 wire \datamem.data_ram[14][22] ;
 wire \datamem.data_ram[14][23] ;
 wire \datamem.data_ram[14][24] ;
 wire \datamem.data_ram[14][25] ;
 wire \datamem.data_ram[14][26] ;
 wire \datamem.data_ram[14][27] ;
 wire \datamem.data_ram[14][28] ;
 wire \datamem.data_ram[14][29] ;
 wire \datamem.data_ram[14][2] ;
 wire \datamem.data_ram[14][30] ;
 wire \datamem.data_ram[14][31] ;
 wire \datamem.data_ram[14][3] ;
 wire \datamem.data_ram[14][4] ;
 wire \datamem.data_ram[14][5] ;
 wire \datamem.data_ram[14][6] ;
 wire \datamem.data_ram[14][7] ;
 wire \datamem.data_ram[14][8] ;
 wire \datamem.data_ram[14][9] ;
 wire \datamem.data_ram[15][0] ;
 wire \datamem.data_ram[15][10] ;
 wire \datamem.data_ram[15][11] ;
 wire \datamem.data_ram[15][12] ;
 wire \datamem.data_ram[15][13] ;
 wire \datamem.data_ram[15][14] ;
 wire \datamem.data_ram[15][15] ;
 wire \datamem.data_ram[15][16] ;
 wire \datamem.data_ram[15][17] ;
 wire \datamem.data_ram[15][18] ;
 wire \datamem.data_ram[15][19] ;
 wire \datamem.data_ram[15][1] ;
 wire \datamem.data_ram[15][20] ;
 wire \datamem.data_ram[15][21] ;
 wire \datamem.data_ram[15][22] ;
 wire \datamem.data_ram[15][23] ;
 wire \datamem.data_ram[15][24] ;
 wire \datamem.data_ram[15][25] ;
 wire \datamem.data_ram[15][26] ;
 wire \datamem.data_ram[15][27] ;
 wire \datamem.data_ram[15][28] ;
 wire \datamem.data_ram[15][29] ;
 wire \datamem.data_ram[15][2] ;
 wire \datamem.data_ram[15][30] ;
 wire \datamem.data_ram[15][31] ;
 wire \datamem.data_ram[15][3] ;
 wire \datamem.data_ram[15][4] ;
 wire \datamem.data_ram[15][5] ;
 wire \datamem.data_ram[15][6] ;
 wire \datamem.data_ram[15][7] ;
 wire \datamem.data_ram[15][8] ;
 wire \datamem.data_ram[15][9] ;
 wire \datamem.data_ram[16][0] ;
 wire \datamem.data_ram[16][10] ;
 wire \datamem.data_ram[16][11] ;
 wire \datamem.data_ram[16][12] ;
 wire \datamem.data_ram[16][13] ;
 wire \datamem.data_ram[16][14] ;
 wire \datamem.data_ram[16][15] ;
 wire \datamem.data_ram[16][16] ;
 wire \datamem.data_ram[16][17] ;
 wire \datamem.data_ram[16][18] ;
 wire \datamem.data_ram[16][19] ;
 wire \datamem.data_ram[16][1] ;
 wire \datamem.data_ram[16][20] ;
 wire \datamem.data_ram[16][21] ;
 wire \datamem.data_ram[16][22] ;
 wire \datamem.data_ram[16][23] ;
 wire \datamem.data_ram[16][24] ;
 wire \datamem.data_ram[16][25] ;
 wire \datamem.data_ram[16][26] ;
 wire \datamem.data_ram[16][27] ;
 wire \datamem.data_ram[16][28] ;
 wire \datamem.data_ram[16][29] ;
 wire \datamem.data_ram[16][2] ;
 wire \datamem.data_ram[16][30] ;
 wire \datamem.data_ram[16][31] ;
 wire \datamem.data_ram[16][3] ;
 wire \datamem.data_ram[16][4] ;
 wire \datamem.data_ram[16][5] ;
 wire \datamem.data_ram[16][6] ;
 wire \datamem.data_ram[16][7] ;
 wire \datamem.data_ram[16][8] ;
 wire \datamem.data_ram[16][9] ;
 wire \datamem.data_ram[17][0] ;
 wire \datamem.data_ram[17][10] ;
 wire \datamem.data_ram[17][11] ;
 wire \datamem.data_ram[17][12] ;
 wire \datamem.data_ram[17][13] ;
 wire \datamem.data_ram[17][14] ;
 wire \datamem.data_ram[17][15] ;
 wire \datamem.data_ram[17][16] ;
 wire \datamem.data_ram[17][17] ;
 wire \datamem.data_ram[17][18] ;
 wire \datamem.data_ram[17][19] ;
 wire \datamem.data_ram[17][1] ;
 wire \datamem.data_ram[17][20] ;
 wire \datamem.data_ram[17][21] ;
 wire \datamem.data_ram[17][22] ;
 wire \datamem.data_ram[17][23] ;
 wire \datamem.data_ram[17][24] ;
 wire \datamem.data_ram[17][25] ;
 wire \datamem.data_ram[17][26] ;
 wire \datamem.data_ram[17][27] ;
 wire \datamem.data_ram[17][28] ;
 wire \datamem.data_ram[17][29] ;
 wire \datamem.data_ram[17][2] ;
 wire \datamem.data_ram[17][30] ;
 wire \datamem.data_ram[17][31] ;
 wire \datamem.data_ram[17][3] ;
 wire \datamem.data_ram[17][4] ;
 wire \datamem.data_ram[17][5] ;
 wire \datamem.data_ram[17][6] ;
 wire \datamem.data_ram[17][7] ;
 wire \datamem.data_ram[17][8] ;
 wire \datamem.data_ram[17][9] ;
 wire \datamem.data_ram[18][0] ;
 wire \datamem.data_ram[18][10] ;
 wire \datamem.data_ram[18][11] ;
 wire \datamem.data_ram[18][12] ;
 wire \datamem.data_ram[18][13] ;
 wire \datamem.data_ram[18][14] ;
 wire \datamem.data_ram[18][15] ;
 wire \datamem.data_ram[18][16] ;
 wire \datamem.data_ram[18][17] ;
 wire \datamem.data_ram[18][18] ;
 wire \datamem.data_ram[18][19] ;
 wire \datamem.data_ram[18][1] ;
 wire \datamem.data_ram[18][20] ;
 wire \datamem.data_ram[18][21] ;
 wire \datamem.data_ram[18][22] ;
 wire \datamem.data_ram[18][23] ;
 wire \datamem.data_ram[18][24] ;
 wire \datamem.data_ram[18][25] ;
 wire \datamem.data_ram[18][26] ;
 wire \datamem.data_ram[18][27] ;
 wire \datamem.data_ram[18][28] ;
 wire \datamem.data_ram[18][29] ;
 wire \datamem.data_ram[18][2] ;
 wire \datamem.data_ram[18][30] ;
 wire \datamem.data_ram[18][31] ;
 wire \datamem.data_ram[18][3] ;
 wire \datamem.data_ram[18][4] ;
 wire \datamem.data_ram[18][5] ;
 wire \datamem.data_ram[18][6] ;
 wire \datamem.data_ram[18][7] ;
 wire \datamem.data_ram[18][8] ;
 wire \datamem.data_ram[18][9] ;
 wire \datamem.data_ram[19][0] ;
 wire \datamem.data_ram[19][10] ;
 wire \datamem.data_ram[19][11] ;
 wire \datamem.data_ram[19][12] ;
 wire \datamem.data_ram[19][13] ;
 wire \datamem.data_ram[19][14] ;
 wire \datamem.data_ram[19][15] ;
 wire \datamem.data_ram[19][16] ;
 wire \datamem.data_ram[19][17] ;
 wire \datamem.data_ram[19][18] ;
 wire \datamem.data_ram[19][19] ;
 wire \datamem.data_ram[19][1] ;
 wire \datamem.data_ram[19][20] ;
 wire \datamem.data_ram[19][21] ;
 wire \datamem.data_ram[19][22] ;
 wire \datamem.data_ram[19][23] ;
 wire \datamem.data_ram[19][24] ;
 wire \datamem.data_ram[19][25] ;
 wire \datamem.data_ram[19][26] ;
 wire \datamem.data_ram[19][27] ;
 wire \datamem.data_ram[19][28] ;
 wire \datamem.data_ram[19][29] ;
 wire \datamem.data_ram[19][2] ;
 wire \datamem.data_ram[19][30] ;
 wire \datamem.data_ram[19][31] ;
 wire \datamem.data_ram[19][3] ;
 wire \datamem.data_ram[19][4] ;
 wire \datamem.data_ram[19][5] ;
 wire \datamem.data_ram[19][6] ;
 wire \datamem.data_ram[19][7] ;
 wire \datamem.data_ram[19][8] ;
 wire \datamem.data_ram[19][9] ;
 wire \datamem.data_ram[1][0] ;
 wire \datamem.data_ram[1][10] ;
 wire \datamem.data_ram[1][11] ;
 wire \datamem.data_ram[1][12] ;
 wire \datamem.data_ram[1][13] ;
 wire \datamem.data_ram[1][14] ;
 wire \datamem.data_ram[1][15] ;
 wire \datamem.data_ram[1][16] ;
 wire \datamem.data_ram[1][17] ;
 wire \datamem.data_ram[1][18] ;
 wire \datamem.data_ram[1][19] ;
 wire \datamem.data_ram[1][1] ;
 wire \datamem.data_ram[1][20] ;
 wire \datamem.data_ram[1][21] ;
 wire \datamem.data_ram[1][22] ;
 wire \datamem.data_ram[1][23] ;
 wire \datamem.data_ram[1][24] ;
 wire \datamem.data_ram[1][25] ;
 wire \datamem.data_ram[1][26] ;
 wire \datamem.data_ram[1][27] ;
 wire \datamem.data_ram[1][28] ;
 wire \datamem.data_ram[1][29] ;
 wire \datamem.data_ram[1][2] ;
 wire \datamem.data_ram[1][30] ;
 wire \datamem.data_ram[1][31] ;
 wire \datamem.data_ram[1][3] ;
 wire \datamem.data_ram[1][4] ;
 wire \datamem.data_ram[1][5] ;
 wire \datamem.data_ram[1][6] ;
 wire \datamem.data_ram[1][7] ;
 wire \datamem.data_ram[1][8] ;
 wire \datamem.data_ram[1][9] ;
 wire \datamem.data_ram[20][0] ;
 wire \datamem.data_ram[20][10] ;
 wire \datamem.data_ram[20][11] ;
 wire \datamem.data_ram[20][12] ;
 wire \datamem.data_ram[20][13] ;
 wire \datamem.data_ram[20][14] ;
 wire \datamem.data_ram[20][15] ;
 wire \datamem.data_ram[20][16] ;
 wire \datamem.data_ram[20][17] ;
 wire \datamem.data_ram[20][18] ;
 wire \datamem.data_ram[20][19] ;
 wire \datamem.data_ram[20][1] ;
 wire \datamem.data_ram[20][20] ;
 wire \datamem.data_ram[20][21] ;
 wire \datamem.data_ram[20][22] ;
 wire \datamem.data_ram[20][23] ;
 wire \datamem.data_ram[20][24] ;
 wire \datamem.data_ram[20][25] ;
 wire \datamem.data_ram[20][26] ;
 wire \datamem.data_ram[20][27] ;
 wire \datamem.data_ram[20][28] ;
 wire \datamem.data_ram[20][29] ;
 wire \datamem.data_ram[20][2] ;
 wire \datamem.data_ram[20][30] ;
 wire \datamem.data_ram[20][31] ;
 wire \datamem.data_ram[20][3] ;
 wire \datamem.data_ram[20][4] ;
 wire \datamem.data_ram[20][5] ;
 wire \datamem.data_ram[20][6] ;
 wire \datamem.data_ram[20][7] ;
 wire \datamem.data_ram[20][8] ;
 wire \datamem.data_ram[20][9] ;
 wire \datamem.data_ram[21][0] ;
 wire \datamem.data_ram[21][10] ;
 wire \datamem.data_ram[21][11] ;
 wire \datamem.data_ram[21][12] ;
 wire \datamem.data_ram[21][13] ;
 wire \datamem.data_ram[21][14] ;
 wire \datamem.data_ram[21][15] ;
 wire \datamem.data_ram[21][16] ;
 wire \datamem.data_ram[21][17] ;
 wire \datamem.data_ram[21][18] ;
 wire \datamem.data_ram[21][19] ;
 wire \datamem.data_ram[21][1] ;
 wire \datamem.data_ram[21][20] ;
 wire \datamem.data_ram[21][21] ;
 wire \datamem.data_ram[21][22] ;
 wire \datamem.data_ram[21][23] ;
 wire \datamem.data_ram[21][24] ;
 wire \datamem.data_ram[21][25] ;
 wire \datamem.data_ram[21][26] ;
 wire \datamem.data_ram[21][27] ;
 wire \datamem.data_ram[21][28] ;
 wire \datamem.data_ram[21][29] ;
 wire \datamem.data_ram[21][2] ;
 wire \datamem.data_ram[21][30] ;
 wire \datamem.data_ram[21][31] ;
 wire \datamem.data_ram[21][3] ;
 wire \datamem.data_ram[21][4] ;
 wire \datamem.data_ram[21][5] ;
 wire \datamem.data_ram[21][6] ;
 wire \datamem.data_ram[21][7] ;
 wire \datamem.data_ram[21][8] ;
 wire \datamem.data_ram[21][9] ;
 wire \datamem.data_ram[22][0] ;
 wire \datamem.data_ram[22][10] ;
 wire \datamem.data_ram[22][11] ;
 wire \datamem.data_ram[22][12] ;
 wire \datamem.data_ram[22][13] ;
 wire \datamem.data_ram[22][14] ;
 wire \datamem.data_ram[22][15] ;
 wire \datamem.data_ram[22][16] ;
 wire \datamem.data_ram[22][17] ;
 wire \datamem.data_ram[22][18] ;
 wire \datamem.data_ram[22][19] ;
 wire \datamem.data_ram[22][1] ;
 wire \datamem.data_ram[22][20] ;
 wire \datamem.data_ram[22][21] ;
 wire \datamem.data_ram[22][22] ;
 wire \datamem.data_ram[22][23] ;
 wire \datamem.data_ram[22][24] ;
 wire \datamem.data_ram[22][25] ;
 wire \datamem.data_ram[22][26] ;
 wire \datamem.data_ram[22][27] ;
 wire \datamem.data_ram[22][28] ;
 wire \datamem.data_ram[22][29] ;
 wire \datamem.data_ram[22][2] ;
 wire \datamem.data_ram[22][30] ;
 wire \datamem.data_ram[22][31] ;
 wire \datamem.data_ram[22][3] ;
 wire \datamem.data_ram[22][4] ;
 wire \datamem.data_ram[22][5] ;
 wire \datamem.data_ram[22][6] ;
 wire \datamem.data_ram[22][7] ;
 wire \datamem.data_ram[22][8] ;
 wire \datamem.data_ram[22][9] ;
 wire \datamem.data_ram[23][0] ;
 wire \datamem.data_ram[23][10] ;
 wire \datamem.data_ram[23][11] ;
 wire \datamem.data_ram[23][12] ;
 wire \datamem.data_ram[23][13] ;
 wire \datamem.data_ram[23][14] ;
 wire \datamem.data_ram[23][15] ;
 wire \datamem.data_ram[23][16] ;
 wire \datamem.data_ram[23][17] ;
 wire \datamem.data_ram[23][18] ;
 wire \datamem.data_ram[23][19] ;
 wire \datamem.data_ram[23][1] ;
 wire \datamem.data_ram[23][20] ;
 wire \datamem.data_ram[23][21] ;
 wire \datamem.data_ram[23][22] ;
 wire \datamem.data_ram[23][23] ;
 wire \datamem.data_ram[23][24] ;
 wire \datamem.data_ram[23][25] ;
 wire \datamem.data_ram[23][26] ;
 wire \datamem.data_ram[23][27] ;
 wire \datamem.data_ram[23][28] ;
 wire \datamem.data_ram[23][29] ;
 wire \datamem.data_ram[23][2] ;
 wire \datamem.data_ram[23][30] ;
 wire \datamem.data_ram[23][31] ;
 wire \datamem.data_ram[23][3] ;
 wire \datamem.data_ram[23][4] ;
 wire \datamem.data_ram[23][5] ;
 wire \datamem.data_ram[23][6] ;
 wire \datamem.data_ram[23][7] ;
 wire \datamem.data_ram[23][8] ;
 wire \datamem.data_ram[23][9] ;
 wire \datamem.data_ram[24][0] ;
 wire \datamem.data_ram[24][10] ;
 wire \datamem.data_ram[24][11] ;
 wire \datamem.data_ram[24][12] ;
 wire \datamem.data_ram[24][13] ;
 wire \datamem.data_ram[24][14] ;
 wire \datamem.data_ram[24][15] ;
 wire \datamem.data_ram[24][16] ;
 wire \datamem.data_ram[24][17] ;
 wire \datamem.data_ram[24][18] ;
 wire \datamem.data_ram[24][19] ;
 wire \datamem.data_ram[24][1] ;
 wire \datamem.data_ram[24][20] ;
 wire \datamem.data_ram[24][21] ;
 wire \datamem.data_ram[24][22] ;
 wire \datamem.data_ram[24][23] ;
 wire \datamem.data_ram[24][24] ;
 wire \datamem.data_ram[24][25] ;
 wire \datamem.data_ram[24][26] ;
 wire \datamem.data_ram[24][27] ;
 wire \datamem.data_ram[24][28] ;
 wire \datamem.data_ram[24][29] ;
 wire \datamem.data_ram[24][2] ;
 wire \datamem.data_ram[24][30] ;
 wire \datamem.data_ram[24][31] ;
 wire \datamem.data_ram[24][3] ;
 wire \datamem.data_ram[24][4] ;
 wire \datamem.data_ram[24][5] ;
 wire \datamem.data_ram[24][6] ;
 wire \datamem.data_ram[24][7] ;
 wire \datamem.data_ram[24][8] ;
 wire \datamem.data_ram[24][9] ;
 wire \datamem.data_ram[25][0] ;
 wire \datamem.data_ram[25][10] ;
 wire \datamem.data_ram[25][11] ;
 wire \datamem.data_ram[25][12] ;
 wire \datamem.data_ram[25][13] ;
 wire \datamem.data_ram[25][14] ;
 wire \datamem.data_ram[25][15] ;
 wire \datamem.data_ram[25][16] ;
 wire \datamem.data_ram[25][17] ;
 wire \datamem.data_ram[25][18] ;
 wire \datamem.data_ram[25][19] ;
 wire \datamem.data_ram[25][1] ;
 wire \datamem.data_ram[25][20] ;
 wire \datamem.data_ram[25][21] ;
 wire \datamem.data_ram[25][22] ;
 wire \datamem.data_ram[25][23] ;
 wire \datamem.data_ram[25][24] ;
 wire \datamem.data_ram[25][25] ;
 wire \datamem.data_ram[25][26] ;
 wire \datamem.data_ram[25][27] ;
 wire \datamem.data_ram[25][28] ;
 wire \datamem.data_ram[25][29] ;
 wire \datamem.data_ram[25][2] ;
 wire \datamem.data_ram[25][30] ;
 wire \datamem.data_ram[25][31] ;
 wire \datamem.data_ram[25][3] ;
 wire \datamem.data_ram[25][4] ;
 wire \datamem.data_ram[25][5] ;
 wire \datamem.data_ram[25][6] ;
 wire \datamem.data_ram[25][7] ;
 wire \datamem.data_ram[25][8] ;
 wire \datamem.data_ram[25][9] ;
 wire \datamem.data_ram[26][0] ;
 wire \datamem.data_ram[26][10] ;
 wire \datamem.data_ram[26][11] ;
 wire \datamem.data_ram[26][12] ;
 wire \datamem.data_ram[26][13] ;
 wire \datamem.data_ram[26][14] ;
 wire \datamem.data_ram[26][15] ;
 wire \datamem.data_ram[26][16] ;
 wire \datamem.data_ram[26][17] ;
 wire \datamem.data_ram[26][18] ;
 wire \datamem.data_ram[26][19] ;
 wire \datamem.data_ram[26][1] ;
 wire \datamem.data_ram[26][20] ;
 wire \datamem.data_ram[26][21] ;
 wire \datamem.data_ram[26][22] ;
 wire \datamem.data_ram[26][23] ;
 wire \datamem.data_ram[26][24] ;
 wire \datamem.data_ram[26][25] ;
 wire \datamem.data_ram[26][26] ;
 wire \datamem.data_ram[26][27] ;
 wire \datamem.data_ram[26][28] ;
 wire \datamem.data_ram[26][29] ;
 wire \datamem.data_ram[26][2] ;
 wire \datamem.data_ram[26][30] ;
 wire \datamem.data_ram[26][31] ;
 wire \datamem.data_ram[26][3] ;
 wire \datamem.data_ram[26][4] ;
 wire \datamem.data_ram[26][5] ;
 wire \datamem.data_ram[26][6] ;
 wire \datamem.data_ram[26][7] ;
 wire \datamem.data_ram[26][8] ;
 wire \datamem.data_ram[26][9] ;
 wire \datamem.data_ram[27][0] ;
 wire \datamem.data_ram[27][10] ;
 wire \datamem.data_ram[27][11] ;
 wire \datamem.data_ram[27][12] ;
 wire \datamem.data_ram[27][13] ;
 wire \datamem.data_ram[27][14] ;
 wire \datamem.data_ram[27][15] ;
 wire \datamem.data_ram[27][16] ;
 wire \datamem.data_ram[27][17] ;
 wire \datamem.data_ram[27][18] ;
 wire \datamem.data_ram[27][19] ;
 wire \datamem.data_ram[27][1] ;
 wire \datamem.data_ram[27][20] ;
 wire \datamem.data_ram[27][21] ;
 wire \datamem.data_ram[27][22] ;
 wire \datamem.data_ram[27][23] ;
 wire \datamem.data_ram[27][24] ;
 wire \datamem.data_ram[27][25] ;
 wire \datamem.data_ram[27][26] ;
 wire \datamem.data_ram[27][27] ;
 wire \datamem.data_ram[27][28] ;
 wire \datamem.data_ram[27][29] ;
 wire \datamem.data_ram[27][2] ;
 wire \datamem.data_ram[27][30] ;
 wire \datamem.data_ram[27][31] ;
 wire \datamem.data_ram[27][3] ;
 wire \datamem.data_ram[27][4] ;
 wire \datamem.data_ram[27][5] ;
 wire \datamem.data_ram[27][6] ;
 wire \datamem.data_ram[27][7] ;
 wire \datamem.data_ram[27][8] ;
 wire \datamem.data_ram[27][9] ;
 wire \datamem.data_ram[28][0] ;
 wire \datamem.data_ram[28][10] ;
 wire \datamem.data_ram[28][11] ;
 wire \datamem.data_ram[28][12] ;
 wire \datamem.data_ram[28][13] ;
 wire \datamem.data_ram[28][14] ;
 wire \datamem.data_ram[28][15] ;
 wire \datamem.data_ram[28][16] ;
 wire \datamem.data_ram[28][17] ;
 wire \datamem.data_ram[28][18] ;
 wire \datamem.data_ram[28][19] ;
 wire \datamem.data_ram[28][1] ;
 wire \datamem.data_ram[28][20] ;
 wire \datamem.data_ram[28][21] ;
 wire \datamem.data_ram[28][22] ;
 wire \datamem.data_ram[28][23] ;
 wire \datamem.data_ram[28][24] ;
 wire \datamem.data_ram[28][25] ;
 wire \datamem.data_ram[28][26] ;
 wire \datamem.data_ram[28][27] ;
 wire \datamem.data_ram[28][28] ;
 wire \datamem.data_ram[28][29] ;
 wire \datamem.data_ram[28][2] ;
 wire \datamem.data_ram[28][30] ;
 wire \datamem.data_ram[28][31] ;
 wire \datamem.data_ram[28][3] ;
 wire \datamem.data_ram[28][4] ;
 wire \datamem.data_ram[28][5] ;
 wire \datamem.data_ram[28][6] ;
 wire \datamem.data_ram[28][7] ;
 wire \datamem.data_ram[28][8] ;
 wire \datamem.data_ram[28][9] ;
 wire \datamem.data_ram[29][0] ;
 wire \datamem.data_ram[29][10] ;
 wire \datamem.data_ram[29][11] ;
 wire \datamem.data_ram[29][12] ;
 wire \datamem.data_ram[29][13] ;
 wire \datamem.data_ram[29][14] ;
 wire \datamem.data_ram[29][15] ;
 wire \datamem.data_ram[29][16] ;
 wire \datamem.data_ram[29][17] ;
 wire \datamem.data_ram[29][18] ;
 wire \datamem.data_ram[29][19] ;
 wire \datamem.data_ram[29][1] ;
 wire \datamem.data_ram[29][20] ;
 wire \datamem.data_ram[29][21] ;
 wire \datamem.data_ram[29][22] ;
 wire \datamem.data_ram[29][23] ;
 wire \datamem.data_ram[29][24] ;
 wire \datamem.data_ram[29][25] ;
 wire \datamem.data_ram[29][26] ;
 wire \datamem.data_ram[29][27] ;
 wire \datamem.data_ram[29][28] ;
 wire \datamem.data_ram[29][29] ;
 wire \datamem.data_ram[29][2] ;
 wire \datamem.data_ram[29][30] ;
 wire \datamem.data_ram[29][31] ;
 wire \datamem.data_ram[29][3] ;
 wire \datamem.data_ram[29][4] ;
 wire \datamem.data_ram[29][5] ;
 wire \datamem.data_ram[29][6] ;
 wire \datamem.data_ram[29][7] ;
 wire \datamem.data_ram[29][8] ;
 wire \datamem.data_ram[29][9] ;
 wire \datamem.data_ram[2][0] ;
 wire \datamem.data_ram[2][10] ;
 wire \datamem.data_ram[2][11] ;
 wire \datamem.data_ram[2][12] ;
 wire \datamem.data_ram[2][13] ;
 wire \datamem.data_ram[2][14] ;
 wire \datamem.data_ram[2][15] ;
 wire \datamem.data_ram[2][16] ;
 wire \datamem.data_ram[2][17] ;
 wire \datamem.data_ram[2][18] ;
 wire \datamem.data_ram[2][19] ;
 wire \datamem.data_ram[2][1] ;
 wire \datamem.data_ram[2][20] ;
 wire \datamem.data_ram[2][21] ;
 wire \datamem.data_ram[2][22] ;
 wire \datamem.data_ram[2][23] ;
 wire \datamem.data_ram[2][24] ;
 wire \datamem.data_ram[2][25] ;
 wire \datamem.data_ram[2][26] ;
 wire \datamem.data_ram[2][27] ;
 wire \datamem.data_ram[2][28] ;
 wire \datamem.data_ram[2][29] ;
 wire \datamem.data_ram[2][2] ;
 wire \datamem.data_ram[2][30] ;
 wire \datamem.data_ram[2][31] ;
 wire \datamem.data_ram[2][3] ;
 wire \datamem.data_ram[2][4] ;
 wire \datamem.data_ram[2][5] ;
 wire \datamem.data_ram[2][6] ;
 wire \datamem.data_ram[2][7] ;
 wire \datamem.data_ram[2][8] ;
 wire \datamem.data_ram[2][9] ;
 wire \datamem.data_ram[30][0] ;
 wire \datamem.data_ram[30][10] ;
 wire \datamem.data_ram[30][11] ;
 wire \datamem.data_ram[30][12] ;
 wire \datamem.data_ram[30][13] ;
 wire \datamem.data_ram[30][14] ;
 wire \datamem.data_ram[30][15] ;
 wire \datamem.data_ram[30][16] ;
 wire \datamem.data_ram[30][17] ;
 wire \datamem.data_ram[30][18] ;
 wire \datamem.data_ram[30][19] ;
 wire \datamem.data_ram[30][1] ;
 wire \datamem.data_ram[30][20] ;
 wire \datamem.data_ram[30][21] ;
 wire \datamem.data_ram[30][22] ;
 wire \datamem.data_ram[30][23] ;
 wire \datamem.data_ram[30][24] ;
 wire \datamem.data_ram[30][25] ;
 wire \datamem.data_ram[30][26] ;
 wire \datamem.data_ram[30][27] ;
 wire \datamem.data_ram[30][28] ;
 wire \datamem.data_ram[30][29] ;
 wire \datamem.data_ram[30][2] ;
 wire \datamem.data_ram[30][30] ;
 wire \datamem.data_ram[30][31] ;
 wire \datamem.data_ram[30][3] ;
 wire \datamem.data_ram[30][4] ;
 wire \datamem.data_ram[30][5] ;
 wire \datamem.data_ram[30][6] ;
 wire \datamem.data_ram[30][7] ;
 wire \datamem.data_ram[30][8] ;
 wire \datamem.data_ram[30][9] ;
 wire \datamem.data_ram[31][0] ;
 wire \datamem.data_ram[31][10] ;
 wire \datamem.data_ram[31][11] ;
 wire \datamem.data_ram[31][12] ;
 wire \datamem.data_ram[31][13] ;
 wire \datamem.data_ram[31][14] ;
 wire \datamem.data_ram[31][15] ;
 wire \datamem.data_ram[31][16] ;
 wire \datamem.data_ram[31][17] ;
 wire \datamem.data_ram[31][18] ;
 wire \datamem.data_ram[31][19] ;
 wire \datamem.data_ram[31][1] ;
 wire \datamem.data_ram[31][20] ;
 wire \datamem.data_ram[31][21] ;
 wire \datamem.data_ram[31][22] ;
 wire \datamem.data_ram[31][23] ;
 wire \datamem.data_ram[31][24] ;
 wire \datamem.data_ram[31][25] ;
 wire \datamem.data_ram[31][26] ;
 wire \datamem.data_ram[31][27] ;
 wire \datamem.data_ram[31][28] ;
 wire \datamem.data_ram[31][29] ;
 wire \datamem.data_ram[31][2] ;
 wire \datamem.data_ram[31][30] ;
 wire \datamem.data_ram[31][31] ;
 wire \datamem.data_ram[31][3] ;
 wire \datamem.data_ram[31][4] ;
 wire \datamem.data_ram[31][5] ;
 wire \datamem.data_ram[31][6] ;
 wire \datamem.data_ram[31][7] ;
 wire \datamem.data_ram[31][8] ;
 wire \datamem.data_ram[31][9] ;
 wire \datamem.data_ram[32][0] ;
 wire \datamem.data_ram[32][10] ;
 wire \datamem.data_ram[32][11] ;
 wire \datamem.data_ram[32][12] ;
 wire \datamem.data_ram[32][13] ;
 wire \datamem.data_ram[32][14] ;
 wire \datamem.data_ram[32][15] ;
 wire \datamem.data_ram[32][16] ;
 wire \datamem.data_ram[32][17] ;
 wire \datamem.data_ram[32][18] ;
 wire \datamem.data_ram[32][19] ;
 wire \datamem.data_ram[32][1] ;
 wire \datamem.data_ram[32][20] ;
 wire \datamem.data_ram[32][21] ;
 wire \datamem.data_ram[32][22] ;
 wire \datamem.data_ram[32][23] ;
 wire \datamem.data_ram[32][24] ;
 wire \datamem.data_ram[32][25] ;
 wire \datamem.data_ram[32][26] ;
 wire \datamem.data_ram[32][27] ;
 wire \datamem.data_ram[32][28] ;
 wire \datamem.data_ram[32][29] ;
 wire \datamem.data_ram[32][2] ;
 wire \datamem.data_ram[32][30] ;
 wire \datamem.data_ram[32][31] ;
 wire \datamem.data_ram[32][3] ;
 wire \datamem.data_ram[32][4] ;
 wire \datamem.data_ram[32][5] ;
 wire \datamem.data_ram[32][6] ;
 wire \datamem.data_ram[32][7] ;
 wire \datamem.data_ram[32][8] ;
 wire \datamem.data_ram[32][9] ;
 wire \datamem.data_ram[33][0] ;
 wire \datamem.data_ram[33][10] ;
 wire \datamem.data_ram[33][11] ;
 wire \datamem.data_ram[33][12] ;
 wire \datamem.data_ram[33][13] ;
 wire \datamem.data_ram[33][14] ;
 wire \datamem.data_ram[33][15] ;
 wire \datamem.data_ram[33][16] ;
 wire \datamem.data_ram[33][17] ;
 wire \datamem.data_ram[33][18] ;
 wire \datamem.data_ram[33][19] ;
 wire \datamem.data_ram[33][1] ;
 wire \datamem.data_ram[33][20] ;
 wire \datamem.data_ram[33][21] ;
 wire \datamem.data_ram[33][22] ;
 wire \datamem.data_ram[33][23] ;
 wire \datamem.data_ram[33][24] ;
 wire \datamem.data_ram[33][25] ;
 wire \datamem.data_ram[33][26] ;
 wire \datamem.data_ram[33][27] ;
 wire \datamem.data_ram[33][28] ;
 wire \datamem.data_ram[33][29] ;
 wire \datamem.data_ram[33][2] ;
 wire \datamem.data_ram[33][30] ;
 wire \datamem.data_ram[33][31] ;
 wire \datamem.data_ram[33][3] ;
 wire \datamem.data_ram[33][4] ;
 wire \datamem.data_ram[33][5] ;
 wire \datamem.data_ram[33][6] ;
 wire \datamem.data_ram[33][7] ;
 wire \datamem.data_ram[33][8] ;
 wire \datamem.data_ram[33][9] ;
 wire \datamem.data_ram[34][0] ;
 wire \datamem.data_ram[34][10] ;
 wire \datamem.data_ram[34][11] ;
 wire \datamem.data_ram[34][12] ;
 wire \datamem.data_ram[34][13] ;
 wire \datamem.data_ram[34][14] ;
 wire \datamem.data_ram[34][15] ;
 wire \datamem.data_ram[34][16] ;
 wire \datamem.data_ram[34][17] ;
 wire \datamem.data_ram[34][18] ;
 wire \datamem.data_ram[34][19] ;
 wire \datamem.data_ram[34][1] ;
 wire \datamem.data_ram[34][20] ;
 wire \datamem.data_ram[34][21] ;
 wire \datamem.data_ram[34][22] ;
 wire \datamem.data_ram[34][23] ;
 wire \datamem.data_ram[34][24] ;
 wire \datamem.data_ram[34][25] ;
 wire \datamem.data_ram[34][26] ;
 wire \datamem.data_ram[34][27] ;
 wire \datamem.data_ram[34][28] ;
 wire \datamem.data_ram[34][29] ;
 wire \datamem.data_ram[34][2] ;
 wire \datamem.data_ram[34][30] ;
 wire \datamem.data_ram[34][31] ;
 wire \datamem.data_ram[34][3] ;
 wire \datamem.data_ram[34][4] ;
 wire \datamem.data_ram[34][5] ;
 wire \datamem.data_ram[34][6] ;
 wire \datamem.data_ram[34][7] ;
 wire \datamem.data_ram[34][8] ;
 wire \datamem.data_ram[34][9] ;
 wire \datamem.data_ram[35][0] ;
 wire \datamem.data_ram[35][10] ;
 wire \datamem.data_ram[35][11] ;
 wire \datamem.data_ram[35][12] ;
 wire \datamem.data_ram[35][13] ;
 wire \datamem.data_ram[35][14] ;
 wire \datamem.data_ram[35][15] ;
 wire \datamem.data_ram[35][16] ;
 wire \datamem.data_ram[35][17] ;
 wire \datamem.data_ram[35][18] ;
 wire \datamem.data_ram[35][19] ;
 wire \datamem.data_ram[35][1] ;
 wire \datamem.data_ram[35][20] ;
 wire \datamem.data_ram[35][21] ;
 wire \datamem.data_ram[35][22] ;
 wire \datamem.data_ram[35][23] ;
 wire \datamem.data_ram[35][24] ;
 wire \datamem.data_ram[35][25] ;
 wire \datamem.data_ram[35][26] ;
 wire \datamem.data_ram[35][27] ;
 wire \datamem.data_ram[35][28] ;
 wire \datamem.data_ram[35][29] ;
 wire \datamem.data_ram[35][2] ;
 wire \datamem.data_ram[35][30] ;
 wire \datamem.data_ram[35][31] ;
 wire \datamem.data_ram[35][3] ;
 wire \datamem.data_ram[35][4] ;
 wire \datamem.data_ram[35][5] ;
 wire \datamem.data_ram[35][6] ;
 wire \datamem.data_ram[35][7] ;
 wire \datamem.data_ram[35][8] ;
 wire \datamem.data_ram[35][9] ;
 wire \datamem.data_ram[36][0] ;
 wire \datamem.data_ram[36][10] ;
 wire \datamem.data_ram[36][11] ;
 wire \datamem.data_ram[36][12] ;
 wire \datamem.data_ram[36][13] ;
 wire \datamem.data_ram[36][14] ;
 wire \datamem.data_ram[36][15] ;
 wire \datamem.data_ram[36][16] ;
 wire \datamem.data_ram[36][17] ;
 wire \datamem.data_ram[36][18] ;
 wire \datamem.data_ram[36][19] ;
 wire \datamem.data_ram[36][1] ;
 wire \datamem.data_ram[36][20] ;
 wire \datamem.data_ram[36][21] ;
 wire \datamem.data_ram[36][22] ;
 wire \datamem.data_ram[36][23] ;
 wire \datamem.data_ram[36][24] ;
 wire \datamem.data_ram[36][25] ;
 wire \datamem.data_ram[36][26] ;
 wire \datamem.data_ram[36][27] ;
 wire \datamem.data_ram[36][28] ;
 wire \datamem.data_ram[36][29] ;
 wire \datamem.data_ram[36][2] ;
 wire \datamem.data_ram[36][30] ;
 wire \datamem.data_ram[36][31] ;
 wire \datamem.data_ram[36][3] ;
 wire \datamem.data_ram[36][4] ;
 wire \datamem.data_ram[36][5] ;
 wire \datamem.data_ram[36][6] ;
 wire \datamem.data_ram[36][7] ;
 wire \datamem.data_ram[36][8] ;
 wire \datamem.data_ram[36][9] ;
 wire \datamem.data_ram[37][0] ;
 wire \datamem.data_ram[37][10] ;
 wire \datamem.data_ram[37][11] ;
 wire \datamem.data_ram[37][12] ;
 wire \datamem.data_ram[37][13] ;
 wire \datamem.data_ram[37][14] ;
 wire \datamem.data_ram[37][15] ;
 wire \datamem.data_ram[37][16] ;
 wire \datamem.data_ram[37][17] ;
 wire \datamem.data_ram[37][18] ;
 wire \datamem.data_ram[37][19] ;
 wire \datamem.data_ram[37][1] ;
 wire \datamem.data_ram[37][20] ;
 wire \datamem.data_ram[37][21] ;
 wire \datamem.data_ram[37][22] ;
 wire \datamem.data_ram[37][23] ;
 wire \datamem.data_ram[37][24] ;
 wire \datamem.data_ram[37][25] ;
 wire \datamem.data_ram[37][26] ;
 wire \datamem.data_ram[37][27] ;
 wire \datamem.data_ram[37][28] ;
 wire \datamem.data_ram[37][29] ;
 wire \datamem.data_ram[37][2] ;
 wire \datamem.data_ram[37][30] ;
 wire \datamem.data_ram[37][31] ;
 wire \datamem.data_ram[37][3] ;
 wire \datamem.data_ram[37][4] ;
 wire \datamem.data_ram[37][5] ;
 wire \datamem.data_ram[37][6] ;
 wire \datamem.data_ram[37][7] ;
 wire \datamem.data_ram[37][8] ;
 wire \datamem.data_ram[37][9] ;
 wire \datamem.data_ram[38][0] ;
 wire \datamem.data_ram[38][10] ;
 wire \datamem.data_ram[38][11] ;
 wire \datamem.data_ram[38][12] ;
 wire \datamem.data_ram[38][13] ;
 wire \datamem.data_ram[38][14] ;
 wire \datamem.data_ram[38][15] ;
 wire \datamem.data_ram[38][16] ;
 wire \datamem.data_ram[38][17] ;
 wire \datamem.data_ram[38][18] ;
 wire \datamem.data_ram[38][19] ;
 wire \datamem.data_ram[38][1] ;
 wire \datamem.data_ram[38][20] ;
 wire \datamem.data_ram[38][21] ;
 wire \datamem.data_ram[38][22] ;
 wire \datamem.data_ram[38][23] ;
 wire \datamem.data_ram[38][24] ;
 wire \datamem.data_ram[38][25] ;
 wire \datamem.data_ram[38][26] ;
 wire \datamem.data_ram[38][27] ;
 wire \datamem.data_ram[38][28] ;
 wire \datamem.data_ram[38][29] ;
 wire \datamem.data_ram[38][2] ;
 wire \datamem.data_ram[38][30] ;
 wire \datamem.data_ram[38][31] ;
 wire \datamem.data_ram[38][3] ;
 wire \datamem.data_ram[38][4] ;
 wire \datamem.data_ram[38][5] ;
 wire \datamem.data_ram[38][6] ;
 wire \datamem.data_ram[38][7] ;
 wire \datamem.data_ram[38][8] ;
 wire \datamem.data_ram[38][9] ;
 wire \datamem.data_ram[39][0] ;
 wire \datamem.data_ram[39][10] ;
 wire \datamem.data_ram[39][11] ;
 wire \datamem.data_ram[39][12] ;
 wire \datamem.data_ram[39][13] ;
 wire \datamem.data_ram[39][14] ;
 wire \datamem.data_ram[39][15] ;
 wire \datamem.data_ram[39][16] ;
 wire \datamem.data_ram[39][17] ;
 wire \datamem.data_ram[39][18] ;
 wire \datamem.data_ram[39][19] ;
 wire \datamem.data_ram[39][1] ;
 wire \datamem.data_ram[39][20] ;
 wire \datamem.data_ram[39][21] ;
 wire \datamem.data_ram[39][22] ;
 wire \datamem.data_ram[39][23] ;
 wire \datamem.data_ram[39][24] ;
 wire \datamem.data_ram[39][25] ;
 wire \datamem.data_ram[39][26] ;
 wire \datamem.data_ram[39][27] ;
 wire \datamem.data_ram[39][28] ;
 wire \datamem.data_ram[39][29] ;
 wire \datamem.data_ram[39][2] ;
 wire \datamem.data_ram[39][30] ;
 wire \datamem.data_ram[39][31] ;
 wire \datamem.data_ram[39][3] ;
 wire \datamem.data_ram[39][4] ;
 wire \datamem.data_ram[39][5] ;
 wire \datamem.data_ram[39][6] ;
 wire \datamem.data_ram[39][7] ;
 wire \datamem.data_ram[39][8] ;
 wire \datamem.data_ram[39][9] ;
 wire \datamem.data_ram[3][0] ;
 wire \datamem.data_ram[3][10] ;
 wire \datamem.data_ram[3][11] ;
 wire \datamem.data_ram[3][12] ;
 wire \datamem.data_ram[3][13] ;
 wire \datamem.data_ram[3][14] ;
 wire \datamem.data_ram[3][15] ;
 wire \datamem.data_ram[3][16] ;
 wire \datamem.data_ram[3][17] ;
 wire \datamem.data_ram[3][18] ;
 wire \datamem.data_ram[3][19] ;
 wire \datamem.data_ram[3][1] ;
 wire \datamem.data_ram[3][20] ;
 wire \datamem.data_ram[3][21] ;
 wire \datamem.data_ram[3][22] ;
 wire \datamem.data_ram[3][23] ;
 wire \datamem.data_ram[3][24] ;
 wire \datamem.data_ram[3][25] ;
 wire \datamem.data_ram[3][26] ;
 wire \datamem.data_ram[3][27] ;
 wire \datamem.data_ram[3][28] ;
 wire \datamem.data_ram[3][29] ;
 wire \datamem.data_ram[3][2] ;
 wire \datamem.data_ram[3][30] ;
 wire \datamem.data_ram[3][31] ;
 wire \datamem.data_ram[3][3] ;
 wire \datamem.data_ram[3][4] ;
 wire \datamem.data_ram[3][5] ;
 wire \datamem.data_ram[3][6] ;
 wire \datamem.data_ram[3][7] ;
 wire \datamem.data_ram[3][8] ;
 wire \datamem.data_ram[3][9] ;
 wire \datamem.data_ram[40][0] ;
 wire \datamem.data_ram[40][10] ;
 wire \datamem.data_ram[40][11] ;
 wire \datamem.data_ram[40][12] ;
 wire \datamem.data_ram[40][13] ;
 wire \datamem.data_ram[40][14] ;
 wire \datamem.data_ram[40][15] ;
 wire \datamem.data_ram[40][16] ;
 wire \datamem.data_ram[40][17] ;
 wire \datamem.data_ram[40][18] ;
 wire \datamem.data_ram[40][19] ;
 wire \datamem.data_ram[40][1] ;
 wire \datamem.data_ram[40][20] ;
 wire \datamem.data_ram[40][21] ;
 wire \datamem.data_ram[40][22] ;
 wire \datamem.data_ram[40][23] ;
 wire \datamem.data_ram[40][24] ;
 wire \datamem.data_ram[40][25] ;
 wire \datamem.data_ram[40][26] ;
 wire \datamem.data_ram[40][27] ;
 wire \datamem.data_ram[40][28] ;
 wire \datamem.data_ram[40][29] ;
 wire \datamem.data_ram[40][2] ;
 wire \datamem.data_ram[40][30] ;
 wire \datamem.data_ram[40][31] ;
 wire \datamem.data_ram[40][3] ;
 wire \datamem.data_ram[40][4] ;
 wire \datamem.data_ram[40][5] ;
 wire \datamem.data_ram[40][6] ;
 wire \datamem.data_ram[40][7] ;
 wire \datamem.data_ram[40][8] ;
 wire \datamem.data_ram[40][9] ;
 wire \datamem.data_ram[41][0] ;
 wire \datamem.data_ram[41][10] ;
 wire \datamem.data_ram[41][11] ;
 wire \datamem.data_ram[41][12] ;
 wire \datamem.data_ram[41][13] ;
 wire \datamem.data_ram[41][14] ;
 wire \datamem.data_ram[41][15] ;
 wire \datamem.data_ram[41][16] ;
 wire \datamem.data_ram[41][17] ;
 wire \datamem.data_ram[41][18] ;
 wire \datamem.data_ram[41][19] ;
 wire \datamem.data_ram[41][1] ;
 wire \datamem.data_ram[41][20] ;
 wire \datamem.data_ram[41][21] ;
 wire \datamem.data_ram[41][22] ;
 wire \datamem.data_ram[41][23] ;
 wire \datamem.data_ram[41][24] ;
 wire \datamem.data_ram[41][25] ;
 wire \datamem.data_ram[41][26] ;
 wire \datamem.data_ram[41][27] ;
 wire \datamem.data_ram[41][28] ;
 wire \datamem.data_ram[41][29] ;
 wire \datamem.data_ram[41][2] ;
 wire \datamem.data_ram[41][30] ;
 wire \datamem.data_ram[41][31] ;
 wire \datamem.data_ram[41][3] ;
 wire \datamem.data_ram[41][4] ;
 wire \datamem.data_ram[41][5] ;
 wire \datamem.data_ram[41][6] ;
 wire \datamem.data_ram[41][7] ;
 wire \datamem.data_ram[41][8] ;
 wire \datamem.data_ram[41][9] ;
 wire \datamem.data_ram[42][0] ;
 wire \datamem.data_ram[42][10] ;
 wire \datamem.data_ram[42][11] ;
 wire \datamem.data_ram[42][12] ;
 wire \datamem.data_ram[42][13] ;
 wire \datamem.data_ram[42][14] ;
 wire \datamem.data_ram[42][15] ;
 wire \datamem.data_ram[42][16] ;
 wire \datamem.data_ram[42][17] ;
 wire \datamem.data_ram[42][18] ;
 wire \datamem.data_ram[42][19] ;
 wire \datamem.data_ram[42][1] ;
 wire \datamem.data_ram[42][20] ;
 wire \datamem.data_ram[42][21] ;
 wire \datamem.data_ram[42][22] ;
 wire \datamem.data_ram[42][23] ;
 wire \datamem.data_ram[42][24] ;
 wire \datamem.data_ram[42][25] ;
 wire \datamem.data_ram[42][26] ;
 wire \datamem.data_ram[42][27] ;
 wire \datamem.data_ram[42][28] ;
 wire \datamem.data_ram[42][29] ;
 wire \datamem.data_ram[42][2] ;
 wire \datamem.data_ram[42][30] ;
 wire \datamem.data_ram[42][31] ;
 wire \datamem.data_ram[42][3] ;
 wire \datamem.data_ram[42][4] ;
 wire \datamem.data_ram[42][5] ;
 wire \datamem.data_ram[42][6] ;
 wire \datamem.data_ram[42][7] ;
 wire \datamem.data_ram[42][8] ;
 wire \datamem.data_ram[42][9] ;
 wire \datamem.data_ram[43][0] ;
 wire \datamem.data_ram[43][10] ;
 wire \datamem.data_ram[43][11] ;
 wire \datamem.data_ram[43][12] ;
 wire \datamem.data_ram[43][13] ;
 wire \datamem.data_ram[43][14] ;
 wire \datamem.data_ram[43][15] ;
 wire \datamem.data_ram[43][16] ;
 wire \datamem.data_ram[43][17] ;
 wire \datamem.data_ram[43][18] ;
 wire \datamem.data_ram[43][19] ;
 wire \datamem.data_ram[43][1] ;
 wire \datamem.data_ram[43][20] ;
 wire \datamem.data_ram[43][21] ;
 wire \datamem.data_ram[43][22] ;
 wire \datamem.data_ram[43][23] ;
 wire \datamem.data_ram[43][24] ;
 wire \datamem.data_ram[43][25] ;
 wire \datamem.data_ram[43][26] ;
 wire \datamem.data_ram[43][27] ;
 wire \datamem.data_ram[43][28] ;
 wire \datamem.data_ram[43][29] ;
 wire \datamem.data_ram[43][2] ;
 wire \datamem.data_ram[43][30] ;
 wire \datamem.data_ram[43][31] ;
 wire \datamem.data_ram[43][3] ;
 wire \datamem.data_ram[43][4] ;
 wire \datamem.data_ram[43][5] ;
 wire \datamem.data_ram[43][6] ;
 wire \datamem.data_ram[43][7] ;
 wire \datamem.data_ram[43][8] ;
 wire \datamem.data_ram[43][9] ;
 wire \datamem.data_ram[44][0] ;
 wire \datamem.data_ram[44][10] ;
 wire \datamem.data_ram[44][11] ;
 wire \datamem.data_ram[44][12] ;
 wire \datamem.data_ram[44][13] ;
 wire \datamem.data_ram[44][14] ;
 wire \datamem.data_ram[44][15] ;
 wire \datamem.data_ram[44][16] ;
 wire \datamem.data_ram[44][17] ;
 wire \datamem.data_ram[44][18] ;
 wire \datamem.data_ram[44][19] ;
 wire \datamem.data_ram[44][1] ;
 wire \datamem.data_ram[44][20] ;
 wire \datamem.data_ram[44][21] ;
 wire \datamem.data_ram[44][22] ;
 wire \datamem.data_ram[44][23] ;
 wire \datamem.data_ram[44][24] ;
 wire \datamem.data_ram[44][25] ;
 wire \datamem.data_ram[44][26] ;
 wire \datamem.data_ram[44][27] ;
 wire \datamem.data_ram[44][28] ;
 wire \datamem.data_ram[44][29] ;
 wire \datamem.data_ram[44][2] ;
 wire \datamem.data_ram[44][30] ;
 wire \datamem.data_ram[44][31] ;
 wire \datamem.data_ram[44][3] ;
 wire \datamem.data_ram[44][4] ;
 wire \datamem.data_ram[44][5] ;
 wire \datamem.data_ram[44][6] ;
 wire \datamem.data_ram[44][7] ;
 wire \datamem.data_ram[44][8] ;
 wire \datamem.data_ram[44][9] ;
 wire \datamem.data_ram[45][0] ;
 wire \datamem.data_ram[45][10] ;
 wire \datamem.data_ram[45][11] ;
 wire \datamem.data_ram[45][12] ;
 wire \datamem.data_ram[45][13] ;
 wire \datamem.data_ram[45][14] ;
 wire \datamem.data_ram[45][15] ;
 wire \datamem.data_ram[45][16] ;
 wire \datamem.data_ram[45][17] ;
 wire \datamem.data_ram[45][18] ;
 wire \datamem.data_ram[45][19] ;
 wire \datamem.data_ram[45][1] ;
 wire \datamem.data_ram[45][20] ;
 wire \datamem.data_ram[45][21] ;
 wire \datamem.data_ram[45][22] ;
 wire \datamem.data_ram[45][23] ;
 wire \datamem.data_ram[45][24] ;
 wire \datamem.data_ram[45][25] ;
 wire \datamem.data_ram[45][26] ;
 wire \datamem.data_ram[45][27] ;
 wire \datamem.data_ram[45][28] ;
 wire \datamem.data_ram[45][29] ;
 wire \datamem.data_ram[45][2] ;
 wire \datamem.data_ram[45][30] ;
 wire \datamem.data_ram[45][31] ;
 wire \datamem.data_ram[45][3] ;
 wire \datamem.data_ram[45][4] ;
 wire \datamem.data_ram[45][5] ;
 wire \datamem.data_ram[45][6] ;
 wire \datamem.data_ram[45][7] ;
 wire \datamem.data_ram[45][8] ;
 wire \datamem.data_ram[45][9] ;
 wire \datamem.data_ram[46][0] ;
 wire \datamem.data_ram[46][10] ;
 wire \datamem.data_ram[46][11] ;
 wire \datamem.data_ram[46][12] ;
 wire \datamem.data_ram[46][13] ;
 wire \datamem.data_ram[46][14] ;
 wire \datamem.data_ram[46][15] ;
 wire \datamem.data_ram[46][16] ;
 wire \datamem.data_ram[46][17] ;
 wire \datamem.data_ram[46][18] ;
 wire \datamem.data_ram[46][19] ;
 wire \datamem.data_ram[46][1] ;
 wire \datamem.data_ram[46][20] ;
 wire \datamem.data_ram[46][21] ;
 wire \datamem.data_ram[46][22] ;
 wire \datamem.data_ram[46][23] ;
 wire \datamem.data_ram[46][24] ;
 wire \datamem.data_ram[46][25] ;
 wire \datamem.data_ram[46][26] ;
 wire \datamem.data_ram[46][27] ;
 wire \datamem.data_ram[46][28] ;
 wire \datamem.data_ram[46][29] ;
 wire \datamem.data_ram[46][2] ;
 wire \datamem.data_ram[46][30] ;
 wire \datamem.data_ram[46][31] ;
 wire \datamem.data_ram[46][3] ;
 wire \datamem.data_ram[46][4] ;
 wire \datamem.data_ram[46][5] ;
 wire \datamem.data_ram[46][6] ;
 wire \datamem.data_ram[46][7] ;
 wire \datamem.data_ram[46][8] ;
 wire \datamem.data_ram[46][9] ;
 wire \datamem.data_ram[47][0] ;
 wire \datamem.data_ram[47][10] ;
 wire \datamem.data_ram[47][11] ;
 wire \datamem.data_ram[47][12] ;
 wire \datamem.data_ram[47][13] ;
 wire \datamem.data_ram[47][14] ;
 wire \datamem.data_ram[47][15] ;
 wire \datamem.data_ram[47][16] ;
 wire \datamem.data_ram[47][17] ;
 wire \datamem.data_ram[47][18] ;
 wire \datamem.data_ram[47][19] ;
 wire \datamem.data_ram[47][1] ;
 wire \datamem.data_ram[47][20] ;
 wire \datamem.data_ram[47][21] ;
 wire \datamem.data_ram[47][22] ;
 wire \datamem.data_ram[47][23] ;
 wire \datamem.data_ram[47][24] ;
 wire \datamem.data_ram[47][25] ;
 wire \datamem.data_ram[47][26] ;
 wire \datamem.data_ram[47][27] ;
 wire \datamem.data_ram[47][28] ;
 wire \datamem.data_ram[47][29] ;
 wire \datamem.data_ram[47][2] ;
 wire \datamem.data_ram[47][30] ;
 wire \datamem.data_ram[47][31] ;
 wire \datamem.data_ram[47][3] ;
 wire \datamem.data_ram[47][4] ;
 wire \datamem.data_ram[47][5] ;
 wire \datamem.data_ram[47][6] ;
 wire \datamem.data_ram[47][7] ;
 wire \datamem.data_ram[47][8] ;
 wire \datamem.data_ram[47][9] ;
 wire \datamem.data_ram[48][0] ;
 wire \datamem.data_ram[48][10] ;
 wire \datamem.data_ram[48][11] ;
 wire \datamem.data_ram[48][12] ;
 wire \datamem.data_ram[48][13] ;
 wire \datamem.data_ram[48][14] ;
 wire \datamem.data_ram[48][15] ;
 wire \datamem.data_ram[48][16] ;
 wire \datamem.data_ram[48][17] ;
 wire \datamem.data_ram[48][18] ;
 wire \datamem.data_ram[48][19] ;
 wire \datamem.data_ram[48][1] ;
 wire \datamem.data_ram[48][20] ;
 wire \datamem.data_ram[48][21] ;
 wire \datamem.data_ram[48][22] ;
 wire \datamem.data_ram[48][23] ;
 wire \datamem.data_ram[48][24] ;
 wire \datamem.data_ram[48][25] ;
 wire \datamem.data_ram[48][26] ;
 wire \datamem.data_ram[48][27] ;
 wire \datamem.data_ram[48][28] ;
 wire \datamem.data_ram[48][29] ;
 wire \datamem.data_ram[48][2] ;
 wire \datamem.data_ram[48][30] ;
 wire \datamem.data_ram[48][31] ;
 wire \datamem.data_ram[48][3] ;
 wire \datamem.data_ram[48][4] ;
 wire \datamem.data_ram[48][5] ;
 wire \datamem.data_ram[48][6] ;
 wire \datamem.data_ram[48][7] ;
 wire \datamem.data_ram[48][8] ;
 wire \datamem.data_ram[48][9] ;
 wire \datamem.data_ram[49][0] ;
 wire \datamem.data_ram[49][10] ;
 wire \datamem.data_ram[49][11] ;
 wire \datamem.data_ram[49][12] ;
 wire \datamem.data_ram[49][13] ;
 wire \datamem.data_ram[49][14] ;
 wire \datamem.data_ram[49][15] ;
 wire \datamem.data_ram[49][16] ;
 wire \datamem.data_ram[49][17] ;
 wire \datamem.data_ram[49][18] ;
 wire \datamem.data_ram[49][19] ;
 wire \datamem.data_ram[49][1] ;
 wire \datamem.data_ram[49][20] ;
 wire \datamem.data_ram[49][21] ;
 wire \datamem.data_ram[49][22] ;
 wire \datamem.data_ram[49][23] ;
 wire \datamem.data_ram[49][24] ;
 wire \datamem.data_ram[49][25] ;
 wire \datamem.data_ram[49][26] ;
 wire \datamem.data_ram[49][27] ;
 wire \datamem.data_ram[49][28] ;
 wire \datamem.data_ram[49][29] ;
 wire \datamem.data_ram[49][2] ;
 wire \datamem.data_ram[49][30] ;
 wire \datamem.data_ram[49][31] ;
 wire \datamem.data_ram[49][3] ;
 wire \datamem.data_ram[49][4] ;
 wire \datamem.data_ram[49][5] ;
 wire \datamem.data_ram[49][6] ;
 wire \datamem.data_ram[49][7] ;
 wire \datamem.data_ram[49][8] ;
 wire \datamem.data_ram[49][9] ;
 wire \datamem.data_ram[4][0] ;
 wire \datamem.data_ram[4][10] ;
 wire \datamem.data_ram[4][11] ;
 wire \datamem.data_ram[4][12] ;
 wire \datamem.data_ram[4][13] ;
 wire \datamem.data_ram[4][14] ;
 wire \datamem.data_ram[4][15] ;
 wire \datamem.data_ram[4][16] ;
 wire \datamem.data_ram[4][17] ;
 wire \datamem.data_ram[4][18] ;
 wire \datamem.data_ram[4][19] ;
 wire \datamem.data_ram[4][1] ;
 wire \datamem.data_ram[4][20] ;
 wire \datamem.data_ram[4][21] ;
 wire \datamem.data_ram[4][22] ;
 wire \datamem.data_ram[4][23] ;
 wire \datamem.data_ram[4][24] ;
 wire \datamem.data_ram[4][25] ;
 wire \datamem.data_ram[4][26] ;
 wire \datamem.data_ram[4][27] ;
 wire \datamem.data_ram[4][28] ;
 wire \datamem.data_ram[4][29] ;
 wire \datamem.data_ram[4][2] ;
 wire \datamem.data_ram[4][30] ;
 wire \datamem.data_ram[4][31] ;
 wire \datamem.data_ram[4][3] ;
 wire \datamem.data_ram[4][4] ;
 wire \datamem.data_ram[4][5] ;
 wire \datamem.data_ram[4][6] ;
 wire \datamem.data_ram[4][7] ;
 wire \datamem.data_ram[4][8] ;
 wire \datamem.data_ram[4][9] ;
 wire \datamem.data_ram[50][0] ;
 wire \datamem.data_ram[50][10] ;
 wire \datamem.data_ram[50][11] ;
 wire \datamem.data_ram[50][12] ;
 wire \datamem.data_ram[50][13] ;
 wire \datamem.data_ram[50][14] ;
 wire \datamem.data_ram[50][15] ;
 wire \datamem.data_ram[50][16] ;
 wire \datamem.data_ram[50][17] ;
 wire \datamem.data_ram[50][18] ;
 wire \datamem.data_ram[50][19] ;
 wire \datamem.data_ram[50][1] ;
 wire \datamem.data_ram[50][20] ;
 wire \datamem.data_ram[50][21] ;
 wire \datamem.data_ram[50][22] ;
 wire \datamem.data_ram[50][23] ;
 wire \datamem.data_ram[50][24] ;
 wire \datamem.data_ram[50][25] ;
 wire \datamem.data_ram[50][26] ;
 wire \datamem.data_ram[50][27] ;
 wire \datamem.data_ram[50][28] ;
 wire \datamem.data_ram[50][29] ;
 wire \datamem.data_ram[50][2] ;
 wire \datamem.data_ram[50][30] ;
 wire \datamem.data_ram[50][31] ;
 wire \datamem.data_ram[50][3] ;
 wire \datamem.data_ram[50][4] ;
 wire \datamem.data_ram[50][5] ;
 wire \datamem.data_ram[50][6] ;
 wire \datamem.data_ram[50][7] ;
 wire \datamem.data_ram[50][8] ;
 wire \datamem.data_ram[50][9] ;
 wire \datamem.data_ram[51][0] ;
 wire \datamem.data_ram[51][10] ;
 wire \datamem.data_ram[51][11] ;
 wire \datamem.data_ram[51][12] ;
 wire \datamem.data_ram[51][13] ;
 wire \datamem.data_ram[51][14] ;
 wire \datamem.data_ram[51][15] ;
 wire \datamem.data_ram[51][16] ;
 wire \datamem.data_ram[51][17] ;
 wire \datamem.data_ram[51][18] ;
 wire \datamem.data_ram[51][19] ;
 wire \datamem.data_ram[51][1] ;
 wire \datamem.data_ram[51][20] ;
 wire \datamem.data_ram[51][21] ;
 wire \datamem.data_ram[51][22] ;
 wire \datamem.data_ram[51][23] ;
 wire \datamem.data_ram[51][24] ;
 wire \datamem.data_ram[51][25] ;
 wire \datamem.data_ram[51][26] ;
 wire \datamem.data_ram[51][27] ;
 wire \datamem.data_ram[51][28] ;
 wire \datamem.data_ram[51][29] ;
 wire \datamem.data_ram[51][2] ;
 wire \datamem.data_ram[51][30] ;
 wire \datamem.data_ram[51][31] ;
 wire \datamem.data_ram[51][3] ;
 wire \datamem.data_ram[51][4] ;
 wire \datamem.data_ram[51][5] ;
 wire \datamem.data_ram[51][6] ;
 wire \datamem.data_ram[51][7] ;
 wire \datamem.data_ram[51][8] ;
 wire \datamem.data_ram[51][9] ;
 wire \datamem.data_ram[52][0] ;
 wire \datamem.data_ram[52][10] ;
 wire \datamem.data_ram[52][11] ;
 wire \datamem.data_ram[52][12] ;
 wire \datamem.data_ram[52][13] ;
 wire \datamem.data_ram[52][14] ;
 wire \datamem.data_ram[52][15] ;
 wire \datamem.data_ram[52][16] ;
 wire \datamem.data_ram[52][17] ;
 wire \datamem.data_ram[52][18] ;
 wire \datamem.data_ram[52][19] ;
 wire \datamem.data_ram[52][1] ;
 wire \datamem.data_ram[52][20] ;
 wire \datamem.data_ram[52][21] ;
 wire \datamem.data_ram[52][22] ;
 wire \datamem.data_ram[52][23] ;
 wire \datamem.data_ram[52][24] ;
 wire \datamem.data_ram[52][25] ;
 wire \datamem.data_ram[52][26] ;
 wire \datamem.data_ram[52][27] ;
 wire \datamem.data_ram[52][28] ;
 wire \datamem.data_ram[52][29] ;
 wire \datamem.data_ram[52][2] ;
 wire \datamem.data_ram[52][30] ;
 wire \datamem.data_ram[52][31] ;
 wire \datamem.data_ram[52][3] ;
 wire \datamem.data_ram[52][4] ;
 wire \datamem.data_ram[52][5] ;
 wire \datamem.data_ram[52][6] ;
 wire \datamem.data_ram[52][7] ;
 wire \datamem.data_ram[52][8] ;
 wire \datamem.data_ram[52][9] ;
 wire \datamem.data_ram[53][0] ;
 wire \datamem.data_ram[53][10] ;
 wire \datamem.data_ram[53][11] ;
 wire \datamem.data_ram[53][12] ;
 wire \datamem.data_ram[53][13] ;
 wire \datamem.data_ram[53][14] ;
 wire \datamem.data_ram[53][15] ;
 wire \datamem.data_ram[53][16] ;
 wire \datamem.data_ram[53][17] ;
 wire \datamem.data_ram[53][18] ;
 wire \datamem.data_ram[53][19] ;
 wire \datamem.data_ram[53][1] ;
 wire \datamem.data_ram[53][20] ;
 wire \datamem.data_ram[53][21] ;
 wire \datamem.data_ram[53][22] ;
 wire \datamem.data_ram[53][23] ;
 wire \datamem.data_ram[53][24] ;
 wire \datamem.data_ram[53][25] ;
 wire \datamem.data_ram[53][26] ;
 wire \datamem.data_ram[53][27] ;
 wire \datamem.data_ram[53][28] ;
 wire \datamem.data_ram[53][29] ;
 wire \datamem.data_ram[53][2] ;
 wire \datamem.data_ram[53][30] ;
 wire \datamem.data_ram[53][31] ;
 wire \datamem.data_ram[53][3] ;
 wire \datamem.data_ram[53][4] ;
 wire \datamem.data_ram[53][5] ;
 wire \datamem.data_ram[53][6] ;
 wire \datamem.data_ram[53][7] ;
 wire \datamem.data_ram[53][8] ;
 wire \datamem.data_ram[53][9] ;
 wire \datamem.data_ram[54][0] ;
 wire \datamem.data_ram[54][10] ;
 wire \datamem.data_ram[54][11] ;
 wire \datamem.data_ram[54][12] ;
 wire \datamem.data_ram[54][13] ;
 wire \datamem.data_ram[54][14] ;
 wire \datamem.data_ram[54][15] ;
 wire \datamem.data_ram[54][16] ;
 wire \datamem.data_ram[54][17] ;
 wire \datamem.data_ram[54][18] ;
 wire \datamem.data_ram[54][19] ;
 wire \datamem.data_ram[54][1] ;
 wire \datamem.data_ram[54][20] ;
 wire \datamem.data_ram[54][21] ;
 wire \datamem.data_ram[54][22] ;
 wire \datamem.data_ram[54][23] ;
 wire \datamem.data_ram[54][24] ;
 wire \datamem.data_ram[54][25] ;
 wire \datamem.data_ram[54][26] ;
 wire \datamem.data_ram[54][27] ;
 wire \datamem.data_ram[54][28] ;
 wire \datamem.data_ram[54][29] ;
 wire \datamem.data_ram[54][2] ;
 wire \datamem.data_ram[54][30] ;
 wire \datamem.data_ram[54][31] ;
 wire \datamem.data_ram[54][3] ;
 wire \datamem.data_ram[54][4] ;
 wire \datamem.data_ram[54][5] ;
 wire \datamem.data_ram[54][6] ;
 wire \datamem.data_ram[54][7] ;
 wire \datamem.data_ram[54][8] ;
 wire \datamem.data_ram[54][9] ;
 wire \datamem.data_ram[55][0] ;
 wire \datamem.data_ram[55][10] ;
 wire \datamem.data_ram[55][11] ;
 wire \datamem.data_ram[55][12] ;
 wire \datamem.data_ram[55][13] ;
 wire \datamem.data_ram[55][14] ;
 wire \datamem.data_ram[55][15] ;
 wire \datamem.data_ram[55][16] ;
 wire \datamem.data_ram[55][17] ;
 wire \datamem.data_ram[55][18] ;
 wire \datamem.data_ram[55][19] ;
 wire \datamem.data_ram[55][1] ;
 wire \datamem.data_ram[55][20] ;
 wire \datamem.data_ram[55][21] ;
 wire \datamem.data_ram[55][22] ;
 wire \datamem.data_ram[55][23] ;
 wire \datamem.data_ram[55][24] ;
 wire \datamem.data_ram[55][25] ;
 wire \datamem.data_ram[55][26] ;
 wire \datamem.data_ram[55][27] ;
 wire \datamem.data_ram[55][28] ;
 wire \datamem.data_ram[55][29] ;
 wire \datamem.data_ram[55][2] ;
 wire \datamem.data_ram[55][30] ;
 wire \datamem.data_ram[55][31] ;
 wire \datamem.data_ram[55][3] ;
 wire \datamem.data_ram[55][4] ;
 wire \datamem.data_ram[55][5] ;
 wire \datamem.data_ram[55][6] ;
 wire \datamem.data_ram[55][7] ;
 wire \datamem.data_ram[55][8] ;
 wire \datamem.data_ram[55][9] ;
 wire \datamem.data_ram[56][0] ;
 wire \datamem.data_ram[56][10] ;
 wire \datamem.data_ram[56][11] ;
 wire \datamem.data_ram[56][12] ;
 wire \datamem.data_ram[56][13] ;
 wire \datamem.data_ram[56][14] ;
 wire \datamem.data_ram[56][15] ;
 wire \datamem.data_ram[56][16] ;
 wire \datamem.data_ram[56][17] ;
 wire \datamem.data_ram[56][18] ;
 wire \datamem.data_ram[56][19] ;
 wire \datamem.data_ram[56][1] ;
 wire \datamem.data_ram[56][20] ;
 wire \datamem.data_ram[56][21] ;
 wire \datamem.data_ram[56][22] ;
 wire \datamem.data_ram[56][23] ;
 wire \datamem.data_ram[56][24] ;
 wire \datamem.data_ram[56][25] ;
 wire \datamem.data_ram[56][26] ;
 wire \datamem.data_ram[56][27] ;
 wire \datamem.data_ram[56][28] ;
 wire \datamem.data_ram[56][29] ;
 wire \datamem.data_ram[56][2] ;
 wire \datamem.data_ram[56][30] ;
 wire \datamem.data_ram[56][31] ;
 wire \datamem.data_ram[56][3] ;
 wire \datamem.data_ram[56][4] ;
 wire \datamem.data_ram[56][5] ;
 wire \datamem.data_ram[56][6] ;
 wire \datamem.data_ram[56][7] ;
 wire \datamem.data_ram[56][8] ;
 wire \datamem.data_ram[56][9] ;
 wire \datamem.data_ram[57][0] ;
 wire \datamem.data_ram[57][10] ;
 wire \datamem.data_ram[57][11] ;
 wire \datamem.data_ram[57][12] ;
 wire \datamem.data_ram[57][13] ;
 wire \datamem.data_ram[57][14] ;
 wire \datamem.data_ram[57][15] ;
 wire \datamem.data_ram[57][16] ;
 wire \datamem.data_ram[57][17] ;
 wire \datamem.data_ram[57][18] ;
 wire \datamem.data_ram[57][19] ;
 wire \datamem.data_ram[57][1] ;
 wire \datamem.data_ram[57][20] ;
 wire \datamem.data_ram[57][21] ;
 wire \datamem.data_ram[57][22] ;
 wire \datamem.data_ram[57][23] ;
 wire \datamem.data_ram[57][24] ;
 wire \datamem.data_ram[57][25] ;
 wire \datamem.data_ram[57][26] ;
 wire \datamem.data_ram[57][27] ;
 wire \datamem.data_ram[57][28] ;
 wire \datamem.data_ram[57][29] ;
 wire \datamem.data_ram[57][2] ;
 wire \datamem.data_ram[57][30] ;
 wire \datamem.data_ram[57][31] ;
 wire \datamem.data_ram[57][3] ;
 wire \datamem.data_ram[57][4] ;
 wire \datamem.data_ram[57][5] ;
 wire \datamem.data_ram[57][6] ;
 wire \datamem.data_ram[57][7] ;
 wire \datamem.data_ram[57][8] ;
 wire \datamem.data_ram[57][9] ;
 wire \datamem.data_ram[58][0] ;
 wire \datamem.data_ram[58][10] ;
 wire \datamem.data_ram[58][11] ;
 wire \datamem.data_ram[58][12] ;
 wire \datamem.data_ram[58][13] ;
 wire \datamem.data_ram[58][14] ;
 wire \datamem.data_ram[58][15] ;
 wire \datamem.data_ram[58][16] ;
 wire \datamem.data_ram[58][17] ;
 wire \datamem.data_ram[58][18] ;
 wire \datamem.data_ram[58][19] ;
 wire \datamem.data_ram[58][1] ;
 wire \datamem.data_ram[58][20] ;
 wire \datamem.data_ram[58][21] ;
 wire \datamem.data_ram[58][22] ;
 wire \datamem.data_ram[58][23] ;
 wire \datamem.data_ram[58][24] ;
 wire \datamem.data_ram[58][25] ;
 wire \datamem.data_ram[58][26] ;
 wire \datamem.data_ram[58][27] ;
 wire \datamem.data_ram[58][28] ;
 wire \datamem.data_ram[58][29] ;
 wire \datamem.data_ram[58][2] ;
 wire \datamem.data_ram[58][30] ;
 wire \datamem.data_ram[58][31] ;
 wire \datamem.data_ram[58][3] ;
 wire \datamem.data_ram[58][4] ;
 wire \datamem.data_ram[58][5] ;
 wire \datamem.data_ram[58][6] ;
 wire \datamem.data_ram[58][7] ;
 wire \datamem.data_ram[58][8] ;
 wire \datamem.data_ram[58][9] ;
 wire \datamem.data_ram[59][0] ;
 wire \datamem.data_ram[59][10] ;
 wire \datamem.data_ram[59][11] ;
 wire \datamem.data_ram[59][12] ;
 wire \datamem.data_ram[59][13] ;
 wire \datamem.data_ram[59][14] ;
 wire \datamem.data_ram[59][15] ;
 wire \datamem.data_ram[59][16] ;
 wire \datamem.data_ram[59][17] ;
 wire \datamem.data_ram[59][18] ;
 wire \datamem.data_ram[59][19] ;
 wire \datamem.data_ram[59][1] ;
 wire \datamem.data_ram[59][20] ;
 wire \datamem.data_ram[59][21] ;
 wire \datamem.data_ram[59][22] ;
 wire \datamem.data_ram[59][23] ;
 wire \datamem.data_ram[59][24] ;
 wire \datamem.data_ram[59][25] ;
 wire \datamem.data_ram[59][26] ;
 wire \datamem.data_ram[59][27] ;
 wire \datamem.data_ram[59][28] ;
 wire \datamem.data_ram[59][29] ;
 wire \datamem.data_ram[59][2] ;
 wire \datamem.data_ram[59][30] ;
 wire \datamem.data_ram[59][31] ;
 wire \datamem.data_ram[59][3] ;
 wire \datamem.data_ram[59][4] ;
 wire \datamem.data_ram[59][5] ;
 wire \datamem.data_ram[59][6] ;
 wire \datamem.data_ram[59][7] ;
 wire \datamem.data_ram[59][8] ;
 wire \datamem.data_ram[59][9] ;
 wire \datamem.data_ram[5][0] ;
 wire \datamem.data_ram[5][10] ;
 wire \datamem.data_ram[5][11] ;
 wire \datamem.data_ram[5][12] ;
 wire \datamem.data_ram[5][13] ;
 wire \datamem.data_ram[5][14] ;
 wire \datamem.data_ram[5][15] ;
 wire \datamem.data_ram[5][16] ;
 wire \datamem.data_ram[5][17] ;
 wire \datamem.data_ram[5][18] ;
 wire \datamem.data_ram[5][19] ;
 wire \datamem.data_ram[5][1] ;
 wire \datamem.data_ram[5][20] ;
 wire \datamem.data_ram[5][21] ;
 wire \datamem.data_ram[5][22] ;
 wire \datamem.data_ram[5][23] ;
 wire \datamem.data_ram[5][24] ;
 wire \datamem.data_ram[5][25] ;
 wire \datamem.data_ram[5][26] ;
 wire \datamem.data_ram[5][27] ;
 wire \datamem.data_ram[5][28] ;
 wire \datamem.data_ram[5][29] ;
 wire \datamem.data_ram[5][2] ;
 wire \datamem.data_ram[5][30] ;
 wire \datamem.data_ram[5][31] ;
 wire \datamem.data_ram[5][3] ;
 wire \datamem.data_ram[5][4] ;
 wire \datamem.data_ram[5][5] ;
 wire \datamem.data_ram[5][6] ;
 wire \datamem.data_ram[5][7] ;
 wire \datamem.data_ram[5][8] ;
 wire \datamem.data_ram[5][9] ;
 wire \datamem.data_ram[60][0] ;
 wire \datamem.data_ram[60][10] ;
 wire \datamem.data_ram[60][11] ;
 wire \datamem.data_ram[60][12] ;
 wire \datamem.data_ram[60][13] ;
 wire \datamem.data_ram[60][14] ;
 wire \datamem.data_ram[60][15] ;
 wire \datamem.data_ram[60][16] ;
 wire \datamem.data_ram[60][17] ;
 wire \datamem.data_ram[60][18] ;
 wire \datamem.data_ram[60][19] ;
 wire \datamem.data_ram[60][1] ;
 wire \datamem.data_ram[60][20] ;
 wire \datamem.data_ram[60][21] ;
 wire \datamem.data_ram[60][22] ;
 wire \datamem.data_ram[60][23] ;
 wire \datamem.data_ram[60][24] ;
 wire \datamem.data_ram[60][25] ;
 wire \datamem.data_ram[60][26] ;
 wire \datamem.data_ram[60][27] ;
 wire \datamem.data_ram[60][28] ;
 wire \datamem.data_ram[60][29] ;
 wire \datamem.data_ram[60][2] ;
 wire \datamem.data_ram[60][30] ;
 wire \datamem.data_ram[60][31] ;
 wire \datamem.data_ram[60][3] ;
 wire \datamem.data_ram[60][4] ;
 wire \datamem.data_ram[60][5] ;
 wire \datamem.data_ram[60][6] ;
 wire \datamem.data_ram[60][7] ;
 wire \datamem.data_ram[60][8] ;
 wire \datamem.data_ram[60][9] ;
 wire \datamem.data_ram[61][0] ;
 wire \datamem.data_ram[61][10] ;
 wire \datamem.data_ram[61][11] ;
 wire \datamem.data_ram[61][12] ;
 wire \datamem.data_ram[61][13] ;
 wire \datamem.data_ram[61][14] ;
 wire \datamem.data_ram[61][15] ;
 wire \datamem.data_ram[61][16] ;
 wire \datamem.data_ram[61][17] ;
 wire \datamem.data_ram[61][18] ;
 wire \datamem.data_ram[61][19] ;
 wire \datamem.data_ram[61][1] ;
 wire \datamem.data_ram[61][20] ;
 wire \datamem.data_ram[61][21] ;
 wire \datamem.data_ram[61][22] ;
 wire \datamem.data_ram[61][23] ;
 wire \datamem.data_ram[61][24] ;
 wire \datamem.data_ram[61][25] ;
 wire \datamem.data_ram[61][26] ;
 wire \datamem.data_ram[61][27] ;
 wire \datamem.data_ram[61][28] ;
 wire \datamem.data_ram[61][29] ;
 wire \datamem.data_ram[61][2] ;
 wire \datamem.data_ram[61][30] ;
 wire \datamem.data_ram[61][31] ;
 wire \datamem.data_ram[61][3] ;
 wire \datamem.data_ram[61][4] ;
 wire \datamem.data_ram[61][5] ;
 wire \datamem.data_ram[61][6] ;
 wire \datamem.data_ram[61][7] ;
 wire \datamem.data_ram[61][8] ;
 wire \datamem.data_ram[61][9] ;
 wire \datamem.data_ram[62][0] ;
 wire \datamem.data_ram[62][10] ;
 wire \datamem.data_ram[62][11] ;
 wire \datamem.data_ram[62][12] ;
 wire \datamem.data_ram[62][13] ;
 wire \datamem.data_ram[62][14] ;
 wire \datamem.data_ram[62][15] ;
 wire \datamem.data_ram[62][16] ;
 wire \datamem.data_ram[62][17] ;
 wire \datamem.data_ram[62][18] ;
 wire \datamem.data_ram[62][19] ;
 wire \datamem.data_ram[62][1] ;
 wire \datamem.data_ram[62][20] ;
 wire \datamem.data_ram[62][21] ;
 wire \datamem.data_ram[62][22] ;
 wire \datamem.data_ram[62][23] ;
 wire \datamem.data_ram[62][24] ;
 wire \datamem.data_ram[62][25] ;
 wire \datamem.data_ram[62][26] ;
 wire \datamem.data_ram[62][27] ;
 wire \datamem.data_ram[62][28] ;
 wire \datamem.data_ram[62][29] ;
 wire \datamem.data_ram[62][2] ;
 wire \datamem.data_ram[62][30] ;
 wire \datamem.data_ram[62][31] ;
 wire \datamem.data_ram[62][3] ;
 wire \datamem.data_ram[62][4] ;
 wire \datamem.data_ram[62][5] ;
 wire \datamem.data_ram[62][6] ;
 wire \datamem.data_ram[62][7] ;
 wire \datamem.data_ram[62][8] ;
 wire \datamem.data_ram[62][9] ;
 wire \datamem.data_ram[63][0] ;
 wire \datamem.data_ram[63][10] ;
 wire \datamem.data_ram[63][11] ;
 wire \datamem.data_ram[63][12] ;
 wire \datamem.data_ram[63][13] ;
 wire \datamem.data_ram[63][14] ;
 wire \datamem.data_ram[63][15] ;
 wire \datamem.data_ram[63][16] ;
 wire \datamem.data_ram[63][17] ;
 wire \datamem.data_ram[63][18] ;
 wire \datamem.data_ram[63][19] ;
 wire \datamem.data_ram[63][1] ;
 wire \datamem.data_ram[63][20] ;
 wire \datamem.data_ram[63][21] ;
 wire \datamem.data_ram[63][22] ;
 wire \datamem.data_ram[63][23] ;
 wire \datamem.data_ram[63][24] ;
 wire \datamem.data_ram[63][25] ;
 wire \datamem.data_ram[63][26] ;
 wire \datamem.data_ram[63][27] ;
 wire \datamem.data_ram[63][28] ;
 wire \datamem.data_ram[63][29] ;
 wire \datamem.data_ram[63][2] ;
 wire \datamem.data_ram[63][30] ;
 wire \datamem.data_ram[63][31] ;
 wire \datamem.data_ram[63][3] ;
 wire \datamem.data_ram[63][4] ;
 wire \datamem.data_ram[63][5] ;
 wire \datamem.data_ram[63][6] ;
 wire \datamem.data_ram[63][7] ;
 wire \datamem.data_ram[63][8] ;
 wire \datamem.data_ram[63][9] ;
 wire \datamem.data_ram[6][0] ;
 wire \datamem.data_ram[6][10] ;
 wire \datamem.data_ram[6][11] ;
 wire \datamem.data_ram[6][12] ;
 wire \datamem.data_ram[6][13] ;
 wire \datamem.data_ram[6][14] ;
 wire \datamem.data_ram[6][15] ;
 wire \datamem.data_ram[6][16] ;
 wire \datamem.data_ram[6][17] ;
 wire \datamem.data_ram[6][18] ;
 wire \datamem.data_ram[6][19] ;
 wire \datamem.data_ram[6][1] ;
 wire \datamem.data_ram[6][20] ;
 wire \datamem.data_ram[6][21] ;
 wire \datamem.data_ram[6][22] ;
 wire \datamem.data_ram[6][23] ;
 wire \datamem.data_ram[6][24] ;
 wire \datamem.data_ram[6][25] ;
 wire \datamem.data_ram[6][26] ;
 wire \datamem.data_ram[6][27] ;
 wire \datamem.data_ram[6][28] ;
 wire \datamem.data_ram[6][29] ;
 wire \datamem.data_ram[6][2] ;
 wire \datamem.data_ram[6][30] ;
 wire \datamem.data_ram[6][31] ;
 wire \datamem.data_ram[6][3] ;
 wire \datamem.data_ram[6][4] ;
 wire \datamem.data_ram[6][5] ;
 wire \datamem.data_ram[6][6] ;
 wire \datamem.data_ram[6][7] ;
 wire \datamem.data_ram[6][8] ;
 wire \datamem.data_ram[6][9] ;
 wire \datamem.data_ram[7][0] ;
 wire \datamem.data_ram[7][10] ;
 wire \datamem.data_ram[7][11] ;
 wire \datamem.data_ram[7][12] ;
 wire \datamem.data_ram[7][13] ;
 wire \datamem.data_ram[7][14] ;
 wire \datamem.data_ram[7][15] ;
 wire \datamem.data_ram[7][16] ;
 wire \datamem.data_ram[7][17] ;
 wire \datamem.data_ram[7][18] ;
 wire \datamem.data_ram[7][19] ;
 wire \datamem.data_ram[7][1] ;
 wire \datamem.data_ram[7][20] ;
 wire \datamem.data_ram[7][21] ;
 wire \datamem.data_ram[7][22] ;
 wire \datamem.data_ram[7][23] ;
 wire \datamem.data_ram[7][24] ;
 wire \datamem.data_ram[7][25] ;
 wire \datamem.data_ram[7][26] ;
 wire \datamem.data_ram[7][27] ;
 wire \datamem.data_ram[7][28] ;
 wire \datamem.data_ram[7][29] ;
 wire \datamem.data_ram[7][2] ;
 wire \datamem.data_ram[7][30] ;
 wire \datamem.data_ram[7][31] ;
 wire \datamem.data_ram[7][3] ;
 wire \datamem.data_ram[7][4] ;
 wire \datamem.data_ram[7][5] ;
 wire \datamem.data_ram[7][6] ;
 wire \datamem.data_ram[7][7] ;
 wire \datamem.data_ram[7][8] ;
 wire \datamem.data_ram[7][9] ;
 wire \datamem.data_ram[8][0] ;
 wire \datamem.data_ram[8][10] ;
 wire \datamem.data_ram[8][11] ;
 wire \datamem.data_ram[8][12] ;
 wire \datamem.data_ram[8][13] ;
 wire \datamem.data_ram[8][14] ;
 wire \datamem.data_ram[8][15] ;
 wire \datamem.data_ram[8][16] ;
 wire \datamem.data_ram[8][17] ;
 wire \datamem.data_ram[8][18] ;
 wire \datamem.data_ram[8][19] ;
 wire \datamem.data_ram[8][1] ;
 wire \datamem.data_ram[8][20] ;
 wire \datamem.data_ram[8][21] ;
 wire \datamem.data_ram[8][22] ;
 wire \datamem.data_ram[8][23] ;
 wire \datamem.data_ram[8][24] ;
 wire \datamem.data_ram[8][25] ;
 wire \datamem.data_ram[8][26] ;
 wire \datamem.data_ram[8][27] ;
 wire \datamem.data_ram[8][28] ;
 wire \datamem.data_ram[8][29] ;
 wire \datamem.data_ram[8][2] ;
 wire \datamem.data_ram[8][30] ;
 wire \datamem.data_ram[8][31] ;
 wire \datamem.data_ram[8][3] ;
 wire \datamem.data_ram[8][4] ;
 wire \datamem.data_ram[8][5] ;
 wire \datamem.data_ram[8][6] ;
 wire \datamem.data_ram[8][7] ;
 wire \datamem.data_ram[8][8] ;
 wire \datamem.data_ram[8][9] ;
 wire \datamem.data_ram[9][0] ;
 wire \datamem.data_ram[9][10] ;
 wire \datamem.data_ram[9][11] ;
 wire \datamem.data_ram[9][12] ;
 wire \datamem.data_ram[9][13] ;
 wire \datamem.data_ram[9][14] ;
 wire \datamem.data_ram[9][15] ;
 wire \datamem.data_ram[9][16] ;
 wire \datamem.data_ram[9][17] ;
 wire \datamem.data_ram[9][18] ;
 wire \datamem.data_ram[9][19] ;
 wire \datamem.data_ram[9][1] ;
 wire \datamem.data_ram[9][20] ;
 wire \datamem.data_ram[9][21] ;
 wire \datamem.data_ram[9][22] ;
 wire \datamem.data_ram[9][23] ;
 wire \datamem.data_ram[9][24] ;
 wire \datamem.data_ram[9][25] ;
 wire \datamem.data_ram[9][26] ;
 wire \datamem.data_ram[9][27] ;
 wire \datamem.data_ram[9][28] ;
 wire \datamem.data_ram[9][29] ;
 wire \datamem.data_ram[9][2] ;
 wire \datamem.data_ram[9][30] ;
 wire \datamem.data_ram[9][31] ;
 wire \datamem.data_ram[9][3] ;
 wire \datamem.data_ram[9][4] ;
 wire \datamem.data_ram[9][5] ;
 wire \datamem.data_ram[9][6] ;
 wire \datamem.data_ram[9][7] ;
 wire \datamem.data_ram[9][8] ;
 wire \datamem.data_ram[9][9] ;
 wire \datamem.rd_data_mem[0] ;
 wire \datamem.rd_data_mem[10] ;
 wire \datamem.rd_data_mem[11] ;
 wire \datamem.rd_data_mem[12] ;
 wire \datamem.rd_data_mem[13] ;
 wire \datamem.rd_data_mem[14] ;
 wire \datamem.rd_data_mem[15] ;
 wire \datamem.rd_data_mem[16] ;
 wire \datamem.rd_data_mem[17] ;
 wire \datamem.rd_data_mem[18] ;
 wire \datamem.rd_data_mem[19] ;
 wire \datamem.rd_data_mem[1] ;
 wire \datamem.rd_data_mem[20] ;
 wire \datamem.rd_data_mem[21] ;
 wire \datamem.rd_data_mem[22] ;
 wire \datamem.rd_data_mem[23] ;
 wire \datamem.rd_data_mem[24] ;
 wire \datamem.rd_data_mem[25] ;
 wire \datamem.rd_data_mem[26] ;
 wire \datamem.rd_data_mem[27] ;
 wire \datamem.rd_data_mem[28] ;
 wire \datamem.rd_data_mem[29] ;
 wire \datamem.rd_data_mem[2] ;
 wire \datamem.rd_data_mem[30] ;
 wire \datamem.rd_data_mem[31] ;
 wire \datamem.rd_data_mem[3] ;
 wire \datamem.rd_data_mem[4] ;
 wire \datamem.rd_data_mem[5] ;
 wire \datamem.rd_data_mem[6] ;
 wire \datamem.rd_data_mem[7] ;
 wire \datamem.rd_data_mem[8] ;
 wire \datamem.rd_data_mem[9] ;
 wire \rvcpu.ALUControl[0] ;
 wire \rvcpu.ALUControl[1] ;
 wire \rvcpu.ALUControl[2] ;
 wire \rvcpu.ALUControl[3] ;
 wire \rvcpu.ALUResultE[0] ;
 wire \rvcpu.ALUResultE[10] ;
 wire \rvcpu.ALUResultE[11] ;
 wire \rvcpu.ALUResultE[12] ;
 wire \rvcpu.ALUResultE[13] ;
 wire \rvcpu.ALUResultE[14] ;
 wire \rvcpu.ALUResultE[15] ;
 wire \rvcpu.ALUResultE[16] ;
 wire \rvcpu.ALUResultE[17] ;
 wire \rvcpu.ALUResultE[18] ;
 wire \rvcpu.ALUResultE[19] ;
 wire \rvcpu.ALUResultE[1] ;
 wire \rvcpu.ALUResultE[20] ;
 wire \rvcpu.ALUResultE[21] ;
 wire \rvcpu.ALUResultE[22] ;
 wire \rvcpu.ALUResultE[23] ;
 wire \rvcpu.ALUResultE[24] ;
 wire \rvcpu.ALUResultE[25] ;
 wire \rvcpu.ALUResultE[26] ;
 wire \rvcpu.ALUResultE[27] ;
 wire \rvcpu.ALUResultE[28] ;
 wire \rvcpu.ALUResultE[29] ;
 wire \rvcpu.ALUResultE[2] ;
 wire \rvcpu.ALUResultE[30] ;
 wire \rvcpu.ALUResultE[31] ;
 wire \rvcpu.ALUResultE[3] ;
 wire \rvcpu.ALUResultE[4] ;
 wire \rvcpu.ALUResultE[5] ;
 wire \rvcpu.ALUResultE[6] ;
 wire \rvcpu.ALUResultE[7] ;
 wire \rvcpu.ALUResultE[8] ;
 wire \rvcpu.ALUResultE[9] ;
 wire \rvcpu.c.ad.funct7b5 ;
 wire \rvcpu.c.ad.opb5 ;
 wire \rvcpu.dp.Cout ;
 wire \rvcpu.dp.SrcBFW_Mux.y[0] ;
 wire \rvcpu.dp.SrcBFW_Mux.y[10] ;
 wire \rvcpu.dp.SrcBFW_Mux.y[11] ;
 wire \rvcpu.dp.SrcBFW_Mux.y[12] ;
 wire \rvcpu.dp.SrcBFW_Mux.y[13] ;
 wire \rvcpu.dp.SrcBFW_Mux.y[14] ;
 wire \rvcpu.dp.SrcBFW_Mux.y[15] ;
 wire \rvcpu.dp.SrcBFW_Mux.y[16] ;
 wire \rvcpu.dp.SrcBFW_Mux.y[17] ;
 wire \rvcpu.dp.SrcBFW_Mux.y[18] ;
 wire \rvcpu.dp.SrcBFW_Mux.y[19] ;
 wire \rvcpu.dp.SrcBFW_Mux.y[1] ;
 wire \rvcpu.dp.SrcBFW_Mux.y[20] ;
 wire \rvcpu.dp.SrcBFW_Mux.y[21] ;
 wire \rvcpu.dp.SrcBFW_Mux.y[22] ;
 wire \rvcpu.dp.SrcBFW_Mux.y[23] ;
 wire \rvcpu.dp.SrcBFW_Mux.y[24] ;
 wire \rvcpu.dp.SrcBFW_Mux.y[25] ;
 wire \rvcpu.dp.SrcBFW_Mux.y[26] ;
 wire \rvcpu.dp.SrcBFW_Mux.y[27] ;
 wire \rvcpu.dp.SrcBFW_Mux.y[28] ;
 wire \rvcpu.dp.SrcBFW_Mux.y[29] ;
 wire \rvcpu.dp.SrcBFW_Mux.y[2] ;
 wire \rvcpu.dp.SrcBFW_Mux.y[30] ;
 wire \rvcpu.dp.SrcBFW_Mux.y[31] ;
 wire \rvcpu.dp.SrcBFW_Mux.y[3] ;
 wire \rvcpu.dp.SrcBFW_Mux.y[4] ;
 wire \rvcpu.dp.SrcBFW_Mux.y[5] ;
 wire \rvcpu.dp.SrcBFW_Mux.y[6] ;
 wire \rvcpu.dp.SrcBFW_Mux.y[7] ;
 wire \rvcpu.dp.SrcBFW_Mux.y[8] ;
 wire \rvcpu.dp.SrcBFW_Mux.y[9] ;
 wire \rvcpu.dp.hu.ResultSrcE0 ;
 wire \rvcpu.dp.lAuiPCE[0] ;
 wire \rvcpu.dp.lAuiPCE[10] ;
 wire \rvcpu.dp.lAuiPCE[11] ;
 wire \rvcpu.dp.lAuiPCE[12] ;
 wire \rvcpu.dp.lAuiPCE[13] ;
 wire \rvcpu.dp.lAuiPCE[14] ;
 wire \rvcpu.dp.lAuiPCE[15] ;
 wire \rvcpu.dp.lAuiPCE[16] ;
 wire \rvcpu.dp.lAuiPCE[17] ;
 wire \rvcpu.dp.lAuiPCE[18] ;
 wire \rvcpu.dp.lAuiPCE[19] ;
 wire \rvcpu.dp.lAuiPCE[1] ;
 wire \rvcpu.dp.lAuiPCE[20] ;
 wire \rvcpu.dp.lAuiPCE[21] ;
 wire \rvcpu.dp.lAuiPCE[22] ;
 wire \rvcpu.dp.lAuiPCE[23] ;
 wire \rvcpu.dp.lAuiPCE[24] ;
 wire \rvcpu.dp.lAuiPCE[25] ;
 wire \rvcpu.dp.lAuiPCE[26] ;
 wire \rvcpu.dp.lAuiPCE[27] ;
 wire \rvcpu.dp.lAuiPCE[28] ;
 wire \rvcpu.dp.lAuiPCE[29] ;
 wire \rvcpu.dp.lAuiPCE[2] ;
 wire \rvcpu.dp.lAuiPCE[30] ;
 wire \rvcpu.dp.lAuiPCE[31] ;
 wire \rvcpu.dp.lAuiPCE[3] ;
 wire \rvcpu.dp.lAuiPCE[4] ;
 wire \rvcpu.dp.lAuiPCE[5] ;
 wire \rvcpu.dp.lAuiPCE[6] ;
 wire \rvcpu.dp.lAuiPCE[7] ;
 wire \rvcpu.dp.lAuiPCE[8] ;
 wire \rvcpu.dp.lAuiPCE[9] ;
 wire \rvcpu.dp.pcreg.q[0] ;
 wire \rvcpu.dp.pcreg.q[10] ;
 wire \rvcpu.dp.pcreg.q[11] ;
 wire \rvcpu.dp.pcreg.q[12] ;
 wire \rvcpu.dp.pcreg.q[13] ;
 wire \rvcpu.dp.pcreg.q[14] ;
 wire \rvcpu.dp.pcreg.q[15] ;
 wire \rvcpu.dp.pcreg.q[16] ;
 wire \rvcpu.dp.pcreg.q[17] ;
 wire \rvcpu.dp.pcreg.q[18] ;
 wire \rvcpu.dp.pcreg.q[19] ;
 wire \rvcpu.dp.pcreg.q[1] ;
 wire \rvcpu.dp.pcreg.q[20] ;
 wire \rvcpu.dp.pcreg.q[21] ;
 wire \rvcpu.dp.pcreg.q[22] ;
 wire \rvcpu.dp.pcreg.q[23] ;
 wire \rvcpu.dp.pcreg.q[24] ;
 wire \rvcpu.dp.pcreg.q[25] ;
 wire \rvcpu.dp.pcreg.q[26] ;
 wire \rvcpu.dp.pcreg.q[27] ;
 wire \rvcpu.dp.pcreg.q[28] ;
 wire \rvcpu.dp.pcreg.q[29] ;
 wire \rvcpu.dp.pcreg.q[2] ;
 wire \rvcpu.dp.pcreg.q[30] ;
 wire \rvcpu.dp.pcreg.q[31] ;
 wire \rvcpu.dp.pcreg.q[3] ;
 wire \rvcpu.dp.pcreg.q[4] ;
 wire \rvcpu.dp.pcreg.q[5] ;
 wire \rvcpu.dp.pcreg.q[6] ;
 wire \rvcpu.dp.pcreg.q[7] ;
 wire \rvcpu.dp.pcreg.q[8] ;
 wire \rvcpu.dp.pcreg.q[9] ;
 wire \rvcpu.dp.plde.ALUControlE[0] ;
 wire \rvcpu.dp.plde.ALUControlE[1] ;
 wire \rvcpu.dp.plde.ALUControlE[2] ;
 wire \rvcpu.dp.plde.ALUControlE[3] ;
 wire \rvcpu.dp.plde.ALUSrcE ;
 wire \rvcpu.dp.plde.BranchE ;
 wire \rvcpu.dp.plde.ImmExtE[0] ;
 wire \rvcpu.dp.plde.ImmExtE[10] ;
 wire \rvcpu.dp.plde.ImmExtE[11] ;
 wire \rvcpu.dp.plde.ImmExtE[12] ;
 wire \rvcpu.dp.plde.ImmExtE[13] ;
 wire \rvcpu.dp.plde.ImmExtE[14] ;
 wire \rvcpu.dp.plde.ImmExtE[15] ;
 wire \rvcpu.dp.plde.ImmExtE[16] ;
 wire \rvcpu.dp.plde.ImmExtE[17] ;
 wire \rvcpu.dp.plde.ImmExtE[18] ;
 wire \rvcpu.dp.plde.ImmExtE[19] ;
 wire \rvcpu.dp.plde.ImmExtE[1] ;
 wire \rvcpu.dp.plde.ImmExtE[20] ;
 wire \rvcpu.dp.plde.ImmExtE[21] ;
 wire \rvcpu.dp.plde.ImmExtE[22] ;
 wire \rvcpu.dp.plde.ImmExtE[23] ;
 wire \rvcpu.dp.plde.ImmExtE[24] ;
 wire \rvcpu.dp.plde.ImmExtE[25] ;
 wire \rvcpu.dp.plde.ImmExtE[26] ;
 wire \rvcpu.dp.plde.ImmExtE[27] ;
 wire \rvcpu.dp.plde.ImmExtE[28] ;
 wire \rvcpu.dp.plde.ImmExtE[29] ;
 wire \rvcpu.dp.plde.ImmExtE[2] ;
 wire \rvcpu.dp.plde.ImmExtE[30] ;
 wire \rvcpu.dp.plde.ImmExtE[31] ;
 wire \rvcpu.dp.plde.ImmExtE[3] ;
 wire \rvcpu.dp.plde.ImmExtE[4] ;
 wire \rvcpu.dp.plde.ImmExtE[5] ;
 wire \rvcpu.dp.plde.ImmExtE[6] ;
 wire \rvcpu.dp.plde.ImmExtE[7] ;
 wire \rvcpu.dp.plde.ImmExtE[8] ;
 wire \rvcpu.dp.plde.ImmExtE[9] ;
 wire \rvcpu.dp.plde.JalrE ;
 wire \rvcpu.dp.plde.JumpE ;
 wire \rvcpu.dp.plde.MemWriteE ;
 wire \rvcpu.dp.plde.PCE[0] ;
 wire \rvcpu.dp.plde.PCE[10] ;
 wire \rvcpu.dp.plde.PCE[11] ;
 wire \rvcpu.dp.plde.PCE[12] ;
 wire \rvcpu.dp.plde.PCE[13] ;
 wire \rvcpu.dp.plde.PCE[14] ;
 wire \rvcpu.dp.plde.PCE[15] ;
 wire \rvcpu.dp.plde.PCE[16] ;
 wire \rvcpu.dp.plde.PCE[17] ;
 wire \rvcpu.dp.plde.PCE[18] ;
 wire \rvcpu.dp.plde.PCE[19] ;
 wire \rvcpu.dp.plde.PCE[1] ;
 wire \rvcpu.dp.plde.PCE[20] ;
 wire \rvcpu.dp.plde.PCE[21] ;
 wire \rvcpu.dp.plde.PCE[22] ;
 wire \rvcpu.dp.plde.PCE[23] ;
 wire \rvcpu.dp.plde.PCE[24] ;
 wire \rvcpu.dp.plde.PCE[25] ;
 wire \rvcpu.dp.plde.PCE[26] ;
 wire \rvcpu.dp.plde.PCE[27] ;
 wire \rvcpu.dp.plde.PCE[28] ;
 wire \rvcpu.dp.plde.PCE[29] ;
 wire \rvcpu.dp.plde.PCE[2] ;
 wire \rvcpu.dp.plde.PCE[30] ;
 wire \rvcpu.dp.plde.PCE[31] ;
 wire \rvcpu.dp.plde.PCE[3] ;
 wire \rvcpu.dp.plde.PCE[4] ;
 wire \rvcpu.dp.plde.PCE[5] ;
 wire \rvcpu.dp.plde.PCE[6] ;
 wire \rvcpu.dp.plde.PCE[7] ;
 wire \rvcpu.dp.plde.PCE[8] ;
 wire \rvcpu.dp.plde.PCE[9] ;
 wire \rvcpu.dp.plde.PCPlus4E[10] ;
 wire \rvcpu.dp.plde.PCPlus4E[11] ;
 wire \rvcpu.dp.plde.PCPlus4E[12] ;
 wire \rvcpu.dp.plde.PCPlus4E[13] ;
 wire \rvcpu.dp.plde.PCPlus4E[14] ;
 wire \rvcpu.dp.plde.PCPlus4E[15] ;
 wire \rvcpu.dp.plde.PCPlus4E[16] ;
 wire \rvcpu.dp.plde.PCPlus4E[17] ;
 wire \rvcpu.dp.plde.PCPlus4E[18] ;
 wire \rvcpu.dp.plde.PCPlus4E[19] ;
 wire \rvcpu.dp.plde.PCPlus4E[20] ;
 wire \rvcpu.dp.plde.PCPlus4E[21] ;
 wire \rvcpu.dp.plde.PCPlus4E[22] ;
 wire \rvcpu.dp.plde.PCPlus4E[23] ;
 wire \rvcpu.dp.plde.PCPlus4E[24] ;
 wire \rvcpu.dp.plde.PCPlus4E[25] ;
 wire \rvcpu.dp.plde.PCPlus4E[26] ;
 wire \rvcpu.dp.plde.PCPlus4E[27] ;
 wire \rvcpu.dp.plde.PCPlus4E[28] ;
 wire \rvcpu.dp.plde.PCPlus4E[29] ;
 wire \rvcpu.dp.plde.PCPlus4E[2] ;
 wire \rvcpu.dp.plde.PCPlus4E[30] ;
 wire \rvcpu.dp.plde.PCPlus4E[31] ;
 wire \rvcpu.dp.plde.PCPlus4E[3] ;
 wire \rvcpu.dp.plde.PCPlus4E[4] ;
 wire \rvcpu.dp.plde.PCPlus4E[5] ;
 wire \rvcpu.dp.plde.PCPlus4E[6] ;
 wire \rvcpu.dp.plde.PCPlus4E[7] ;
 wire \rvcpu.dp.plde.PCPlus4E[8] ;
 wire \rvcpu.dp.plde.PCPlus4E[9] ;
 wire \rvcpu.dp.plde.RD1E[0] ;
 wire \rvcpu.dp.plde.RD1E[10] ;
 wire \rvcpu.dp.plde.RD1E[11] ;
 wire \rvcpu.dp.plde.RD1E[12] ;
 wire \rvcpu.dp.plde.RD1E[13] ;
 wire \rvcpu.dp.plde.RD1E[14] ;
 wire \rvcpu.dp.plde.RD1E[15] ;
 wire \rvcpu.dp.plde.RD1E[16] ;
 wire \rvcpu.dp.plde.RD1E[17] ;
 wire \rvcpu.dp.plde.RD1E[18] ;
 wire \rvcpu.dp.plde.RD1E[19] ;
 wire \rvcpu.dp.plde.RD1E[1] ;
 wire \rvcpu.dp.plde.RD1E[20] ;
 wire \rvcpu.dp.plde.RD1E[21] ;
 wire \rvcpu.dp.plde.RD1E[22] ;
 wire \rvcpu.dp.plde.RD1E[23] ;
 wire \rvcpu.dp.plde.RD1E[24] ;
 wire \rvcpu.dp.plde.RD1E[25] ;
 wire \rvcpu.dp.plde.RD1E[26] ;
 wire \rvcpu.dp.plde.RD1E[27] ;
 wire \rvcpu.dp.plde.RD1E[28] ;
 wire \rvcpu.dp.plde.RD1E[29] ;
 wire \rvcpu.dp.plde.RD1E[2] ;
 wire \rvcpu.dp.plde.RD1E[30] ;
 wire \rvcpu.dp.plde.RD1E[31] ;
 wire \rvcpu.dp.plde.RD1E[3] ;
 wire \rvcpu.dp.plde.RD1E[4] ;
 wire \rvcpu.dp.plde.RD1E[5] ;
 wire \rvcpu.dp.plde.RD1E[6] ;
 wire \rvcpu.dp.plde.RD1E[7] ;
 wire \rvcpu.dp.plde.RD1E[8] ;
 wire \rvcpu.dp.plde.RD1E[9] ;
 wire \rvcpu.dp.plde.RD2E[0] ;
 wire \rvcpu.dp.plde.RD2E[10] ;
 wire \rvcpu.dp.plde.RD2E[11] ;
 wire \rvcpu.dp.plde.RD2E[12] ;
 wire \rvcpu.dp.plde.RD2E[13] ;
 wire \rvcpu.dp.plde.RD2E[14] ;
 wire \rvcpu.dp.plde.RD2E[15] ;
 wire \rvcpu.dp.plde.RD2E[16] ;
 wire \rvcpu.dp.plde.RD2E[17] ;
 wire \rvcpu.dp.plde.RD2E[18] ;
 wire \rvcpu.dp.plde.RD2E[19] ;
 wire \rvcpu.dp.plde.RD2E[1] ;
 wire \rvcpu.dp.plde.RD2E[20] ;
 wire \rvcpu.dp.plde.RD2E[21] ;
 wire \rvcpu.dp.plde.RD2E[22] ;
 wire \rvcpu.dp.plde.RD2E[23] ;
 wire \rvcpu.dp.plde.RD2E[24] ;
 wire \rvcpu.dp.plde.RD2E[25] ;
 wire \rvcpu.dp.plde.RD2E[26] ;
 wire \rvcpu.dp.plde.RD2E[27] ;
 wire \rvcpu.dp.plde.RD2E[28] ;
 wire \rvcpu.dp.plde.RD2E[29] ;
 wire \rvcpu.dp.plde.RD2E[2] ;
 wire \rvcpu.dp.plde.RD2E[30] ;
 wire \rvcpu.dp.plde.RD2E[31] ;
 wire \rvcpu.dp.plde.RD2E[3] ;
 wire \rvcpu.dp.plde.RD2E[4] ;
 wire \rvcpu.dp.plde.RD2E[5] ;
 wire \rvcpu.dp.plde.RD2E[6] ;
 wire \rvcpu.dp.plde.RD2E[7] ;
 wire \rvcpu.dp.plde.RD2E[8] ;
 wire \rvcpu.dp.plde.RD2E[9] ;
 wire \rvcpu.dp.plde.RdE[0] ;
 wire \rvcpu.dp.plde.RdE[1] ;
 wire \rvcpu.dp.plde.RdE[2] ;
 wire \rvcpu.dp.plde.RdE[3] ;
 wire \rvcpu.dp.plde.RdE[4] ;
 wire \rvcpu.dp.plde.RegWriteE ;
 wire \rvcpu.dp.plde.ResultSrcE[1] ;
 wire \rvcpu.dp.plde.Rs1E[0] ;
 wire \rvcpu.dp.plde.Rs1E[1] ;
 wire \rvcpu.dp.plde.Rs1E[2] ;
 wire \rvcpu.dp.plde.Rs1E[3] ;
 wire \rvcpu.dp.plde.Rs1E[4] ;
 wire \rvcpu.dp.plde.Rs2E[0] ;
 wire \rvcpu.dp.plde.Rs2E[1] ;
 wire \rvcpu.dp.plde.Rs2E[2] ;
 wire \rvcpu.dp.plde.Rs2E[3] ;
 wire \rvcpu.dp.plde.Rs2E[4] ;
 wire \rvcpu.dp.plde.funct3E[0] ;
 wire \rvcpu.dp.plde.funct3E[1] ;
 wire \rvcpu.dp.plde.funct3E[2] ;
 wire \rvcpu.dp.plde.luiE ;
 wire \rvcpu.dp.plde.unsignE ;
 wire \rvcpu.dp.plem.ALUResultM[0] ;
 wire \rvcpu.dp.plem.ALUResultM[10] ;
 wire \rvcpu.dp.plem.ALUResultM[11] ;
 wire \rvcpu.dp.plem.ALUResultM[12] ;
 wire \rvcpu.dp.plem.ALUResultM[13] ;
 wire \rvcpu.dp.plem.ALUResultM[14] ;
 wire \rvcpu.dp.plem.ALUResultM[15] ;
 wire \rvcpu.dp.plem.ALUResultM[16] ;
 wire \rvcpu.dp.plem.ALUResultM[17] ;
 wire \rvcpu.dp.plem.ALUResultM[18] ;
 wire \rvcpu.dp.plem.ALUResultM[19] ;
 wire \rvcpu.dp.plem.ALUResultM[1] ;
 wire \rvcpu.dp.plem.ALUResultM[20] ;
 wire \rvcpu.dp.plem.ALUResultM[21] ;
 wire \rvcpu.dp.plem.ALUResultM[22] ;
 wire \rvcpu.dp.plem.ALUResultM[23] ;
 wire \rvcpu.dp.plem.ALUResultM[24] ;
 wire \rvcpu.dp.plem.ALUResultM[25] ;
 wire \rvcpu.dp.plem.ALUResultM[26] ;
 wire \rvcpu.dp.plem.ALUResultM[27] ;
 wire \rvcpu.dp.plem.ALUResultM[28] ;
 wire \rvcpu.dp.plem.ALUResultM[29] ;
 wire \rvcpu.dp.plem.ALUResultM[2] ;
 wire \rvcpu.dp.plem.ALUResultM[30] ;
 wire \rvcpu.dp.plem.ALUResultM[31] ;
 wire \rvcpu.dp.plem.ALUResultM[3] ;
 wire \rvcpu.dp.plem.ALUResultM[4] ;
 wire \rvcpu.dp.plem.ALUResultM[5] ;
 wire \rvcpu.dp.plem.ALUResultM[6] ;
 wire \rvcpu.dp.plem.ALUResultM[7] ;
 wire \rvcpu.dp.plem.ALUResultM[8] ;
 wire \rvcpu.dp.plem.ALUResultM[9] ;
 wire \rvcpu.dp.plem.MemWriteM ;
 wire \rvcpu.dp.plem.PCPlus4M[0] ;
 wire \rvcpu.dp.plem.PCPlus4M[10] ;
 wire \rvcpu.dp.plem.PCPlus4M[11] ;
 wire \rvcpu.dp.plem.PCPlus4M[12] ;
 wire \rvcpu.dp.plem.PCPlus4M[13] ;
 wire \rvcpu.dp.plem.PCPlus4M[14] ;
 wire \rvcpu.dp.plem.PCPlus4M[15] ;
 wire \rvcpu.dp.plem.PCPlus4M[16] ;
 wire \rvcpu.dp.plem.PCPlus4M[17] ;
 wire \rvcpu.dp.plem.PCPlus4M[18] ;
 wire \rvcpu.dp.plem.PCPlus4M[19] ;
 wire \rvcpu.dp.plem.PCPlus4M[1] ;
 wire \rvcpu.dp.plem.PCPlus4M[20] ;
 wire \rvcpu.dp.plem.PCPlus4M[21] ;
 wire \rvcpu.dp.plem.PCPlus4M[22] ;
 wire \rvcpu.dp.plem.PCPlus4M[23] ;
 wire \rvcpu.dp.plem.PCPlus4M[24] ;
 wire \rvcpu.dp.plem.PCPlus4M[25] ;
 wire \rvcpu.dp.plem.PCPlus4M[26] ;
 wire \rvcpu.dp.plem.PCPlus4M[27] ;
 wire \rvcpu.dp.plem.PCPlus4M[28] ;
 wire \rvcpu.dp.plem.PCPlus4M[29] ;
 wire \rvcpu.dp.plem.PCPlus4M[2] ;
 wire \rvcpu.dp.plem.PCPlus4M[30] ;
 wire \rvcpu.dp.plem.PCPlus4M[31] ;
 wire \rvcpu.dp.plem.PCPlus4M[3] ;
 wire \rvcpu.dp.plem.PCPlus4M[4] ;
 wire \rvcpu.dp.plem.PCPlus4M[5] ;
 wire \rvcpu.dp.plem.PCPlus4M[6] ;
 wire \rvcpu.dp.plem.PCPlus4M[7] ;
 wire \rvcpu.dp.plem.PCPlus4M[8] ;
 wire \rvcpu.dp.plem.PCPlus4M[9] ;
 wire \rvcpu.dp.plem.RdM[0] ;
 wire \rvcpu.dp.plem.RdM[1] ;
 wire \rvcpu.dp.plem.RdM[2] ;
 wire \rvcpu.dp.plem.RdM[3] ;
 wire \rvcpu.dp.plem.RdM[4] ;
 wire \rvcpu.dp.plem.RegWriteM ;
 wire \rvcpu.dp.plem.ResultSrcM[0] ;
 wire \rvcpu.dp.plem.ResultSrcM[1] ;
 wire \rvcpu.dp.plem.WriteDataM[0] ;
 wire \rvcpu.dp.plem.WriteDataM[10] ;
 wire \rvcpu.dp.plem.WriteDataM[11] ;
 wire \rvcpu.dp.plem.WriteDataM[12] ;
 wire \rvcpu.dp.plem.WriteDataM[13] ;
 wire \rvcpu.dp.plem.WriteDataM[14] ;
 wire \rvcpu.dp.plem.WriteDataM[15] ;
 wire \rvcpu.dp.plem.WriteDataM[16] ;
 wire \rvcpu.dp.plem.WriteDataM[17] ;
 wire \rvcpu.dp.plem.WriteDataM[18] ;
 wire \rvcpu.dp.plem.WriteDataM[19] ;
 wire \rvcpu.dp.plem.WriteDataM[1] ;
 wire \rvcpu.dp.plem.WriteDataM[20] ;
 wire \rvcpu.dp.plem.WriteDataM[21] ;
 wire \rvcpu.dp.plem.WriteDataM[22] ;
 wire \rvcpu.dp.plem.WriteDataM[23] ;
 wire \rvcpu.dp.plem.WriteDataM[24] ;
 wire \rvcpu.dp.plem.WriteDataM[25] ;
 wire \rvcpu.dp.plem.WriteDataM[26] ;
 wire \rvcpu.dp.plem.WriteDataM[27] ;
 wire \rvcpu.dp.plem.WriteDataM[28] ;
 wire \rvcpu.dp.plem.WriteDataM[29] ;
 wire \rvcpu.dp.plem.WriteDataM[2] ;
 wire \rvcpu.dp.plem.WriteDataM[30] ;
 wire \rvcpu.dp.plem.WriteDataM[31] ;
 wire \rvcpu.dp.plem.WriteDataM[3] ;
 wire \rvcpu.dp.plem.WriteDataM[4] ;
 wire \rvcpu.dp.plem.WriteDataM[5] ;
 wire \rvcpu.dp.plem.WriteDataM[6] ;
 wire \rvcpu.dp.plem.WriteDataM[7] ;
 wire \rvcpu.dp.plem.WriteDataM[8] ;
 wire \rvcpu.dp.plem.WriteDataM[9] ;
 wire \rvcpu.dp.plem.funct3M[0] ;
 wire \rvcpu.dp.plem.funct3M[1] ;
 wire \rvcpu.dp.plem.funct3M[2] ;
 wire \rvcpu.dp.plem.lAuiPCM[0] ;
 wire \rvcpu.dp.plem.lAuiPCM[10] ;
 wire \rvcpu.dp.plem.lAuiPCM[11] ;
 wire \rvcpu.dp.plem.lAuiPCM[12] ;
 wire \rvcpu.dp.plem.lAuiPCM[13] ;
 wire \rvcpu.dp.plem.lAuiPCM[14] ;
 wire \rvcpu.dp.plem.lAuiPCM[15] ;
 wire \rvcpu.dp.plem.lAuiPCM[16] ;
 wire \rvcpu.dp.plem.lAuiPCM[17] ;
 wire \rvcpu.dp.plem.lAuiPCM[18] ;
 wire \rvcpu.dp.plem.lAuiPCM[19] ;
 wire \rvcpu.dp.plem.lAuiPCM[1] ;
 wire \rvcpu.dp.plem.lAuiPCM[20] ;
 wire \rvcpu.dp.plem.lAuiPCM[21] ;
 wire \rvcpu.dp.plem.lAuiPCM[22] ;
 wire \rvcpu.dp.plem.lAuiPCM[23] ;
 wire \rvcpu.dp.plem.lAuiPCM[24] ;
 wire \rvcpu.dp.plem.lAuiPCM[25] ;
 wire \rvcpu.dp.plem.lAuiPCM[26] ;
 wire \rvcpu.dp.plem.lAuiPCM[27] ;
 wire \rvcpu.dp.plem.lAuiPCM[28] ;
 wire \rvcpu.dp.plem.lAuiPCM[29] ;
 wire \rvcpu.dp.plem.lAuiPCM[2] ;
 wire \rvcpu.dp.plem.lAuiPCM[30] ;
 wire \rvcpu.dp.plem.lAuiPCM[31] ;
 wire \rvcpu.dp.plem.lAuiPCM[3] ;
 wire \rvcpu.dp.plem.lAuiPCM[4] ;
 wire \rvcpu.dp.plem.lAuiPCM[5] ;
 wire \rvcpu.dp.plem.lAuiPCM[6] ;
 wire \rvcpu.dp.plem.lAuiPCM[7] ;
 wire \rvcpu.dp.plem.lAuiPCM[8] ;
 wire \rvcpu.dp.plem.lAuiPCM[9] ;
 wire \rvcpu.dp.plfd.InstrD[0] ;
 wire \rvcpu.dp.plfd.InstrD[10] ;
 wire \rvcpu.dp.plfd.InstrD[11] ;
 wire \rvcpu.dp.plfd.InstrD[12] ;
 wire \rvcpu.dp.plfd.InstrD[13] ;
 wire \rvcpu.dp.plfd.InstrD[14] ;
 wire \rvcpu.dp.plfd.InstrD[15] ;
 wire \rvcpu.dp.plfd.InstrD[16] ;
 wire \rvcpu.dp.plfd.InstrD[17] ;
 wire \rvcpu.dp.plfd.InstrD[18] ;
 wire \rvcpu.dp.plfd.InstrD[19] ;
 wire \rvcpu.dp.plfd.InstrD[20] ;
 wire \rvcpu.dp.plfd.InstrD[21] ;
 wire \rvcpu.dp.plfd.InstrD[22] ;
 wire \rvcpu.dp.plfd.InstrD[23] ;
 wire \rvcpu.dp.plfd.InstrD[24] ;
 wire \rvcpu.dp.plfd.InstrD[25] ;
 wire \rvcpu.dp.plfd.InstrD[26] ;
 wire \rvcpu.dp.plfd.InstrD[27] ;
 wire \rvcpu.dp.plfd.InstrD[28] ;
 wire \rvcpu.dp.plfd.InstrD[29] ;
 wire \rvcpu.dp.plfd.InstrD[2] ;
 wire \rvcpu.dp.plfd.InstrD[31] ;
 wire \rvcpu.dp.plfd.InstrD[3] ;
 wire \rvcpu.dp.plfd.InstrD[4] ;
 wire \rvcpu.dp.plfd.InstrD[6] ;
 wire \rvcpu.dp.plfd.InstrD[7] ;
 wire \rvcpu.dp.plfd.InstrD[8] ;
 wire \rvcpu.dp.plfd.InstrD[9] ;
 wire \rvcpu.dp.plfd.PCD[0] ;
 wire \rvcpu.dp.plfd.PCD[10] ;
 wire \rvcpu.dp.plfd.PCD[11] ;
 wire \rvcpu.dp.plfd.PCD[12] ;
 wire \rvcpu.dp.plfd.PCD[13] ;
 wire \rvcpu.dp.plfd.PCD[14] ;
 wire \rvcpu.dp.plfd.PCD[15] ;
 wire \rvcpu.dp.plfd.PCD[16] ;
 wire \rvcpu.dp.plfd.PCD[17] ;
 wire \rvcpu.dp.plfd.PCD[18] ;
 wire \rvcpu.dp.plfd.PCD[19] ;
 wire \rvcpu.dp.plfd.PCD[1] ;
 wire \rvcpu.dp.plfd.PCD[20] ;
 wire \rvcpu.dp.plfd.PCD[21] ;
 wire \rvcpu.dp.plfd.PCD[22] ;
 wire \rvcpu.dp.plfd.PCD[23] ;
 wire \rvcpu.dp.plfd.PCD[24] ;
 wire \rvcpu.dp.plfd.PCD[25] ;
 wire \rvcpu.dp.plfd.PCD[26] ;
 wire \rvcpu.dp.plfd.PCD[27] ;
 wire \rvcpu.dp.plfd.PCD[28] ;
 wire \rvcpu.dp.plfd.PCD[29] ;
 wire \rvcpu.dp.plfd.PCD[2] ;
 wire \rvcpu.dp.plfd.PCD[30] ;
 wire \rvcpu.dp.plfd.PCD[31] ;
 wire \rvcpu.dp.plfd.PCD[3] ;
 wire \rvcpu.dp.plfd.PCD[4] ;
 wire \rvcpu.dp.plfd.PCD[5] ;
 wire \rvcpu.dp.plfd.PCD[6] ;
 wire \rvcpu.dp.plfd.PCD[7] ;
 wire \rvcpu.dp.plfd.PCD[8] ;
 wire \rvcpu.dp.plfd.PCD[9] ;
 wire \rvcpu.dp.plfd.PCPlus4D[10] ;
 wire \rvcpu.dp.plfd.PCPlus4D[11] ;
 wire \rvcpu.dp.plfd.PCPlus4D[12] ;
 wire \rvcpu.dp.plfd.PCPlus4D[13] ;
 wire \rvcpu.dp.plfd.PCPlus4D[14] ;
 wire \rvcpu.dp.plfd.PCPlus4D[15] ;
 wire \rvcpu.dp.plfd.PCPlus4D[16] ;
 wire \rvcpu.dp.plfd.PCPlus4D[17] ;
 wire \rvcpu.dp.plfd.PCPlus4D[18] ;
 wire \rvcpu.dp.plfd.PCPlus4D[19] ;
 wire \rvcpu.dp.plfd.PCPlus4D[20] ;
 wire \rvcpu.dp.plfd.PCPlus4D[21] ;
 wire \rvcpu.dp.plfd.PCPlus4D[22] ;
 wire \rvcpu.dp.plfd.PCPlus4D[23] ;
 wire \rvcpu.dp.plfd.PCPlus4D[24] ;
 wire \rvcpu.dp.plfd.PCPlus4D[25] ;
 wire \rvcpu.dp.plfd.PCPlus4D[26] ;
 wire \rvcpu.dp.plfd.PCPlus4D[27] ;
 wire \rvcpu.dp.plfd.PCPlus4D[28] ;
 wire \rvcpu.dp.plfd.PCPlus4D[29] ;
 wire \rvcpu.dp.plfd.PCPlus4D[2] ;
 wire \rvcpu.dp.plfd.PCPlus4D[30] ;
 wire \rvcpu.dp.plfd.PCPlus4D[31] ;
 wire \rvcpu.dp.plfd.PCPlus4D[3] ;
 wire \rvcpu.dp.plfd.PCPlus4D[4] ;
 wire \rvcpu.dp.plfd.PCPlus4D[5] ;
 wire \rvcpu.dp.plfd.PCPlus4D[6] ;
 wire \rvcpu.dp.plfd.PCPlus4D[7] ;
 wire \rvcpu.dp.plfd.PCPlus4D[8] ;
 wire \rvcpu.dp.plfd.PCPlus4D[9] ;
 wire \rvcpu.dp.plmw.ALUResultW[0] ;
 wire \rvcpu.dp.plmw.ALUResultW[10] ;
 wire \rvcpu.dp.plmw.ALUResultW[11] ;
 wire \rvcpu.dp.plmw.ALUResultW[12] ;
 wire \rvcpu.dp.plmw.ALUResultW[13] ;
 wire \rvcpu.dp.plmw.ALUResultW[14] ;
 wire \rvcpu.dp.plmw.ALUResultW[15] ;
 wire \rvcpu.dp.plmw.ALUResultW[16] ;
 wire \rvcpu.dp.plmw.ALUResultW[17] ;
 wire \rvcpu.dp.plmw.ALUResultW[18] ;
 wire \rvcpu.dp.plmw.ALUResultW[19] ;
 wire \rvcpu.dp.plmw.ALUResultW[1] ;
 wire \rvcpu.dp.plmw.ALUResultW[20] ;
 wire \rvcpu.dp.plmw.ALUResultW[21] ;
 wire \rvcpu.dp.plmw.ALUResultW[22] ;
 wire \rvcpu.dp.plmw.ALUResultW[23] ;
 wire \rvcpu.dp.plmw.ALUResultW[24] ;
 wire \rvcpu.dp.plmw.ALUResultW[25] ;
 wire \rvcpu.dp.plmw.ALUResultW[26] ;
 wire \rvcpu.dp.plmw.ALUResultW[27] ;
 wire \rvcpu.dp.plmw.ALUResultW[28] ;
 wire \rvcpu.dp.plmw.ALUResultW[29] ;
 wire \rvcpu.dp.plmw.ALUResultW[2] ;
 wire \rvcpu.dp.plmw.ALUResultW[30] ;
 wire \rvcpu.dp.plmw.ALUResultW[31] ;
 wire \rvcpu.dp.plmw.ALUResultW[3] ;
 wire \rvcpu.dp.plmw.ALUResultW[4] ;
 wire \rvcpu.dp.plmw.ALUResultW[5] ;
 wire \rvcpu.dp.plmw.ALUResultW[6] ;
 wire \rvcpu.dp.plmw.ALUResultW[7] ;
 wire \rvcpu.dp.plmw.ALUResultW[8] ;
 wire \rvcpu.dp.plmw.ALUResultW[9] ;
 wire \rvcpu.dp.plmw.PCPlus4W[0] ;
 wire \rvcpu.dp.plmw.PCPlus4W[10] ;
 wire \rvcpu.dp.plmw.PCPlus4W[11] ;
 wire \rvcpu.dp.plmw.PCPlus4W[12] ;
 wire \rvcpu.dp.plmw.PCPlus4W[13] ;
 wire \rvcpu.dp.plmw.PCPlus4W[14] ;
 wire \rvcpu.dp.plmw.PCPlus4W[15] ;
 wire \rvcpu.dp.plmw.PCPlus4W[16] ;
 wire \rvcpu.dp.plmw.PCPlus4W[17] ;
 wire \rvcpu.dp.plmw.PCPlus4W[18] ;
 wire \rvcpu.dp.plmw.PCPlus4W[19] ;
 wire \rvcpu.dp.plmw.PCPlus4W[1] ;
 wire \rvcpu.dp.plmw.PCPlus4W[20] ;
 wire \rvcpu.dp.plmw.PCPlus4W[21] ;
 wire \rvcpu.dp.plmw.PCPlus4W[22] ;
 wire \rvcpu.dp.plmw.PCPlus4W[23] ;
 wire \rvcpu.dp.plmw.PCPlus4W[24] ;
 wire \rvcpu.dp.plmw.PCPlus4W[25] ;
 wire \rvcpu.dp.plmw.PCPlus4W[26] ;
 wire \rvcpu.dp.plmw.PCPlus4W[27] ;
 wire \rvcpu.dp.plmw.PCPlus4W[28] ;
 wire \rvcpu.dp.plmw.PCPlus4W[29] ;
 wire \rvcpu.dp.plmw.PCPlus4W[2] ;
 wire \rvcpu.dp.plmw.PCPlus4W[30] ;
 wire \rvcpu.dp.plmw.PCPlus4W[31] ;
 wire \rvcpu.dp.plmw.PCPlus4W[3] ;
 wire \rvcpu.dp.plmw.PCPlus4W[4] ;
 wire \rvcpu.dp.plmw.PCPlus4W[5] ;
 wire \rvcpu.dp.plmw.PCPlus4W[6] ;
 wire \rvcpu.dp.plmw.PCPlus4W[7] ;
 wire \rvcpu.dp.plmw.PCPlus4W[8] ;
 wire \rvcpu.dp.plmw.PCPlus4W[9] ;
 wire \rvcpu.dp.plmw.RdW[0] ;
 wire \rvcpu.dp.plmw.RdW[1] ;
 wire \rvcpu.dp.plmw.RdW[2] ;
 wire \rvcpu.dp.plmw.RdW[3] ;
 wire \rvcpu.dp.plmw.RdW[4] ;
 wire \rvcpu.dp.plmw.ReadDataW[0] ;
 wire \rvcpu.dp.plmw.ReadDataW[10] ;
 wire \rvcpu.dp.plmw.ReadDataW[11] ;
 wire \rvcpu.dp.plmw.ReadDataW[12] ;
 wire \rvcpu.dp.plmw.ReadDataW[13] ;
 wire \rvcpu.dp.plmw.ReadDataW[14] ;
 wire \rvcpu.dp.plmw.ReadDataW[15] ;
 wire \rvcpu.dp.plmw.ReadDataW[16] ;
 wire \rvcpu.dp.plmw.ReadDataW[17] ;
 wire \rvcpu.dp.plmw.ReadDataW[18] ;
 wire \rvcpu.dp.plmw.ReadDataW[19] ;
 wire \rvcpu.dp.plmw.ReadDataW[1] ;
 wire \rvcpu.dp.plmw.ReadDataW[20] ;
 wire \rvcpu.dp.plmw.ReadDataW[21] ;
 wire \rvcpu.dp.plmw.ReadDataW[22] ;
 wire \rvcpu.dp.plmw.ReadDataW[23] ;
 wire \rvcpu.dp.plmw.ReadDataW[24] ;
 wire \rvcpu.dp.plmw.ReadDataW[25] ;
 wire \rvcpu.dp.plmw.ReadDataW[26] ;
 wire \rvcpu.dp.plmw.ReadDataW[27] ;
 wire \rvcpu.dp.plmw.ReadDataW[28] ;
 wire \rvcpu.dp.plmw.ReadDataW[29] ;
 wire \rvcpu.dp.plmw.ReadDataW[2] ;
 wire \rvcpu.dp.plmw.ReadDataW[30] ;
 wire \rvcpu.dp.plmw.ReadDataW[31] ;
 wire \rvcpu.dp.plmw.ReadDataW[3] ;
 wire \rvcpu.dp.plmw.ReadDataW[4] ;
 wire \rvcpu.dp.plmw.ReadDataW[5] ;
 wire \rvcpu.dp.plmw.ReadDataW[6] ;
 wire \rvcpu.dp.plmw.ReadDataW[7] ;
 wire \rvcpu.dp.plmw.ReadDataW[8] ;
 wire \rvcpu.dp.plmw.ReadDataW[9] ;
 wire \rvcpu.dp.plmw.RegWriteW ;
 wire \rvcpu.dp.plmw.ResultSrcW[0] ;
 wire \rvcpu.dp.plmw.ResultSrcW[1] ;
 wire \rvcpu.dp.plmw.lAuiPCW[0] ;
 wire \rvcpu.dp.plmw.lAuiPCW[10] ;
 wire \rvcpu.dp.plmw.lAuiPCW[11] ;
 wire \rvcpu.dp.plmw.lAuiPCW[12] ;
 wire \rvcpu.dp.plmw.lAuiPCW[13] ;
 wire \rvcpu.dp.plmw.lAuiPCW[14] ;
 wire \rvcpu.dp.plmw.lAuiPCW[15] ;
 wire \rvcpu.dp.plmw.lAuiPCW[16] ;
 wire \rvcpu.dp.plmw.lAuiPCW[17] ;
 wire \rvcpu.dp.plmw.lAuiPCW[18] ;
 wire \rvcpu.dp.plmw.lAuiPCW[19] ;
 wire \rvcpu.dp.plmw.lAuiPCW[1] ;
 wire \rvcpu.dp.plmw.lAuiPCW[20] ;
 wire \rvcpu.dp.plmw.lAuiPCW[21] ;
 wire \rvcpu.dp.plmw.lAuiPCW[22] ;
 wire \rvcpu.dp.plmw.lAuiPCW[23] ;
 wire \rvcpu.dp.plmw.lAuiPCW[24] ;
 wire \rvcpu.dp.plmw.lAuiPCW[25] ;
 wire \rvcpu.dp.plmw.lAuiPCW[26] ;
 wire \rvcpu.dp.plmw.lAuiPCW[27] ;
 wire \rvcpu.dp.plmw.lAuiPCW[28] ;
 wire \rvcpu.dp.plmw.lAuiPCW[29] ;
 wire \rvcpu.dp.plmw.lAuiPCW[2] ;
 wire \rvcpu.dp.plmw.lAuiPCW[30] ;
 wire \rvcpu.dp.plmw.lAuiPCW[31] ;
 wire \rvcpu.dp.plmw.lAuiPCW[3] ;
 wire \rvcpu.dp.plmw.lAuiPCW[4] ;
 wire \rvcpu.dp.plmw.lAuiPCW[5] ;
 wire \rvcpu.dp.plmw.lAuiPCW[6] ;
 wire \rvcpu.dp.plmw.lAuiPCW[7] ;
 wire \rvcpu.dp.plmw.lAuiPCW[8] ;
 wire \rvcpu.dp.plmw.lAuiPCW[9] ;
 wire \rvcpu.dp.rf.reg_file_arr[0][0] ;
 wire \rvcpu.dp.rf.reg_file_arr[0][10] ;
 wire \rvcpu.dp.rf.reg_file_arr[0][11] ;
 wire \rvcpu.dp.rf.reg_file_arr[0][12] ;
 wire \rvcpu.dp.rf.reg_file_arr[0][13] ;
 wire \rvcpu.dp.rf.reg_file_arr[0][14] ;
 wire \rvcpu.dp.rf.reg_file_arr[0][15] ;
 wire \rvcpu.dp.rf.reg_file_arr[0][16] ;
 wire \rvcpu.dp.rf.reg_file_arr[0][17] ;
 wire \rvcpu.dp.rf.reg_file_arr[0][18] ;
 wire \rvcpu.dp.rf.reg_file_arr[0][19] ;
 wire \rvcpu.dp.rf.reg_file_arr[0][1] ;
 wire \rvcpu.dp.rf.reg_file_arr[0][20] ;
 wire \rvcpu.dp.rf.reg_file_arr[0][21] ;
 wire \rvcpu.dp.rf.reg_file_arr[0][22] ;
 wire \rvcpu.dp.rf.reg_file_arr[0][23] ;
 wire \rvcpu.dp.rf.reg_file_arr[0][24] ;
 wire \rvcpu.dp.rf.reg_file_arr[0][25] ;
 wire \rvcpu.dp.rf.reg_file_arr[0][26] ;
 wire \rvcpu.dp.rf.reg_file_arr[0][27] ;
 wire \rvcpu.dp.rf.reg_file_arr[0][28] ;
 wire \rvcpu.dp.rf.reg_file_arr[0][29] ;
 wire \rvcpu.dp.rf.reg_file_arr[0][2] ;
 wire \rvcpu.dp.rf.reg_file_arr[0][30] ;
 wire \rvcpu.dp.rf.reg_file_arr[0][31] ;
 wire \rvcpu.dp.rf.reg_file_arr[0][3] ;
 wire \rvcpu.dp.rf.reg_file_arr[0][4] ;
 wire \rvcpu.dp.rf.reg_file_arr[0][5] ;
 wire \rvcpu.dp.rf.reg_file_arr[0][6] ;
 wire \rvcpu.dp.rf.reg_file_arr[0][7] ;
 wire \rvcpu.dp.rf.reg_file_arr[0][8] ;
 wire \rvcpu.dp.rf.reg_file_arr[0][9] ;
 wire \rvcpu.dp.rf.reg_file_arr[10][0] ;
 wire \rvcpu.dp.rf.reg_file_arr[10][10] ;
 wire \rvcpu.dp.rf.reg_file_arr[10][11] ;
 wire \rvcpu.dp.rf.reg_file_arr[10][12] ;
 wire \rvcpu.dp.rf.reg_file_arr[10][13] ;
 wire \rvcpu.dp.rf.reg_file_arr[10][14] ;
 wire \rvcpu.dp.rf.reg_file_arr[10][15] ;
 wire \rvcpu.dp.rf.reg_file_arr[10][16] ;
 wire \rvcpu.dp.rf.reg_file_arr[10][17] ;
 wire \rvcpu.dp.rf.reg_file_arr[10][18] ;
 wire \rvcpu.dp.rf.reg_file_arr[10][19] ;
 wire \rvcpu.dp.rf.reg_file_arr[10][1] ;
 wire \rvcpu.dp.rf.reg_file_arr[10][20] ;
 wire \rvcpu.dp.rf.reg_file_arr[10][21] ;
 wire \rvcpu.dp.rf.reg_file_arr[10][22] ;
 wire \rvcpu.dp.rf.reg_file_arr[10][23] ;
 wire \rvcpu.dp.rf.reg_file_arr[10][24] ;
 wire \rvcpu.dp.rf.reg_file_arr[10][25] ;
 wire \rvcpu.dp.rf.reg_file_arr[10][26] ;
 wire \rvcpu.dp.rf.reg_file_arr[10][27] ;
 wire \rvcpu.dp.rf.reg_file_arr[10][28] ;
 wire \rvcpu.dp.rf.reg_file_arr[10][29] ;
 wire \rvcpu.dp.rf.reg_file_arr[10][2] ;
 wire \rvcpu.dp.rf.reg_file_arr[10][30] ;
 wire \rvcpu.dp.rf.reg_file_arr[10][31] ;
 wire \rvcpu.dp.rf.reg_file_arr[10][3] ;
 wire \rvcpu.dp.rf.reg_file_arr[10][4] ;
 wire \rvcpu.dp.rf.reg_file_arr[10][5] ;
 wire \rvcpu.dp.rf.reg_file_arr[10][6] ;
 wire \rvcpu.dp.rf.reg_file_arr[10][7] ;
 wire \rvcpu.dp.rf.reg_file_arr[10][8] ;
 wire \rvcpu.dp.rf.reg_file_arr[10][9] ;
 wire \rvcpu.dp.rf.reg_file_arr[11][0] ;
 wire \rvcpu.dp.rf.reg_file_arr[11][10] ;
 wire \rvcpu.dp.rf.reg_file_arr[11][11] ;
 wire \rvcpu.dp.rf.reg_file_arr[11][12] ;
 wire \rvcpu.dp.rf.reg_file_arr[11][13] ;
 wire \rvcpu.dp.rf.reg_file_arr[11][14] ;
 wire \rvcpu.dp.rf.reg_file_arr[11][15] ;
 wire \rvcpu.dp.rf.reg_file_arr[11][16] ;
 wire \rvcpu.dp.rf.reg_file_arr[11][17] ;
 wire \rvcpu.dp.rf.reg_file_arr[11][18] ;
 wire \rvcpu.dp.rf.reg_file_arr[11][19] ;
 wire \rvcpu.dp.rf.reg_file_arr[11][1] ;
 wire \rvcpu.dp.rf.reg_file_arr[11][20] ;
 wire \rvcpu.dp.rf.reg_file_arr[11][21] ;
 wire \rvcpu.dp.rf.reg_file_arr[11][22] ;
 wire \rvcpu.dp.rf.reg_file_arr[11][23] ;
 wire \rvcpu.dp.rf.reg_file_arr[11][24] ;
 wire \rvcpu.dp.rf.reg_file_arr[11][25] ;
 wire \rvcpu.dp.rf.reg_file_arr[11][26] ;
 wire \rvcpu.dp.rf.reg_file_arr[11][27] ;
 wire \rvcpu.dp.rf.reg_file_arr[11][28] ;
 wire \rvcpu.dp.rf.reg_file_arr[11][29] ;
 wire \rvcpu.dp.rf.reg_file_arr[11][2] ;
 wire \rvcpu.dp.rf.reg_file_arr[11][30] ;
 wire \rvcpu.dp.rf.reg_file_arr[11][31] ;
 wire \rvcpu.dp.rf.reg_file_arr[11][3] ;
 wire \rvcpu.dp.rf.reg_file_arr[11][4] ;
 wire \rvcpu.dp.rf.reg_file_arr[11][5] ;
 wire \rvcpu.dp.rf.reg_file_arr[11][6] ;
 wire \rvcpu.dp.rf.reg_file_arr[11][7] ;
 wire \rvcpu.dp.rf.reg_file_arr[11][8] ;
 wire \rvcpu.dp.rf.reg_file_arr[11][9] ;
 wire \rvcpu.dp.rf.reg_file_arr[12][0] ;
 wire \rvcpu.dp.rf.reg_file_arr[12][10] ;
 wire \rvcpu.dp.rf.reg_file_arr[12][11] ;
 wire \rvcpu.dp.rf.reg_file_arr[12][12] ;
 wire \rvcpu.dp.rf.reg_file_arr[12][13] ;
 wire \rvcpu.dp.rf.reg_file_arr[12][14] ;
 wire \rvcpu.dp.rf.reg_file_arr[12][15] ;
 wire \rvcpu.dp.rf.reg_file_arr[12][16] ;
 wire \rvcpu.dp.rf.reg_file_arr[12][17] ;
 wire \rvcpu.dp.rf.reg_file_arr[12][18] ;
 wire \rvcpu.dp.rf.reg_file_arr[12][19] ;
 wire \rvcpu.dp.rf.reg_file_arr[12][1] ;
 wire \rvcpu.dp.rf.reg_file_arr[12][20] ;
 wire \rvcpu.dp.rf.reg_file_arr[12][21] ;
 wire \rvcpu.dp.rf.reg_file_arr[12][22] ;
 wire \rvcpu.dp.rf.reg_file_arr[12][23] ;
 wire \rvcpu.dp.rf.reg_file_arr[12][24] ;
 wire \rvcpu.dp.rf.reg_file_arr[12][25] ;
 wire \rvcpu.dp.rf.reg_file_arr[12][26] ;
 wire \rvcpu.dp.rf.reg_file_arr[12][27] ;
 wire \rvcpu.dp.rf.reg_file_arr[12][28] ;
 wire \rvcpu.dp.rf.reg_file_arr[12][29] ;
 wire \rvcpu.dp.rf.reg_file_arr[12][2] ;
 wire \rvcpu.dp.rf.reg_file_arr[12][30] ;
 wire \rvcpu.dp.rf.reg_file_arr[12][31] ;
 wire \rvcpu.dp.rf.reg_file_arr[12][3] ;
 wire \rvcpu.dp.rf.reg_file_arr[12][4] ;
 wire \rvcpu.dp.rf.reg_file_arr[12][5] ;
 wire \rvcpu.dp.rf.reg_file_arr[12][6] ;
 wire \rvcpu.dp.rf.reg_file_arr[12][7] ;
 wire \rvcpu.dp.rf.reg_file_arr[12][8] ;
 wire \rvcpu.dp.rf.reg_file_arr[12][9] ;
 wire \rvcpu.dp.rf.reg_file_arr[13][0] ;
 wire \rvcpu.dp.rf.reg_file_arr[13][10] ;
 wire \rvcpu.dp.rf.reg_file_arr[13][11] ;
 wire \rvcpu.dp.rf.reg_file_arr[13][12] ;
 wire \rvcpu.dp.rf.reg_file_arr[13][13] ;
 wire \rvcpu.dp.rf.reg_file_arr[13][14] ;
 wire \rvcpu.dp.rf.reg_file_arr[13][15] ;
 wire \rvcpu.dp.rf.reg_file_arr[13][16] ;
 wire \rvcpu.dp.rf.reg_file_arr[13][17] ;
 wire \rvcpu.dp.rf.reg_file_arr[13][18] ;
 wire \rvcpu.dp.rf.reg_file_arr[13][19] ;
 wire \rvcpu.dp.rf.reg_file_arr[13][1] ;
 wire \rvcpu.dp.rf.reg_file_arr[13][20] ;
 wire \rvcpu.dp.rf.reg_file_arr[13][21] ;
 wire \rvcpu.dp.rf.reg_file_arr[13][22] ;
 wire \rvcpu.dp.rf.reg_file_arr[13][23] ;
 wire \rvcpu.dp.rf.reg_file_arr[13][24] ;
 wire \rvcpu.dp.rf.reg_file_arr[13][25] ;
 wire \rvcpu.dp.rf.reg_file_arr[13][26] ;
 wire \rvcpu.dp.rf.reg_file_arr[13][27] ;
 wire \rvcpu.dp.rf.reg_file_arr[13][28] ;
 wire \rvcpu.dp.rf.reg_file_arr[13][29] ;
 wire \rvcpu.dp.rf.reg_file_arr[13][2] ;
 wire \rvcpu.dp.rf.reg_file_arr[13][30] ;
 wire \rvcpu.dp.rf.reg_file_arr[13][31] ;
 wire \rvcpu.dp.rf.reg_file_arr[13][3] ;
 wire \rvcpu.dp.rf.reg_file_arr[13][4] ;
 wire \rvcpu.dp.rf.reg_file_arr[13][5] ;
 wire \rvcpu.dp.rf.reg_file_arr[13][6] ;
 wire \rvcpu.dp.rf.reg_file_arr[13][7] ;
 wire \rvcpu.dp.rf.reg_file_arr[13][8] ;
 wire \rvcpu.dp.rf.reg_file_arr[13][9] ;
 wire \rvcpu.dp.rf.reg_file_arr[14][0] ;
 wire \rvcpu.dp.rf.reg_file_arr[14][10] ;
 wire \rvcpu.dp.rf.reg_file_arr[14][11] ;
 wire \rvcpu.dp.rf.reg_file_arr[14][12] ;
 wire \rvcpu.dp.rf.reg_file_arr[14][13] ;
 wire \rvcpu.dp.rf.reg_file_arr[14][14] ;
 wire \rvcpu.dp.rf.reg_file_arr[14][15] ;
 wire \rvcpu.dp.rf.reg_file_arr[14][16] ;
 wire \rvcpu.dp.rf.reg_file_arr[14][17] ;
 wire \rvcpu.dp.rf.reg_file_arr[14][18] ;
 wire \rvcpu.dp.rf.reg_file_arr[14][19] ;
 wire \rvcpu.dp.rf.reg_file_arr[14][1] ;
 wire \rvcpu.dp.rf.reg_file_arr[14][20] ;
 wire \rvcpu.dp.rf.reg_file_arr[14][21] ;
 wire \rvcpu.dp.rf.reg_file_arr[14][22] ;
 wire \rvcpu.dp.rf.reg_file_arr[14][23] ;
 wire \rvcpu.dp.rf.reg_file_arr[14][24] ;
 wire \rvcpu.dp.rf.reg_file_arr[14][25] ;
 wire \rvcpu.dp.rf.reg_file_arr[14][26] ;
 wire \rvcpu.dp.rf.reg_file_arr[14][27] ;
 wire \rvcpu.dp.rf.reg_file_arr[14][28] ;
 wire \rvcpu.dp.rf.reg_file_arr[14][29] ;
 wire \rvcpu.dp.rf.reg_file_arr[14][2] ;
 wire \rvcpu.dp.rf.reg_file_arr[14][30] ;
 wire \rvcpu.dp.rf.reg_file_arr[14][31] ;
 wire \rvcpu.dp.rf.reg_file_arr[14][3] ;
 wire \rvcpu.dp.rf.reg_file_arr[14][4] ;
 wire \rvcpu.dp.rf.reg_file_arr[14][5] ;
 wire \rvcpu.dp.rf.reg_file_arr[14][6] ;
 wire \rvcpu.dp.rf.reg_file_arr[14][7] ;
 wire \rvcpu.dp.rf.reg_file_arr[14][8] ;
 wire \rvcpu.dp.rf.reg_file_arr[14][9] ;
 wire \rvcpu.dp.rf.reg_file_arr[15][0] ;
 wire \rvcpu.dp.rf.reg_file_arr[15][10] ;
 wire \rvcpu.dp.rf.reg_file_arr[15][11] ;
 wire \rvcpu.dp.rf.reg_file_arr[15][12] ;
 wire \rvcpu.dp.rf.reg_file_arr[15][13] ;
 wire \rvcpu.dp.rf.reg_file_arr[15][14] ;
 wire \rvcpu.dp.rf.reg_file_arr[15][15] ;
 wire \rvcpu.dp.rf.reg_file_arr[15][16] ;
 wire \rvcpu.dp.rf.reg_file_arr[15][17] ;
 wire \rvcpu.dp.rf.reg_file_arr[15][18] ;
 wire \rvcpu.dp.rf.reg_file_arr[15][19] ;
 wire \rvcpu.dp.rf.reg_file_arr[15][1] ;
 wire \rvcpu.dp.rf.reg_file_arr[15][20] ;
 wire \rvcpu.dp.rf.reg_file_arr[15][21] ;
 wire \rvcpu.dp.rf.reg_file_arr[15][22] ;
 wire \rvcpu.dp.rf.reg_file_arr[15][23] ;
 wire \rvcpu.dp.rf.reg_file_arr[15][24] ;
 wire \rvcpu.dp.rf.reg_file_arr[15][25] ;
 wire \rvcpu.dp.rf.reg_file_arr[15][26] ;
 wire \rvcpu.dp.rf.reg_file_arr[15][27] ;
 wire \rvcpu.dp.rf.reg_file_arr[15][28] ;
 wire \rvcpu.dp.rf.reg_file_arr[15][29] ;
 wire \rvcpu.dp.rf.reg_file_arr[15][2] ;
 wire \rvcpu.dp.rf.reg_file_arr[15][30] ;
 wire \rvcpu.dp.rf.reg_file_arr[15][31] ;
 wire \rvcpu.dp.rf.reg_file_arr[15][3] ;
 wire \rvcpu.dp.rf.reg_file_arr[15][4] ;
 wire \rvcpu.dp.rf.reg_file_arr[15][5] ;
 wire \rvcpu.dp.rf.reg_file_arr[15][6] ;
 wire \rvcpu.dp.rf.reg_file_arr[15][7] ;
 wire \rvcpu.dp.rf.reg_file_arr[15][8] ;
 wire \rvcpu.dp.rf.reg_file_arr[15][9] ;
 wire \rvcpu.dp.rf.reg_file_arr[16][0] ;
 wire \rvcpu.dp.rf.reg_file_arr[16][10] ;
 wire \rvcpu.dp.rf.reg_file_arr[16][11] ;
 wire \rvcpu.dp.rf.reg_file_arr[16][12] ;
 wire \rvcpu.dp.rf.reg_file_arr[16][13] ;
 wire \rvcpu.dp.rf.reg_file_arr[16][14] ;
 wire \rvcpu.dp.rf.reg_file_arr[16][15] ;
 wire \rvcpu.dp.rf.reg_file_arr[16][16] ;
 wire \rvcpu.dp.rf.reg_file_arr[16][17] ;
 wire \rvcpu.dp.rf.reg_file_arr[16][18] ;
 wire \rvcpu.dp.rf.reg_file_arr[16][19] ;
 wire \rvcpu.dp.rf.reg_file_arr[16][1] ;
 wire \rvcpu.dp.rf.reg_file_arr[16][20] ;
 wire \rvcpu.dp.rf.reg_file_arr[16][21] ;
 wire \rvcpu.dp.rf.reg_file_arr[16][22] ;
 wire \rvcpu.dp.rf.reg_file_arr[16][23] ;
 wire \rvcpu.dp.rf.reg_file_arr[16][24] ;
 wire \rvcpu.dp.rf.reg_file_arr[16][25] ;
 wire \rvcpu.dp.rf.reg_file_arr[16][26] ;
 wire \rvcpu.dp.rf.reg_file_arr[16][27] ;
 wire \rvcpu.dp.rf.reg_file_arr[16][28] ;
 wire \rvcpu.dp.rf.reg_file_arr[16][29] ;
 wire \rvcpu.dp.rf.reg_file_arr[16][2] ;
 wire \rvcpu.dp.rf.reg_file_arr[16][30] ;
 wire \rvcpu.dp.rf.reg_file_arr[16][31] ;
 wire \rvcpu.dp.rf.reg_file_arr[16][3] ;
 wire \rvcpu.dp.rf.reg_file_arr[16][4] ;
 wire \rvcpu.dp.rf.reg_file_arr[16][5] ;
 wire \rvcpu.dp.rf.reg_file_arr[16][6] ;
 wire \rvcpu.dp.rf.reg_file_arr[16][7] ;
 wire \rvcpu.dp.rf.reg_file_arr[16][8] ;
 wire \rvcpu.dp.rf.reg_file_arr[16][9] ;
 wire \rvcpu.dp.rf.reg_file_arr[17][0] ;
 wire \rvcpu.dp.rf.reg_file_arr[17][10] ;
 wire \rvcpu.dp.rf.reg_file_arr[17][11] ;
 wire \rvcpu.dp.rf.reg_file_arr[17][12] ;
 wire \rvcpu.dp.rf.reg_file_arr[17][13] ;
 wire \rvcpu.dp.rf.reg_file_arr[17][14] ;
 wire \rvcpu.dp.rf.reg_file_arr[17][15] ;
 wire \rvcpu.dp.rf.reg_file_arr[17][16] ;
 wire \rvcpu.dp.rf.reg_file_arr[17][17] ;
 wire \rvcpu.dp.rf.reg_file_arr[17][18] ;
 wire \rvcpu.dp.rf.reg_file_arr[17][19] ;
 wire \rvcpu.dp.rf.reg_file_arr[17][1] ;
 wire \rvcpu.dp.rf.reg_file_arr[17][20] ;
 wire \rvcpu.dp.rf.reg_file_arr[17][21] ;
 wire \rvcpu.dp.rf.reg_file_arr[17][22] ;
 wire \rvcpu.dp.rf.reg_file_arr[17][23] ;
 wire \rvcpu.dp.rf.reg_file_arr[17][24] ;
 wire \rvcpu.dp.rf.reg_file_arr[17][25] ;
 wire \rvcpu.dp.rf.reg_file_arr[17][26] ;
 wire \rvcpu.dp.rf.reg_file_arr[17][27] ;
 wire \rvcpu.dp.rf.reg_file_arr[17][28] ;
 wire \rvcpu.dp.rf.reg_file_arr[17][29] ;
 wire \rvcpu.dp.rf.reg_file_arr[17][2] ;
 wire \rvcpu.dp.rf.reg_file_arr[17][30] ;
 wire \rvcpu.dp.rf.reg_file_arr[17][31] ;
 wire \rvcpu.dp.rf.reg_file_arr[17][3] ;
 wire \rvcpu.dp.rf.reg_file_arr[17][4] ;
 wire \rvcpu.dp.rf.reg_file_arr[17][5] ;
 wire \rvcpu.dp.rf.reg_file_arr[17][6] ;
 wire \rvcpu.dp.rf.reg_file_arr[17][7] ;
 wire \rvcpu.dp.rf.reg_file_arr[17][8] ;
 wire \rvcpu.dp.rf.reg_file_arr[17][9] ;
 wire \rvcpu.dp.rf.reg_file_arr[18][0] ;
 wire \rvcpu.dp.rf.reg_file_arr[18][10] ;
 wire \rvcpu.dp.rf.reg_file_arr[18][11] ;
 wire \rvcpu.dp.rf.reg_file_arr[18][12] ;
 wire \rvcpu.dp.rf.reg_file_arr[18][13] ;
 wire \rvcpu.dp.rf.reg_file_arr[18][14] ;
 wire \rvcpu.dp.rf.reg_file_arr[18][15] ;
 wire \rvcpu.dp.rf.reg_file_arr[18][16] ;
 wire \rvcpu.dp.rf.reg_file_arr[18][17] ;
 wire \rvcpu.dp.rf.reg_file_arr[18][18] ;
 wire \rvcpu.dp.rf.reg_file_arr[18][19] ;
 wire \rvcpu.dp.rf.reg_file_arr[18][1] ;
 wire \rvcpu.dp.rf.reg_file_arr[18][20] ;
 wire \rvcpu.dp.rf.reg_file_arr[18][21] ;
 wire \rvcpu.dp.rf.reg_file_arr[18][22] ;
 wire \rvcpu.dp.rf.reg_file_arr[18][23] ;
 wire \rvcpu.dp.rf.reg_file_arr[18][24] ;
 wire \rvcpu.dp.rf.reg_file_arr[18][25] ;
 wire \rvcpu.dp.rf.reg_file_arr[18][26] ;
 wire \rvcpu.dp.rf.reg_file_arr[18][27] ;
 wire \rvcpu.dp.rf.reg_file_arr[18][28] ;
 wire \rvcpu.dp.rf.reg_file_arr[18][29] ;
 wire \rvcpu.dp.rf.reg_file_arr[18][2] ;
 wire \rvcpu.dp.rf.reg_file_arr[18][30] ;
 wire \rvcpu.dp.rf.reg_file_arr[18][31] ;
 wire \rvcpu.dp.rf.reg_file_arr[18][3] ;
 wire \rvcpu.dp.rf.reg_file_arr[18][4] ;
 wire \rvcpu.dp.rf.reg_file_arr[18][5] ;
 wire \rvcpu.dp.rf.reg_file_arr[18][6] ;
 wire \rvcpu.dp.rf.reg_file_arr[18][7] ;
 wire \rvcpu.dp.rf.reg_file_arr[18][8] ;
 wire \rvcpu.dp.rf.reg_file_arr[18][9] ;
 wire \rvcpu.dp.rf.reg_file_arr[19][0] ;
 wire \rvcpu.dp.rf.reg_file_arr[19][10] ;
 wire \rvcpu.dp.rf.reg_file_arr[19][11] ;
 wire \rvcpu.dp.rf.reg_file_arr[19][12] ;
 wire \rvcpu.dp.rf.reg_file_arr[19][13] ;
 wire \rvcpu.dp.rf.reg_file_arr[19][14] ;
 wire \rvcpu.dp.rf.reg_file_arr[19][15] ;
 wire \rvcpu.dp.rf.reg_file_arr[19][16] ;
 wire \rvcpu.dp.rf.reg_file_arr[19][17] ;
 wire \rvcpu.dp.rf.reg_file_arr[19][18] ;
 wire \rvcpu.dp.rf.reg_file_arr[19][19] ;
 wire \rvcpu.dp.rf.reg_file_arr[19][1] ;
 wire \rvcpu.dp.rf.reg_file_arr[19][20] ;
 wire \rvcpu.dp.rf.reg_file_arr[19][21] ;
 wire \rvcpu.dp.rf.reg_file_arr[19][22] ;
 wire \rvcpu.dp.rf.reg_file_arr[19][23] ;
 wire \rvcpu.dp.rf.reg_file_arr[19][24] ;
 wire \rvcpu.dp.rf.reg_file_arr[19][25] ;
 wire \rvcpu.dp.rf.reg_file_arr[19][26] ;
 wire \rvcpu.dp.rf.reg_file_arr[19][27] ;
 wire \rvcpu.dp.rf.reg_file_arr[19][28] ;
 wire \rvcpu.dp.rf.reg_file_arr[19][29] ;
 wire \rvcpu.dp.rf.reg_file_arr[19][2] ;
 wire \rvcpu.dp.rf.reg_file_arr[19][30] ;
 wire \rvcpu.dp.rf.reg_file_arr[19][31] ;
 wire \rvcpu.dp.rf.reg_file_arr[19][3] ;
 wire \rvcpu.dp.rf.reg_file_arr[19][4] ;
 wire \rvcpu.dp.rf.reg_file_arr[19][5] ;
 wire \rvcpu.dp.rf.reg_file_arr[19][6] ;
 wire \rvcpu.dp.rf.reg_file_arr[19][7] ;
 wire \rvcpu.dp.rf.reg_file_arr[19][8] ;
 wire \rvcpu.dp.rf.reg_file_arr[19][9] ;
 wire \rvcpu.dp.rf.reg_file_arr[1][0] ;
 wire \rvcpu.dp.rf.reg_file_arr[1][10] ;
 wire \rvcpu.dp.rf.reg_file_arr[1][11] ;
 wire \rvcpu.dp.rf.reg_file_arr[1][12] ;
 wire \rvcpu.dp.rf.reg_file_arr[1][13] ;
 wire \rvcpu.dp.rf.reg_file_arr[1][14] ;
 wire \rvcpu.dp.rf.reg_file_arr[1][15] ;
 wire \rvcpu.dp.rf.reg_file_arr[1][16] ;
 wire \rvcpu.dp.rf.reg_file_arr[1][17] ;
 wire \rvcpu.dp.rf.reg_file_arr[1][18] ;
 wire \rvcpu.dp.rf.reg_file_arr[1][19] ;
 wire \rvcpu.dp.rf.reg_file_arr[1][1] ;
 wire \rvcpu.dp.rf.reg_file_arr[1][20] ;
 wire \rvcpu.dp.rf.reg_file_arr[1][21] ;
 wire \rvcpu.dp.rf.reg_file_arr[1][22] ;
 wire \rvcpu.dp.rf.reg_file_arr[1][23] ;
 wire \rvcpu.dp.rf.reg_file_arr[1][24] ;
 wire \rvcpu.dp.rf.reg_file_arr[1][25] ;
 wire \rvcpu.dp.rf.reg_file_arr[1][26] ;
 wire \rvcpu.dp.rf.reg_file_arr[1][27] ;
 wire \rvcpu.dp.rf.reg_file_arr[1][28] ;
 wire \rvcpu.dp.rf.reg_file_arr[1][29] ;
 wire \rvcpu.dp.rf.reg_file_arr[1][2] ;
 wire \rvcpu.dp.rf.reg_file_arr[1][30] ;
 wire \rvcpu.dp.rf.reg_file_arr[1][31] ;
 wire \rvcpu.dp.rf.reg_file_arr[1][3] ;
 wire \rvcpu.dp.rf.reg_file_arr[1][4] ;
 wire \rvcpu.dp.rf.reg_file_arr[1][5] ;
 wire \rvcpu.dp.rf.reg_file_arr[1][6] ;
 wire \rvcpu.dp.rf.reg_file_arr[1][7] ;
 wire \rvcpu.dp.rf.reg_file_arr[1][8] ;
 wire \rvcpu.dp.rf.reg_file_arr[1][9] ;
 wire \rvcpu.dp.rf.reg_file_arr[20][0] ;
 wire \rvcpu.dp.rf.reg_file_arr[20][10] ;
 wire \rvcpu.dp.rf.reg_file_arr[20][11] ;
 wire \rvcpu.dp.rf.reg_file_arr[20][12] ;
 wire \rvcpu.dp.rf.reg_file_arr[20][13] ;
 wire \rvcpu.dp.rf.reg_file_arr[20][14] ;
 wire \rvcpu.dp.rf.reg_file_arr[20][15] ;
 wire \rvcpu.dp.rf.reg_file_arr[20][16] ;
 wire \rvcpu.dp.rf.reg_file_arr[20][17] ;
 wire \rvcpu.dp.rf.reg_file_arr[20][18] ;
 wire \rvcpu.dp.rf.reg_file_arr[20][19] ;
 wire \rvcpu.dp.rf.reg_file_arr[20][1] ;
 wire \rvcpu.dp.rf.reg_file_arr[20][20] ;
 wire \rvcpu.dp.rf.reg_file_arr[20][21] ;
 wire \rvcpu.dp.rf.reg_file_arr[20][22] ;
 wire \rvcpu.dp.rf.reg_file_arr[20][23] ;
 wire \rvcpu.dp.rf.reg_file_arr[20][24] ;
 wire \rvcpu.dp.rf.reg_file_arr[20][25] ;
 wire \rvcpu.dp.rf.reg_file_arr[20][26] ;
 wire \rvcpu.dp.rf.reg_file_arr[20][27] ;
 wire \rvcpu.dp.rf.reg_file_arr[20][28] ;
 wire \rvcpu.dp.rf.reg_file_arr[20][29] ;
 wire \rvcpu.dp.rf.reg_file_arr[20][2] ;
 wire \rvcpu.dp.rf.reg_file_arr[20][30] ;
 wire \rvcpu.dp.rf.reg_file_arr[20][31] ;
 wire \rvcpu.dp.rf.reg_file_arr[20][3] ;
 wire \rvcpu.dp.rf.reg_file_arr[20][4] ;
 wire \rvcpu.dp.rf.reg_file_arr[20][5] ;
 wire \rvcpu.dp.rf.reg_file_arr[20][6] ;
 wire \rvcpu.dp.rf.reg_file_arr[20][7] ;
 wire \rvcpu.dp.rf.reg_file_arr[20][8] ;
 wire \rvcpu.dp.rf.reg_file_arr[20][9] ;
 wire \rvcpu.dp.rf.reg_file_arr[21][0] ;
 wire \rvcpu.dp.rf.reg_file_arr[21][10] ;
 wire \rvcpu.dp.rf.reg_file_arr[21][11] ;
 wire \rvcpu.dp.rf.reg_file_arr[21][12] ;
 wire \rvcpu.dp.rf.reg_file_arr[21][13] ;
 wire \rvcpu.dp.rf.reg_file_arr[21][14] ;
 wire \rvcpu.dp.rf.reg_file_arr[21][15] ;
 wire \rvcpu.dp.rf.reg_file_arr[21][16] ;
 wire \rvcpu.dp.rf.reg_file_arr[21][17] ;
 wire \rvcpu.dp.rf.reg_file_arr[21][18] ;
 wire \rvcpu.dp.rf.reg_file_arr[21][19] ;
 wire \rvcpu.dp.rf.reg_file_arr[21][1] ;
 wire \rvcpu.dp.rf.reg_file_arr[21][20] ;
 wire \rvcpu.dp.rf.reg_file_arr[21][21] ;
 wire \rvcpu.dp.rf.reg_file_arr[21][22] ;
 wire \rvcpu.dp.rf.reg_file_arr[21][23] ;
 wire \rvcpu.dp.rf.reg_file_arr[21][24] ;
 wire \rvcpu.dp.rf.reg_file_arr[21][25] ;
 wire \rvcpu.dp.rf.reg_file_arr[21][26] ;
 wire \rvcpu.dp.rf.reg_file_arr[21][27] ;
 wire \rvcpu.dp.rf.reg_file_arr[21][28] ;
 wire \rvcpu.dp.rf.reg_file_arr[21][29] ;
 wire \rvcpu.dp.rf.reg_file_arr[21][2] ;
 wire \rvcpu.dp.rf.reg_file_arr[21][30] ;
 wire \rvcpu.dp.rf.reg_file_arr[21][31] ;
 wire \rvcpu.dp.rf.reg_file_arr[21][3] ;
 wire \rvcpu.dp.rf.reg_file_arr[21][4] ;
 wire \rvcpu.dp.rf.reg_file_arr[21][5] ;
 wire \rvcpu.dp.rf.reg_file_arr[21][6] ;
 wire \rvcpu.dp.rf.reg_file_arr[21][7] ;
 wire \rvcpu.dp.rf.reg_file_arr[21][8] ;
 wire \rvcpu.dp.rf.reg_file_arr[21][9] ;
 wire \rvcpu.dp.rf.reg_file_arr[22][0] ;
 wire \rvcpu.dp.rf.reg_file_arr[22][10] ;
 wire \rvcpu.dp.rf.reg_file_arr[22][11] ;
 wire \rvcpu.dp.rf.reg_file_arr[22][12] ;
 wire \rvcpu.dp.rf.reg_file_arr[22][13] ;
 wire \rvcpu.dp.rf.reg_file_arr[22][14] ;
 wire \rvcpu.dp.rf.reg_file_arr[22][15] ;
 wire \rvcpu.dp.rf.reg_file_arr[22][16] ;
 wire \rvcpu.dp.rf.reg_file_arr[22][17] ;
 wire \rvcpu.dp.rf.reg_file_arr[22][18] ;
 wire \rvcpu.dp.rf.reg_file_arr[22][19] ;
 wire \rvcpu.dp.rf.reg_file_arr[22][1] ;
 wire \rvcpu.dp.rf.reg_file_arr[22][20] ;
 wire \rvcpu.dp.rf.reg_file_arr[22][21] ;
 wire \rvcpu.dp.rf.reg_file_arr[22][22] ;
 wire \rvcpu.dp.rf.reg_file_arr[22][23] ;
 wire \rvcpu.dp.rf.reg_file_arr[22][24] ;
 wire \rvcpu.dp.rf.reg_file_arr[22][25] ;
 wire \rvcpu.dp.rf.reg_file_arr[22][26] ;
 wire \rvcpu.dp.rf.reg_file_arr[22][27] ;
 wire \rvcpu.dp.rf.reg_file_arr[22][28] ;
 wire \rvcpu.dp.rf.reg_file_arr[22][29] ;
 wire \rvcpu.dp.rf.reg_file_arr[22][2] ;
 wire \rvcpu.dp.rf.reg_file_arr[22][30] ;
 wire \rvcpu.dp.rf.reg_file_arr[22][31] ;
 wire \rvcpu.dp.rf.reg_file_arr[22][3] ;
 wire \rvcpu.dp.rf.reg_file_arr[22][4] ;
 wire \rvcpu.dp.rf.reg_file_arr[22][5] ;
 wire \rvcpu.dp.rf.reg_file_arr[22][6] ;
 wire \rvcpu.dp.rf.reg_file_arr[22][7] ;
 wire \rvcpu.dp.rf.reg_file_arr[22][8] ;
 wire \rvcpu.dp.rf.reg_file_arr[22][9] ;
 wire \rvcpu.dp.rf.reg_file_arr[23][0] ;
 wire \rvcpu.dp.rf.reg_file_arr[23][10] ;
 wire \rvcpu.dp.rf.reg_file_arr[23][11] ;
 wire \rvcpu.dp.rf.reg_file_arr[23][12] ;
 wire \rvcpu.dp.rf.reg_file_arr[23][13] ;
 wire \rvcpu.dp.rf.reg_file_arr[23][14] ;
 wire \rvcpu.dp.rf.reg_file_arr[23][15] ;
 wire \rvcpu.dp.rf.reg_file_arr[23][16] ;
 wire \rvcpu.dp.rf.reg_file_arr[23][17] ;
 wire \rvcpu.dp.rf.reg_file_arr[23][18] ;
 wire \rvcpu.dp.rf.reg_file_arr[23][19] ;
 wire \rvcpu.dp.rf.reg_file_arr[23][1] ;
 wire \rvcpu.dp.rf.reg_file_arr[23][20] ;
 wire \rvcpu.dp.rf.reg_file_arr[23][21] ;
 wire \rvcpu.dp.rf.reg_file_arr[23][22] ;
 wire \rvcpu.dp.rf.reg_file_arr[23][23] ;
 wire \rvcpu.dp.rf.reg_file_arr[23][24] ;
 wire \rvcpu.dp.rf.reg_file_arr[23][25] ;
 wire \rvcpu.dp.rf.reg_file_arr[23][26] ;
 wire \rvcpu.dp.rf.reg_file_arr[23][27] ;
 wire \rvcpu.dp.rf.reg_file_arr[23][28] ;
 wire \rvcpu.dp.rf.reg_file_arr[23][29] ;
 wire \rvcpu.dp.rf.reg_file_arr[23][2] ;
 wire \rvcpu.dp.rf.reg_file_arr[23][30] ;
 wire \rvcpu.dp.rf.reg_file_arr[23][31] ;
 wire \rvcpu.dp.rf.reg_file_arr[23][3] ;
 wire \rvcpu.dp.rf.reg_file_arr[23][4] ;
 wire \rvcpu.dp.rf.reg_file_arr[23][5] ;
 wire \rvcpu.dp.rf.reg_file_arr[23][6] ;
 wire \rvcpu.dp.rf.reg_file_arr[23][7] ;
 wire \rvcpu.dp.rf.reg_file_arr[23][8] ;
 wire \rvcpu.dp.rf.reg_file_arr[23][9] ;
 wire \rvcpu.dp.rf.reg_file_arr[24][0] ;
 wire \rvcpu.dp.rf.reg_file_arr[24][10] ;
 wire \rvcpu.dp.rf.reg_file_arr[24][11] ;
 wire \rvcpu.dp.rf.reg_file_arr[24][12] ;
 wire \rvcpu.dp.rf.reg_file_arr[24][13] ;
 wire \rvcpu.dp.rf.reg_file_arr[24][14] ;
 wire \rvcpu.dp.rf.reg_file_arr[24][15] ;
 wire \rvcpu.dp.rf.reg_file_arr[24][16] ;
 wire \rvcpu.dp.rf.reg_file_arr[24][17] ;
 wire \rvcpu.dp.rf.reg_file_arr[24][18] ;
 wire \rvcpu.dp.rf.reg_file_arr[24][19] ;
 wire \rvcpu.dp.rf.reg_file_arr[24][1] ;
 wire \rvcpu.dp.rf.reg_file_arr[24][20] ;
 wire \rvcpu.dp.rf.reg_file_arr[24][21] ;
 wire \rvcpu.dp.rf.reg_file_arr[24][22] ;
 wire \rvcpu.dp.rf.reg_file_arr[24][23] ;
 wire \rvcpu.dp.rf.reg_file_arr[24][24] ;
 wire \rvcpu.dp.rf.reg_file_arr[24][25] ;
 wire \rvcpu.dp.rf.reg_file_arr[24][26] ;
 wire \rvcpu.dp.rf.reg_file_arr[24][27] ;
 wire \rvcpu.dp.rf.reg_file_arr[24][28] ;
 wire \rvcpu.dp.rf.reg_file_arr[24][29] ;
 wire \rvcpu.dp.rf.reg_file_arr[24][2] ;
 wire \rvcpu.dp.rf.reg_file_arr[24][30] ;
 wire \rvcpu.dp.rf.reg_file_arr[24][31] ;
 wire \rvcpu.dp.rf.reg_file_arr[24][3] ;
 wire \rvcpu.dp.rf.reg_file_arr[24][4] ;
 wire \rvcpu.dp.rf.reg_file_arr[24][5] ;
 wire \rvcpu.dp.rf.reg_file_arr[24][6] ;
 wire \rvcpu.dp.rf.reg_file_arr[24][7] ;
 wire \rvcpu.dp.rf.reg_file_arr[24][8] ;
 wire \rvcpu.dp.rf.reg_file_arr[24][9] ;
 wire \rvcpu.dp.rf.reg_file_arr[25][0] ;
 wire \rvcpu.dp.rf.reg_file_arr[25][10] ;
 wire \rvcpu.dp.rf.reg_file_arr[25][11] ;
 wire \rvcpu.dp.rf.reg_file_arr[25][12] ;
 wire \rvcpu.dp.rf.reg_file_arr[25][13] ;
 wire \rvcpu.dp.rf.reg_file_arr[25][14] ;
 wire \rvcpu.dp.rf.reg_file_arr[25][15] ;
 wire \rvcpu.dp.rf.reg_file_arr[25][16] ;
 wire \rvcpu.dp.rf.reg_file_arr[25][17] ;
 wire \rvcpu.dp.rf.reg_file_arr[25][18] ;
 wire \rvcpu.dp.rf.reg_file_arr[25][19] ;
 wire \rvcpu.dp.rf.reg_file_arr[25][1] ;
 wire \rvcpu.dp.rf.reg_file_arr[25][20] ;
 wire \rvcpu.dp.rf.reg_file_arr[25][21] ;
 wire \rvcpu.dp.rf.reg_file_arr[25][22] ;
 wire \rvcpu.dp.rf.reg_file_arr[25][23] ;
 wire \rvcpu.dp.rf.reg_file_arr[25][24] ;
 wire \rvcpu.dp.rf.reg_file_arr[25][25] ;
 wire \rvcpu.dp.rf.reg_file_arr[25][26] ;
 wire \rvcpu.dp.rf.reg_file_arr[25][27] ;
 wire \rvcpu.dp.rf.reg_file_arr[25][28] ;
 wire \rvcpu.dp.rf.reg_file_arr[25][29] ;
 wire \rvcpu.dp.rf.reg_file_arr[25][2] ;
 wire \rvcpu.dp.rf.reg_file_arr[25][30] ;
 wire \rvcpu.dp.rf.reg_file_arr[25][31] ;
 wire \rvcpu.dp.rf.reg_file_arr[25][3] ;
 wire \rvcpu.dp.rf.reg_file_arr[25][4] ;
 wire \rvcpu.dp.rf.reg_file_arr[25][5] ;
 wire \rvcpu.dp.rf.reg_file_arr[25][6] ;
 wire \rvcpu.dp.rf.reg_file_arr[25][7] ;
 wire \rvcpu.dp.rf.reg_file_arr[25][8] ;
 wire \rvcpu.dp.rf.reg_file_arr[25][9] ;
 wire \rvcpu.dp.rf.reg_file_arr[26][0] ;
 wire \rvcpu.dp.rf.reg_file_arr[26][10] ;
 wire \rvcpu.dp.rf.reg_file_arr[26][11] ;
 wire \rvcpu.dp.rf.reg_file_arr[26][12] ;
 wire \rvcpu.dp.rf.reg_file_arr[26][13] ;
 wire \rvcpu.dp.rf.reg_file_arr[26][14] ;
 wire \rvcpu.dp.rf.reg_file_arr[26][15] ;
 wire \rvcpu.dp.rf.reg_file_arr[26][16] ;
 wire \rvcpu.dp.rf.reg_file_arr[26][17] ;
 wire \rvcpu.dp.rf.reg_file_arr[26][18] ;
 wire \rvcpu.dp.rf.reg_file_arr[26][19] ;
 wire \rvcpu.dp.rf.reg_file_arr[26][1] ;
 wire \rvcpu.dp.rf.reg_file_arr[26][20] ;
 wire \rvcpu.dp.rf.reg_file_arr[26][21] ;
 wire \rvcpu.dp.rf.reg_file_arr[26][22] ;
 wire \rvcpu.dp.rf.reg_file_arr[26][23] ;
 wire \rvcpu.dp.rf.reg_file_arr[26][24] ;
 wire \rvcpu.dp.rf.reg_file_arr[26][25] ;
 wire \rvcpu.dp.rf.reg_file_arr[26][26] ;
 wire \rvcpu.dp.rf.reg_file_arr[26][27] ;
 wire \rvcpu.dp.rf.reg_file_arr[26][28] ;
 wire \rvcpu.dp.rf.reg_file_arr[26][29] ;
 wire \rvcpu.dp.rf.reg_file_arr[26][2] ;
 wire \rvcpu.dp.rf.reg_file_arr[26][30] ;
 wire \rvcpu.dp.rf.reg_file_arr[26][31] ;
 wire \rvcpu.dp.rf.reg_file_arr[26][3] ;
 wire \rvcpu.dp.rf.reg_file_arr[26][4] ;
 wire \rvcpu.dp.rf.reg_file_arr[26][5] ;
 wire \rvcpu.dp.rf.reg_file_arr[26][6] ;
 wire \rvcpu.dp.rf.reg_file_arr[26][7] ;
 wire \rvcpu.dp.rf.reg_file_arr[26][8] ;
 wire \rvcpu.dp.rf.reg_file_arr[26][9] ;
 wire \rvcpu.dp.rf.reg_file_arr[27][0] ;
 wire \rvcpu.dp.rf.reg_file_arr[27][10] ;
 wire \rvcpu.dp.rf.reg_file_arr[27][11] ;
 wire \rvcpu.dp.rf.reg_file_arr[27][12] ;
 wire \rvcpu.dp.rf.reg_file_arr[27][13] ;
 wire \rvcpu.dp.rf.reg_file_arr[27][14] ;
 wire \rvcpu.dp.rf.reg_file_arr[27][15] ;
 wire \rvcpu.dp.rf.reg_file_arr[27][16] ;
 wire \rvcpu.dp.rf.reg_file_arr[27][17] ;
 wire \rvcpu.dp.rf.reg_file_arr[27][18] ;
 wire \rvcpu.dp.rf.reg_file_arr[27][19] ;
 wire \rvcpu.dp.rf.reg_file_arr[27][1] ;
 wire \rvcpu.dp.rf.reg_file_arr[27][20] ;
 wire \rvcpu.dp.rf.reg_file_arr[27][21] ;
 wire \rvcpu.dp.rf.reg_file_arr[27][22] ;
 wire \rvcpu.dp.rf.reg_file_arr[27][23] ;
 wire \rvcpu.dp.rf.reg_file_arr[27][24] ;
 wire \rvcpu.dp.rf.reg_file_arr[27][25] ;
 wire \rvcpu.dp.rf.reg_file_arr[27][26] ;
 wire \rvcpu.dp.rf.reg_file_arr[27][27] ;
 wire \rvcpu.dp.rf.reg_file_arr[27][28] ;
 wire \rvcpu.dp.rf.reg_file_arr[27][29] ;
 wire \rvcpu.dp.rf.reg_file_arr[27][2] ;
 wire \rvcpu.dp.rf.reg_file_arr[27][30] ;
 wire \rvcpu.dp.rf.reg_file_arr[27][31] ;
 wire \rvcpu.dp.rf.reg_file_arr[27][3] ;
 wire \rvcpu.dp.rf.reg_file_arr[27][4] ;
 wire \rvcpu.dp.rf.reg_file_arr[27][5] ;
 wire \rvcpu.dp.rf.reg_file_arr[27][6] ;
 wire \rvcpu.dp.rf.reg_file_arr[27][7] ;
 wire \rvcpu.dp.rf.reg_file_arr[27][8] ;
 wire \rvcpu.dp.rf.reg_file_arr[27][9] ;
 wire \rvcpu.dp.rf.reg_file_arr[28][0] ;
 wire \rvcpu.dp.rf.reg_file_arr[28][10] ;
 wire \rvcpu.dp.rf.reg_file_arr[28][11] ;
 wire \rvcpu.dp.rf.reg_file_arr[28][12] ;
 wire \rvcpu.dp.rf.reg_file_arr[28][13] ;
 wire \rvcpu.dp.rf.reg_file_arr[28][14] ;
 wire \rvcpu.dp.rf.reg_file_arr[28][15] ;
 wire \rvcpu.dp.rf.reg_file_arr[28][16] ;
 wire \rvcpu.dp.rf.reg_file_arr[28][17] ;
 wire \rvcpu.dp.rf.reg_file_arr[28][18] ;
 wire \rvcpu.dp.rf.reg_file_arr[28][19] ;
 wire \rvcpu.dp.rf.reg_file_arr[28][1] ;
 wire \rvcpu.dp.rf.reg_file_arr[28][20] ;
 wire \rvcpu.dp.rf.reg_file_arr[28][21] ;
 wire \rvcpu.dp.rf.reg_file_arr[28][22] ;
 wire \rvcpu.dp.rf.reg_file_arr[28][23] ;
 wire \rvcpu.dp.rf.reg_file_arr[28][24] ;
 wire \rvcpu.dp.rf.reg_file_arr[28][25] ;
 wire \rvcpu.dp.rf.reg_file_arr[28][26] ;
 wire \rvcpu.dp.rf.reg_file_arr[28][27] ;
 wire \rvcpu.dp.rf.reg_file_arr[28][28] ;
 wire \rvcpu.dp.rf.reg_file_arr[28][29] ;
 wire \rvcpu.dp.rf.reg_file_arr[28][2] ;
 wire \rvcpu.dp.rf.reg_file_arr[28][30] ;
 wire \rvcpu.dp.rf.reg_file_arr[28][31] ;
 wire \rvcpu.dp.rf.reg_file_arr[28][3] ;
 wire \rvcpu.dp.rf.reg_file_arr[28][4] ;
 wire \rvcpu.dp.rf.reg_file_arr[28][5] ;
 wire \rvcpu.dp.rf.reg_file_arr[28][6] ;
 wire \rvcpu.dp.rf.reg_file_arr[28][7] ;
 wire \rvcpu.dp.rf.reg_file_arr[28][8] ;
 wire \rvcpu.dp.rf.reg_file_arr[28][9] ;
 wire \rvcpu.dp.rf.reg_file_arr[29][0] ;
 wire \rvcpu.dp.rf.reg_file_arr[29][10] ;
 wire \rvcpu.dp.rf.reg_file_arr[29][11] ;
 wire \rvcpu.dp.rf.reg_file_arr[29][12] ;
 wire \rvcpu.dp.rf.reg_file_arr[29][13] ;
 wire \rvcpu.dp.rf.reg_file_arr[29][14] ;
 wire \rvcpu.dp.rf.reg_file_arr[29][15] ;
 wire \rvcpu.dp.rf.reg_file_arr[29][16] ;
 wire \rvcpu.dp.rf.reg_file_arr[29][17] ;
 wire \rvcpu.dp.rf.reg_file_arr[29][18] ;
 wire \rvcpu.dp.rf.reg_file_arr[29][19] ;
 wire \rvcpu.dp.rf.reg_file_arr[29][1] ;
 wire \rvcpu.dp.rf.reg_file_arr[29][20] ;
 wire \rvcpu.dp.rf.reg_file_arr[29][21] ;
 wire \rvcpu.dp.rf.reg_file_arr[29][22] ;
 wire \rvcpu.dp.rf.reg_file_arr[29][23] ;
 wire \rvcpu.dp.rf.reg_file_arr[29][24] ;
 wire \rvcpu.dp.rf.reg_file_arr[29][25] ;
 wire \rvcpu.dp.rf.reg_file_arr[29][26] ;
 wire \rvcpu.dp.rf.reg_file_arr[29][27] ;
 wire \rvcpu.dp.rf.reg_file_arr[29][28] ;
 wire \rvcpu.dp.rf.reg_file_arr[29][29] ;
 wire \rvcpu.dp.rf.reg_file_arr[29][2] ;
 wire \rvcpu.dp.rf.reg_file_arr[29][30] ;
 wire \rvcpu.dp.rf.reg_file_arr[29][31] ;
 wire \rvcpu.dp.rf.reg_file_arr[29][3] ;
 wire \rvcpu.dp.rf.reg_file_arr[29][4] ;
 wire \rvcpu.dp.rf.reg_file_arr[29][5] ;
 wire \rvcpu.dp.rf.reg_file_arr[29][6] ;
 wire \rvcpu.dp.rf.reg_file_arr[29][7] ;
 wire \rvcpu.dp.rf.reg_file_arr[29][8] ;
 wire \rvcpu.dp.rf.reg_file_arr[29][9] ;
 wire \rvcpu.dp.rf.reg_file_arr[2][0] ;
 wire \rvcpu.dp.rf.reg_file_arr[2][10] ;
 wire \rvcpu.dp.rf.reg_file_arr[2][11] ;
 wire \rvcpu.dp.rf.reg_file_arr[2][12] ;
 wire \rvcpu.dp.rf.reg_file_arr[2][13] ;
 wire \rvcpu.dp.rf.reg_file_arr[2][14] ;
 wire \rvcpu.dp.rf.reg_file_arr[2][15] ;
 wire \rvcpu.dp.rf.reg_file_arr[2][16] ;
 wire \rvcpu.dp.rf.reg_file_arr[2][17] ;
 wire \rvcpu.dp.rf.reg_file_arr[2][18] ;
 wire \rvcpu.dp.rf.reg_file_arr[2][19] ;
 wire \rvcpu.dp.rf.reg_file_arr[2][1] ;
 wire \rvcpu.dp.rf.reg_file_arr[2][20] ;
 wire \rvcpu.dp.rf.reg_file_arr[2][21] ;
 wire \rvcpu.dp.rf.reg_file_arr[2][22] ;
 wire \rvcpu.dp.rf.reg_file_arr[2][23] ;
 wire \rvcpu.dp.rf.reg_file_arr[2][24] ;
 wire \rvcpu.dp.rf.reg_file_arr[2][25] ;
 wire \rvcpu.dp.rf.reg_file_arr[2][26] ;
 wire \rvcpu.dp.rf.reg_file_arr[2][27] ;
 wire \rvcpu.dp.rf.reg_file_arr[2][28] ;
 wire \rvcpu.dp.rf.reg_file_arr[2][29] ;
 wire \rvcpu.dp.rf.reg_file_arr[2][2] ;
 wire \rvcpu.dp.rf.reg_file_arr[2][30] ;
 wire \rvcpu.dp.rf.reg_file_arr[2][31] ;
 wire \rvcpu.dp.rf.reg_file_arr[2][3] ;
 wire \rvcpu.dp.rf.reg_file_arr[2][4] ;
 wire \rvcpu.dp.rf.reg_file_arr[2][5] ;
 wire \rvcpu.dp.rf.reg_file_arr[2][6] ;
 wire \rvcpu.dp.rf.reg_file_arr[2][7] ;
 wire \rvcpu.dp.rf.reg_file_arr[2][8] ;
 wire \rvcpu.dp.rf.reg_file_arr[2][9] ;
 wire \rvcpu.dp.rf.reg_file_arr[30][0] ;
 wire \rvcpu.dp.rf.reg_file_arr[30][10] ;
 wire \rvcpu.dp.rf.reg_file_arr[30][11] ;
 wire \rvcpu.dp.rf.reg_file_arr[30][12] ;
 wire \rvcpu.dp.rf.reg_file_arr[30][13] ;
 wire \rvcpu.dp.rf.reg_file_arr[30][14] ;
 wire \rvcpu.dp.rf.reg_file_arr[30][15] ;
 wire \rvcpu.dp.rf.reg_file_arr[30][16] ;
 wire \rvcpu.dp.rf.reg_file_arr[30][17] ;
 wire \rvcpu.dp.rf.reg_file_arr[30][18] ;
 wire \rvcpu.dp.rf.reg_file_arr[30][19] ;
 wire \rvcpu.dp.rf.reg_file_arr[30][1] ;
 wire \rvcpu.dp.rf.reg_file_arr[30][20] ;
 wire \rvcpu.dp.rf.reg_file_arr[30][21] ;
 wire \rvcpu.dp.rf.reg_file_arr[30][22] ;
 wire \rvcpu.dp.rf.reg_file_arr[30][23] ;
 wire \rvcpu.dp.rf.reg_file_arr[30][24] ;
 wire \rvcpu.dp.rf.reg_file_arr[30][25] ;
 wire \rvcpu.dp.rf.reg_file_arr[30][26] ;
 wire \rvcpu.dp.rf.reg_file_arr[30][27] ;
 wire \rvcpu.dp.rf.reg_file_arr[30][28] ;
 wire \rvcpu.dp.rf.reg_file_arr[30][29] ;
 wire \rvcpu.dp.rf.reg_file_arr[30][2] ;
 wire \rvcpu.dp.rf.reg_file_arr[30][30] ;
 wire \rvcpu.dp.rf.reg_file_arr[30][31] ;
 wire \rvcpu.dp.rf.reg_file_arr[30][3] ;
 wire \rvcpu.dp.rf.reg_file_arr[30][4] ;
 wire \rvcpu.dp.rf.reg_file_arr[30][5] ;
 wire \rvcpu.dp.rf.reg_file_arr[30][6] ;
 wire \rvcpu.dp.rf.reg_file_arr[30][7] ;
 wire \rvcpu.dp.rf.reg_file_arr[30][8] ;
 wire \rvcpu.dp.rf.reg_file_arr[30][9] ;
 wire \rvcpu.dp.rf.reg_file_arr[31][0] ;
 wire \rvcpu.dp.rf.reg_file_arr[31][10] ;
 wire \rvcpu.dp.rf.reg_file_arr[31][11] ;
 wire \rvcpu.dp.rf.reg_file_arr[31][12] ;
 wire \rvcpu.dp.rf.reg_file_arr[31][13] ;
 wire \rvcpu.dp.rf.reg_file_arr[31][14] ;
 wire \rvcpu.dp.rf.reg_file_arr[31][15] ;
 wire \rvcpu.dp.rf.reg_file_arr[31][16] ;
 wire \rvcpu.dp.rf.reg_file_arr[31][17] ;
 wire \rvcpu.dp.rf.reg_file_arr[31][18] ;
 wire \rvcpu.dp.rf.reg_file_arr[31][19] ;
 wire \rvcpu.dp.rf.reg_file_arr[31][1] ;
 wire \rvcpu.dp.rf.reg_file_arr[31][20] ;
 wire \rvcpu.dp.rf.reg_file_arr[31][21] ;
 wire \rvcpu.dp.rf.reg_file_arr[31][22] ;
 wire \rvcpu.dp.rf.reg_file_arr[31][23] ;
 wire \rvcpu.dp.rf.reg_file_arr[31][24] ;
 wire \rvcpu.dp.rf.reg_file_arr[31][25] ;
 wire \rvcpu.dp.rf.reg_file_arr[31][26] ;
 wire \rvcpu.dp.rf.reg_file_arr[31][27] ;
 wire \rvcpu.dp.rf.reg_file_arr[31][28] ;
 wire \rvcpu.dp.rf.reg_file_arr[31][29] ;
 wire \rvcpu.dp.rf.reg_file_arr[31][2] ;
 wire \rvcpu.dp.rf.reg_file_arr[31][30] ;
 wire \rvcpu.dp.rf.reg_file_arr[31][31] ;
 wire \rvcpu.dp.rf.reg_file_arr[31][3] ;
 wire \rvcpu.dp.rf.reg_file_arr[31][4] ;
 wire \rvcpu.dp.rf.reg_file_arr[31][5] ;
 wire \rvcpu.dp.rf.reg_file_arr[31][6] ;
 wire \rvcpu.dp.rf.reg_file_arr[31][7] ;
 wire \rvcpu.dp.rf.reg_file_arr[31][8] ;
 wire \rvcpu.dp.rf.reg_file_arr[31][9] ;
 wire \rvcpu.dp.rf.reg_file_arr[3][0] ;
 wire \rvcpu.dp.rf.reg_file_arr[3][10] ;
 wire \rvcpu.dp.rf.reg_file_arr[3][11] ;
 wire \rvcpu.dp.rf.reg_file_arr[3][12] ;
 wire \rvcpu.dp.rf.reg_file_arr[3][13] ;
 wire \rvcpu.dp.rf.reg_file_arr[3][14] ;
 wire \rvcpu.dp.rf.reg_file_arr[3][15] ;
 wire \rvcpu.dp.rf.reg_file_arr[3][16] ;
 wire \rvcpu.dp.rf.reg_file_arr[3][17] ;
 wire \rvcpu.dp.rf.reg_file_arr[3][18] ;
 wire \rvcpu.dp.rf.reg_file_arr[3][19] ;
 wire \rvcpu.dp.rf.reg_file_arr[3][1] ;
 wire \rvcpu.dp.rf.reg_file_arr[3][20] ;
 wire \rvcpu.dp.rf.reg_file_arr[3][21] ;
 wire \rvcpu.dp.rf.reg_file_arr[3][22] ;
 wire \rvcpu.dp.rf.reg_file_arr[3][23] ;
 wire \rvcpu.dp.rf.reg_file_arr[3][24] ;
 wire \rvcpu.dp.rf.reg_file_arr[3][25] ;
 wire \rvcpu.dp.rf.reg_file_arr[3][26] ;
 wire \rvcpu.dp.rf.reg_file_arr[3][27] ;
 wire \rvcpu.dp.rf.reg_file_arr[3][28] ;
 wire \rvcpu.dp.rf.reg_file_arr[3][29] ;
 wire \rvcpu.dp.rf.reg_file_arr[3][2] ;
 wire \rvcpu.dp.rf.reg_file_arr[3][30] ;
 wire \rvcpu.dp.rf.reg_file_arr[3][31] ;
 wire \rvcpu.dp.rf.reg_file_arr[3][3] ;
 wire \rvcpu.dp.rf.reg_file_arr[3][4] ;
 wire \rvcpu.dp.rf.reg_file_arr[3][5] ;
 wire \rvcpu.dp.rf.reg_file_arr[3][6] ;
 wire \rvcpu.dp.rf.reg_file_arr[3][7] ;
 wire \rvcpu.dp.rf.reg_file_arr[3][8] ;
 wire \rvcpu.dp.rf.reg_file_arr[3][9] ;
 wire \rvcpu.dp.rf.reg_file_arr[4][0] ;
 wire \rvcpu.dp.rf.reg_file_arr[4][10] ;
 wire \rvcpu.dp.rf.reg_file_arr[4][11] ;
 wire \rvcpu.dp.rf.reg_file_arr[4][12] ;
 wire \rvcpu.dp.rf.reg_file_arr[4][13] ;
 wire \rvcpu.dp.rf.reg_file_arr[4][14] ;
 wire \rvcpu.dp.rf.reg_file_arr[4][15] ;
 wire \rvcpu.dp.rf.reg_file_arr[4][16] ;
 wire \rvcpu.dp.rf.reg_file_arr[4][17] ;
 wire \rvcpu.dp.rf.reg_file_arr[4][18] ;
 wire \rvcpu.dp.rf.reg_file_arr[4][19] ;
 wire \rvcpu.dp.rf.reg_file_arr[4][1] ;
 wire \rvcpu.dp.rf.reg_file_arr[4][20] ;
 wire \rvcpu.dp.rf.reg_file_arr[4][21] ;
 wire \rvcpu.dp.rf.reg_file_arr[4][22] ;
 wire \rvcpu.dp.rf.reg_file_arr[4][23] ;
 wire \rvcpu.dp.rf.reg_file_arr[4][24] ;
 wire \rvcpu.dp.rf.reg_file_arr[4][25] ;
 wire \rvcpu.dp.rf.reg_file_arr[4][26] ;
 wire \rvcpu.dp.rf.reg_file_arr[4][27] ;
 wire \rvcpu.dp.rf.reg_file_arr[4][28] ;
 wire \rvcpu.dp.rf.reg_file_arr[4][29] ;
 wire \rvcpu.dp.rf.reg_file_arr[4][2] ;
 wire \rvcpu.dp.rf.reg_file_arr[4][30] ;
 wire \rvcpu.dp.rf.reg_file_arr[4][31] ;
 wire \rvcpu.dp.rf.reg_file_arr[4][3] ;
 wire \rvcpu.dp.rf.reg_file_arr[4][4] ;
 wire \rvcpu.dp.rf.reg_file_arr[4][5] ;
 wire \rvcpu.dp.rf.reg_file_arr[4][6] ;
 wire \rvcpu.dp.rf.reg_file_arr[4][7] ;
 wire \rvcpu.dp.rf.reg_file_arr[4][8] ;
 wire \rvcpu.dp.rf.reg_file_arr[4][9] ;
 wire \rvcpu.dp.rf.reg_file_arr[5][0] ;
 wire \rvcpu.dp.rf.reg_file_arr[5][10] ;
 wire \rvcpu.dp.rf.reg_file_arr[5][11] ;
 wire \rvcpu.dp.rf.reg_file_arr[5][12] ;
 wire \rvcpu.dp.rf.reg_file_arr[5][13] ;
 wire \rvcpu.dp.rf.reg_file_arr[5][14] ;
 wire \rvcpu.dp.rf.reg_file_arr[5][15] ;
 wire \rvcpu.dp.rf.reg_file_arr[5][16] ;
 wire \rvcpu.dp.rf.reg_file_arr[5][17] ;
 wire \rvcpu.dp.rf.reg_file_arr[5][18] ;
 wire \rvcpu.dp.rf.reg_file_arr[5][19] ;
 wire \rvcpu.dp.rf.reg_file_arr[5][1] ;
 wire \rvcpu.dp.rf.reg_file_arr[5][20] ;
 wire \rvcpu.dp.rf.reg_file_arr[5][21] ;
 wire \rvcpu.dp.rf.reg_file_arr[5][22] ;
 wire \rvcpu.dp.rf.reg_file_arr[5][23] ;
 wire \rvcpu.dp.rf.reg_file_arr[5][24] ;
 wire \rvcpu.dp.rf.reg_file_arr[5][25] ;
 wire \rvcpu.dp.rf.reg_file_arr[5][26] ;
 wire \rvcpu.dp.rf.reg_file_arr[5][27] ;
 wire \rvcpu.dp.rf.reg_file_arr[5][28] ;
 wire \rvcpu.dp.rf.reg_file_arr[5][29] ;
 wire \rvcpu.dp.rf.reg_file_arr[5][2] ;
 wire \rvcpu.dp.rf.reg_file_arr[5][30] ;
 wire \rvcpu.dp.rf.reg_file_arr[5][31] ;
 wire \rvcpu.dp.rf.reg_file_arr[5][3] ;
 wire \rvcpu.dp.rf.reg_file_arr[5][4] ;
 wire \rvcpu.dp.rf.reg_file_arr[5][5] ;
 wire \rvcpu.dp.rf.reg_file_arr[5][6] ;
 wire \rvcpu.dp.rf.reg_file_arr[5][7] ;
 wire \rvcpu.dp.rf.reg_file_arr[5][8] ;
 wire \rvcpu.dp.rf.reg_file_arr[5][9] ;
 wire \rvcpu.dp.rf.reg_file_arr[6][0] ;
 wire \rvcpu.dp.rf.reg_file_arr[6][10] ;
 wire \rvcpu.dp.rf.reg_file_arr[6][11] ;
 wire \rvcpu.dp.rf.reg_file_arr[6][12] ;
 wire \rvcpu.dp.rf.reg_file_arr[6][13] ;
 wire \rvcpu.dp.rf.reg_file_arr[6][14] ;
 wire \rvcpu.dp.rf.reg_file_arr[6][15] ;
 wire \rvcpu.dp.rf.reg_file_arr[6][16] ;
 wire \rvcpu.dp.rf.reg_file_arr[6][17] ;
 wire \rvcpu.dp.rf.reg_file_arr[6][18] ;
 wire \rvcpu.dp.rf.reg_file_arr[6][19] ;
 wire \rvcpu.dp.rf.reg_file_arr[6][1] ;
 wire \rvcpu.dp.rf.reg_file_arr[6][20] ;
 wire \rvcpu.dp.rf.reg_file_arr[6][21] ;
 wire \rvcpu.dp.rf.reg_file_arr[6][22] ;
 wire \rvcpu.dp.rf.reg_file_arr[6][23] ;
 wire \rvcpu.dp.rf.reg_file_arr[6][24] ;
 wire \rvcpu.dp.rf.reg_file_arr[6][25] ;
 wire \rvcpu.dp.rf.reg_file_arr[6][26] ;
 wire \rvcpu.dp.rf.reg_file_arr[6][27] ;
 wire \rvcpu.dp.rf.reg_file_arr[6][28] ;
 wire \rvcpu.dp.rf.reg_file_arr[6][29] ;
 wire \rvcpu.dp.rf.reg_file_arr[6][2] ;
 wire \rvcpu.dp.rf.reg_file_arr[6][30] ;
 wire \rvcpu.dp.rf.reg_file_arr[6][31] ;
 wire \rvcpu.dp.rf.reg_file_arr[6][3] ;
 wire \rvcpu.dp.rf.reg_file_arr[6][4] ;
 wire \rvcpu.dp.rf.reg_file_arr[6][5] ;
 wire \rvcpu.dp.rf.reg_file_arr[6][6] ;
 wire \rvcpu.dp.rf.reg_file_arr[6][7] ;
 wire \rvcpu.dp.rf.reg_file_arr[6][8] ;
 wire \rvcpu.dp.rf.reg_file_arr[6][9] ;
 wire \rvcpu.dp.rf.reg_file_arr[7][0] ;
 wire \rvcpu.dp.rf.reg_file_arr[7][10] ;
 wire \rvcpu.dp.rf.reg_file_arr[7][11] ;
 wire \rvcpu.dp.rf.reg_file_arr[7][12] ;
 wire \rvcpu.dp.rf.reg_file_arr[7][13] ;
 wire \rvcpu.dp.rf.reg_file_arr[7][14] ;
 wire \rvcpu.dp.rf.reg_file_arr[7][15] ;
 wire \rvcpu.dp.rf.reg_file_arr[7][16] ;
 wire \rvcpu.dp.rf.reg_file_arr[7][17] ;
 wire \rvcpu.dp.rf.reg_file_arr[7][18] ;
 wire \rvcpu.dp.rf.reg_file_arr[7][19] ;
 wire \rvcpu.dp.rf.reg_file_arr[7][1] ;
 wire \rvcpu.dp.rf.reg_file_arr[7][20] ;
 wire \rvcpu.dp.rf.reg_file_arr[7][21] ;
 wire \rvcpu.dp.rf.reg_file_arr[7][22] ;
 wire \rvcpu.dp.rf.reg_file_arr[7][23] ;
 wire \rvcpu.dp.rf.reg_file_arr[7][24] ;
 wire \rvcpu.dp.rf.reg_file_arr[7][25] ;
 wire \rvcpu.dp.rf.reg_file_arr[7][26] ;
 wire \rvcpu.dp.rf.reg_file_arr[7][27] ;
 wire \rvcpu.dp.rf.reg_file_arr[7][28] ;
 wire \rvcpu.dp.rf.reg_file_arr[7][29] ;
 wire \rvcpu.dp.rf.reg_file_arr[7][2] ;
 wire \rvcpu.dp.rf.reg_file_arr[7][30] ;
 wire \rvcpu.dp.rf.reg_file_arr[7][31] ;
 wire \rvcpu.dp.rf.reg_file_arr[7][3] ;
 wire \rvcpu.dp.rf.reg_file_arr[7][4] ;
 wire \rvcpu.dp.rf.reg_file_arr[7][5] ;
 wire \rvcpu.dp.rf.reg_file_arr[7][6] ;
 wire \rvcpu.dp.rf.reg_file_arr[7][7] ;
 wire \rvcpu.dp.rf.reg_file_arr[7][8] ;
 wire \rvcpu.dp.rf.reg_file_arr[7][9] ;
 wire \rvcpu.dp.rf.reg_file_arr[8][0] ;
 wire \rvcpu.dp.rf.reg_file_arr[8][10] ;
 wire \rvcpu.dp.rf.reg_file_arr[8][11] ;
 wire \rvcpu.dp.rf.reg_file_arr[8][12] ;
 wire \rvcpu.dp.rf.reg_file_arr[8][13] ;
 wire \rvcpu.dp.rf.reg_file_arr[8][14] ;
 wire \rvcpu.dp.rf.reg_file_arr[8][15] ;
 wire \rvcpu.dp.rf.reg_file_arr[8][16] ;
 wire \rvcpu.dp.rf.reg_file_arr[8][17] ;
 wire \rvcpu.dp.rf.reg_file_arr[8][18] ;
 wire \rvcpu.dp.rf.reg_file_arr[8][19] ;
 wire \rvcpu.dp.rf.reg_file_arr[8][1] ;
 wire \rvcpu.dp.rf.reg_file_arr[8][20] ;
 wire \rvcpu.dp.rf.reg_file_arr[8][21] ;
 wire \rvcpu.dp.rf.reg_file_arr[8][22] ;
 wire \rvcpu.dp.rf.reg_file_arr[8][23] ;
 wire \rvcpu.dp.rf.reg_file_arr[8][24] ;
 wire \rvcpu.dp.rf.reg_file_arr[8][25] ;
 wire \rvcpu.dp.rf.reg_file_arr[8][26] ;
 wire \rvcpu.dp.rf.reg_file_arr[8][27] ;
 wire \rvcpu.dp.rf.reg_file_arr[8][28] ;
 wire \rvcpu.dp.rf.reg_file_arr[8][29] ;
 wire \rvcpu.dp.rf.reg_file_arr[8][2] ;
 wire \rvcpu.dp.rf.reg_file_arr[8][30] ;
 wire \rvcpu.dp.rf.reg_file_arr[8][31] ;
 wire \rvcpu.dp.rf.reg_file_arr[8][3] ;
 wire \rvcpu.dp.rf.reg_file_arr[8][4] ;
 wire \rvcpu.dp.rf.reg_file_arr[8][5] ;
 wire \rvcpu.dp.rf.reg_file_arr[8][6] ;
 wire \rvcpu.dp.rf.reg_file_arr[8][7] ;
 wire \rvcpu.dp.rf.reg_file_arr[8][8] ;
 wire \rvcpu.dp.rf.reg_file_arr[8][9] ;
 wire \rvcpu.dp.rf.reg_file_arr[9][0] ;
 wire \rvcpu.dp.rf.reg_file_arr[9][10] ;
 wire \rvcpu.dp.rf.reg_file_arr[9][11] ;
 wire \rvcpu.dp.rf.reg_file_arr[9][12] ;
 wire \rvcpu.dp.rf.reg_file_arr[9][13] ;
 wire \rvcpu.dp.rf.reg_file_arr[9][14] ;
 wire \rvcpu.dp.rf.reg_file_arr[9][15] ;
 wire \rvcpu.dp.rf.reg_file_arr[9][16] ;
 wire \rvcpu.dp.rf.reg_file_arr[9][17] ;
 wire \rvcpu.dp.rf.reg_file_arr[9][18] ;
 wire \rvcpu.dp.rf.reg_file_arr[9][19] ;
 wire \rvcpu.dp.rf.reg_file_arr[9][1] ;
 wire \rvcpu.dp.rf.reg_file_arr[9][20] ;
 wire \rvcpu.dp.rf.reg_file_arr[9][21] ;
 wire \rvcpu.dp.rf.reg_file_arr[9][22] ;
 wire \rvcpu.dp.rf.reg_file_arr[9][23] ;
 wire \rvcpu.dp.rf.reg_file_arr[9][24] ;
 wire \rvcpu.dp.rf.reg_file_arr[9][25] ;
 wire \rvcpu.dp.rf.reg_file_arr[9][26] ;
 wire \rvcpu.dp.rf.reg_file_arr[9][27] ;
 wire \rvcpu.dp.rf.reg_file_arr[9][28] ;
 wire \rvcpu.dp.rf.reg_file_arr[9][29] ;
 wire \rvcpu.dp.rf.reg_file_arr[9][2] ;
 wire \rvcpu.dp.rf.reg_file_arr[9][30] ;
 wire \rvcpu.dp.rf.reg_file_arr[9][31] ;
 wire \rvcpu.dp.rf.reg_file_arr[9][3] ;
 wire \rvcpu.dp.rf.reg_file_arr[9][4] ;
 wire \rvcpu.dp.rf.reg_file_arr[9][5] ;
 wire \rvcpu.dp.rf.reg_file_arr[9][6] ;
 wire \rvcpu.dp.rf.reg_file_arr[9][7] ;
 wire \rvcpu.dp.rf.reg_file_arr[9][8] ;
 wire \rvcpu.dp.rf.reg_file_arr[9][9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;

 sky130_fd_sc_hd__clkbuf_8 _14583_ (.A(\rvcpu.dp.plmw.ResultSrcW[0] ),
    .X(_13168_));
 sky130_fd_sc_hd__clkbuf_8 _14584_ (.A(_13168_),
    .X(_13169_));
 sky130_fd_sc_hd__buf_4 _14585_ (.A(\rvcpu.dp.plmw.ResultSrcW[1] ),
    .X(_13170_));
 sky130_fd_sc_hd__clkbuf_4 _14586_ (.A(_13170_),
    .X(_13171_));
 sky130_fd_sc_hd__mux4_2 _14587_ (.A0(\rvcpu.dp.plmw.ALUResultW[31] ),
    .A1(\rvcpu.dp.plmw.ReadDataW[31] ),
    .A2(\rvcpu.dp.plmw.PCPlus4W[31] ),
    .A3(\rvcpu.dp.plmw.lAuiPCW[31] ),
    .S0(_13169_),
    .S1(_13171_),
    .X(_13172_));
 sky130_fd_sc_hd__buf_4 _14588_ (.A(_13172_),
    .X(_13173_));
 sky130_fd_sc_hd__clkbuf_4 _14589_ (.A(\rvcpu.dp.plmw.RdW[2] ),
    .X(_13174_));
 sky130_fd_sc_hd__inv_2 _14590_ (.A(\rvcpu.dp.plmw.RdW[3] ),
    .Y(_13175_));
 sky130_fd_sc_hd__clkbuf_4 _14591_ (.A(\rvcpu.dp.plmw.RdW[4] ),
    .X(_13176_));
 sky130_fd_sc_hd__or3_4 _14592_ (.A(_13174_),
    .B(_13175_),
    .C(_13176_),
    .X(_13177_));
 sky130_fd_sc_hd__nand2_2 _14593_ (.A(\rvcpu.dp.plmw.RegWriteW ),
    .B(\rvcpu.dp.plmw.RdW[0] ),
    .Y(_13178_));
 sky130_fd_sc_hd__or2_4 _14594_ (.A(\rvcpu.dp.plmw.RdW[1] ),
    .B(_13178_),
    .X(_13179_));
 sky130_fd_sc_hd__nor2_2 _14595_ (.A(_13177_),
    .B(_13179_),
    .Y(_13180_));
 sky130_fd_sc_hd__buf_4 _14596_ (.A(_13180_),
    .X(_13181_));
 sky130_fd_sc_hd__mux2_1 _14597_ (.A0(\rvcpu.dp.rf.reg_file_arr[9][31] ),
    .A1(_13173_),
    .S(_13181_),
    .X(_13182_));
 sky130_fd_sc_hd__clkbuf_1 _14598_ (.A(_13182_),
    .X(_03203_));
 sky130_fd_sc_hd__mux4_2 _14599_ (.A0(\rvcpu.dp.plmw.ALUResultW[30] ),
    .A1(\rvcpu.dp.plmw.ReadDataW[30] ),
    .A2(\rvcpu.dp.plmw.PCPlus4W[30] ),
    .A3(\rvcpu.dp.plmw.lAuiPCW[30] ),
    .S0(_13168_),
    .S1(_13170_),
    .X(_13183_));
 sky130_fd_sc_hd__buf_4 _14600_ (.A(_13183_),
    .X(_13184_));
 sky130_fd_sc_hd__mux2_1 _14601_ (.A0(\rvcpu.dp.rf.reg_file_arr[9][30] ),
    .A1(_13184_),
    .S(_13181_),
    .X(_13185_));
 sky130_fd_sc_hd__clkbuf_1 _14602_ (.A(_13185_),
    .X(_03202_));
 sky130_fd_sc_hd__mux4_2 _14603_ (.A0(\rvcpu.dp.plmw.ALUResultW[29] ),
    .A1(\rvcpu.dp.plmw.ReadDataW[29] ),
    .A2(\rvcpu.dp.plmw.PCPlus4W[29] ),
    .A3(\rvcpu.dp.plmw.lAuiPCW[29] ),
    .S0(_13168_),
    .S1(_13170_),
    .X(_13186_));
 sky130_fd_sc_hd__buf_4 _14604_ (.A(_13186_),
    .X(_13187_));
 sky130_fd_sc_hd__mux2_1 _14605_ (.A0(\rvcpu.dp.rf.reg_file_arr[9][29] ),
    .A1(_13187_),
    .S(_13181_),
    .X(_13188_));
 sky130_fd_sc_hd__clkbuf_1 _14606_ (.A(_13188_),
    .X(_03201_));
 sky130_fd_sc_hd__mux4_2 _14607_ (.A0(\rvcpu.dp.plmw.ALUResultW[28] ),
    .A1(\rvcpu.dp.plmw.ReadDataW[28] ),
    .A2(\rvcpu.dp.plmw.PCPlus4W[28] ),
    .A3(\rvcpu.dp.plmw.lAuiPCW[28] ),
    .S0(_13168_),
    .S1(_13170_),
    .X(_13189_));
 sky130_fd_sc_hd__buf_4 _14608_ (.A(_13189_),
    .X(_13190_));
 sky130_fd_sc_hd__mux2_1 _14609_ (.A0(\rvcpu.dp.rf.reg_file_arr[9][28] ),
    .A1(_13190_),
    .S(_13181_),
    .X(_13191_));
 sky130_fd_sc_hd__clkbuf_1 _14610_ (.A(_13191_),
    .X(_03200_));
 sky130_fd_sc_hd__clkbuf_8 _14611_ (.A(_13168_),
    .X(_13192_));
 sky130_fd_sc_hd__buf_4 _14612_ (.A(_13170_),
    .X(_13193_));
 sky130_fd_sc_hd__mux4_2 _14613_ (.A0(\rvcpu.dp.plmw.ALUResultW[27] ),
    .A1(\rvcpu.dp.plmw.ReadDataW[27] ),
    .A2(\rvcpu.dp.plmw.PCPlus4W[27] ),
    .A3(\rvcpu.dp.plmw.lAuiPCW[27] ),
    .S0(_13192_),
    .S1(_13193_),
    .X(_13194_));
 sky130_fd_sc_hd__buf_4 _14614_ (.A(_13194_),
    .X(_13195_));
 sky130_fd_sc_hd__mux2_1 _14615_ (.A0(\rvcpu.dp.rf.reg_file_arr[9][27] ),
    .A1(_13195_),
    .S(_13181_),
    .X(_13196_));
 sky130_fd_sc_hd__clkbuf_1 _14616_ (.A(_13196_),
    .X(_03199_));
 sky130_fd_sc_hd__mux4_2 _14617_ (.A0(\rvcpu.dp.plmw.ALUResultW[26] ),
    .A1(\rvcpu.dp.plmw.ReadDataW[26] ),
    .A2(\rvcpu.dp.plmw.PCPlus4W[26] ),
    .A3(\rvcpu.dp.plmw.lAuiPCW[26] ),
    .S0(_13192_),
    .S1(_13193_),
    .X(_13197_));
 sky130_fd_sc_hd__buf_4 _14618_ (.A(_13197_),
    .X(_13198_));
 sky130_fd_sc_hd__mux2_1 _14619_ (.A0(\rvcpu.dp.rf.reg_file_arr[9][26] ),
    .A1(_13198_),
    .S(_13181_),
    .X(_13199_));
 sky130_fd_sc_hd__clkbuf_1 _14620_ (.A(_13199_),
    .X(_03198_));
 sky130_fd_sc_hd__mux4_2 _14621_ (.A0(\rvcpu.dp.plmw.ALUResultW[25] ),
    .A1(\rvcpu.dp.plmw.ReadDataW[25] ),
    .A2(\rvcpu.dp.plmw.PCPlus4W[25] ),
    .A3(\rvcpu.dp.plmw.lAuiPCW[25] ),
    .S0(_13192_),
    .S1(_13193_),
    .X(_13200_));
 sky130_fd_sc_hd__buf_4 _14622_ (.A(_13200_),
    .X(_13201_));
 sky130_fd_sc_hd__mux2_1 _14623_ (.A0(\rvcpu.dp.rf.reg_file_arr[9][25] ),
    .A1(_13201_),
    .S(_13181_),
    .X(_13202_));
 sky130_fd_sc_hd__clkbuf_1 _14624_ (.A(_13202_),
    .X(_03197_));
 sky130_fd_sc_hd__mux4_2 _14625_ (.A0(\rvcpu.dp.plmw.ALUResultW[24] ),
    .A1(\rvcpu.dp.plmw.ReadDataW[24] ),
    .A2(\rvcpu.dp.plmw.PCPlus4W[24] ),
    .A3(\rvcpu.dp.plmw.lAuiPCW[24] ),
    .S0(_13192_),
    .S1(_13193_),
    .X(_13203_));
 sky130_fd_sc_hd__buf_4 _14626_ (.A(_13203_),
    .X(_13204_));
 sky130_fd_sc_hd__mux2_1 _14627_ (.A0(\rvcpu.dp.rf.reg_file_arr[9][24] ),
    .A1(_13204_),
    .S(_13181_),
    .X(_13205_));
 sky130_fd_sc_hd__clkbuf_1 _14628_ (.A(_13205_),
    .X(_03196_));
 sky130_fd_sc_hd__mux4_2 _14629_ (.A0(\rvcpu.dp.plmw.ALUResultW[23] ),
    .A1(\rvcpu.dp.plmw.ReadDataW[23] ),
    .A2(\rvcpu.dp.plmw.PCPlus4W[23] ),
    .A3(\rvcpu.dp.plmw.lAuiPCW[23] ),
    .S0(_13169_),
    .S1(_13171_),
    .X(_13206_));
 sky130_fd_sc_hd__buf_4 _14630_ (.A(_13206_),
    .X(_13207_));
 sky130_fd_sc_hd__mux2_1 _14631_ (.A0(\rvcpu.dp.rf.reg_file_arr[9][23] ),
    .A1(_13207_),
    .S(_13181_),
    .X(_13208_));
 sky130_fd_sc_hd__clkbuf_1 _14632_ (.A(_13208_),
    .X(_03195_));
 sky130_fd_sc_hd__mux4_2 _14633_ (.A0(\rvcpu.dp.plmw.ALUResultW[22] ),
    .A1(\rvcpu.dp.plmw.ReadDataW[22] ),
    .A2(\rvcpu.dp.plmw.PCPlus4W[22] ),
    .A3(\rvcpu.dp.plmw.lAuiPCW[22] ),
    .S0(_13169_),
    .S1(_13171_),
    .X(_13209_));
 sky130_fd_sc_hd__buf_4 _14634_ (.A(_13209_),
    .X(_13210_));
 sky130_fd_sc_hd__mux2_1 _14635_ (.A0(\rvcpu.dp.rf.reg_file_arr[9][22] ),
    .A1(_13210_),
    .S(_13181_),
    .X(_13211_));
 sky130_fd_sc_hd__clkbuf_1 _14636_ (.A(_13211_),
    .X(_03194_));
 sky130_fd_sc_hd__mux4_2 _14637_ (.A0(\rvcpu.dp.plmw.ALUResultW[21] ),
    .A1(\rvcpu.dp.plmw.ReadDataW[21] ),
    .A2(\rvcpu.dp.plmw.PCPlus4W[21] ),
    .A3(\rvcpu.dp.plmw.lAuiPCW[21] ),
    .S0(_13169_),
    .S1(_13171_),
    .X(_13212_));
 sky130_fd_sc_hd__clkbuf_8 _14638_ (.A(_13212_),
    .X(_13213_));
 sky130_fd_sc_hd__clkbuf_4 _14639_ (.A(_13180_),
    .X(_13214_));
 sky130_fd_sc_hd__mux2_1 _14640_ (.A0(\rvcpu.dp.rf.reg_file_arr[9][21] ),
    .A1(_13213_),
    .S(_13214_),
    .X(_13215_));
 sky130_fd_sc_hd__clkbuf_1 _14641_ (.A(_13215_),
    .X(_03193_));
 sky130_fd_sc_hd__mux4_2 _14642_ (.A0(\rvcpu.dp.plmw.ALUResultW[20] ),
    .A1(\rvcpu.dp.plmw.ReadDataW[20] ),
    .A2(\rvcpu.dp.plmw.PCPlus4W[20] ),
    .A3(\rvcpu.dp.plmw.lAuiPCW[20] ),
    .S0(_13169_),
    .S1(_13171_),
    .X(_13216_));
 sky130_fd_sc_hd__clkbuf_8 _14643_ (.A(_13216_),
    .X(_13217_));
 sky130_fd_sc_hd__mux2_1 _14644_ (.A0(\rvcpu.dp.rf.reg_file_arr[9][20] ),
    .A1(_13217_),
    .S(_13214_),
    .X(_13218_));
 sky130_fd_sc_hd__clkbuf_1 _14645_ (.A(_13218_),
    .X(_03192_));
 sky130_fd_sc_hd__mux4_2 _14646_ (.A0(\rvcpu.dp.plmw.ALUResultW[19] ),
    .A1(\rvcpu.dp.plmw.ReadDataW[19] ),
    .A2(\rvcpu.dp.plmw.PCPlus4W[19] ),
    .A3(\rvcpu.dp.plmw.lAuiPCW[19] ),
    .S0(_13169_),
    .S1(_13171_),
    .X(_13219_));
 sky130_fd_sc_hd__clkbuf_8 _14647_ (.A(_13219_),
    .X(_13220_));
 sky130_fd_sc_hd__mux2_1 _14648_ (.A0(\rvcpu.dp.rf.reg_file_arr[9][19] ),
    .A1(_13220_),
    .S(_13214_),
    .X(_13221_));
 sky130_fd_sc_hd__clkbuf_1 _14649_ (.A(_13221_),
    .X(_03191_));
 sky130_fd_sc_hd__mux4_2 _14650_ (.A0(\rvcpu.dp.plmw.ALUResultW[18] ),
    .A1(\rvcpu.dp.plmw.ReadDataW[18] ),
    .A2(\rvcpu.dp.plmw.PCPlus4W[18] ),
    .A3(\rvcpu.dp.plmw.lAuiPCW[18] ),
    .S0(_13192_),
    .S1(_13193_),
    .X(_13222_));
 sky130_fd_sc_hd__clkbuf_8 _14651_ (.A(_13222_),
    .X(_13223_));
 sky130_fd_sc_hd__mux2_1 _14652_ (.A0(\rvcpu.dp.rf.reg_file_arr[9][18] ),
    .A1(_13223_),
    .S(_13214_),
    .X(_13224_));
 sky130_fd_sc_hd__clkbuf_1 _14653_ (.A(_13224_),
    .X(_03190_));
 sky130_fd_sc_hd__mux4_2 _14654_ (.A0(\rvcpu.dp.plmw.ALUResultW[17] ),
    .A1(\rvcpu.dp.plmw.ReadDataW[17] ),
    .A2(\rvcpu.dp.plmw.PCPlus4W[17] ),
    .A3(\rvcpu.dp.plmw.lAuiPCW[17] ),
    .S0(_13169_),
    .S1(_13171_),
    .X(_13225_));
 sky130_fd_sc_hd__buf_4 _14655_ (.A(_13225_),
    .X(_13226_));
 sky130_fd_sc_hd__mux2_1 _14656_ (.A0(\rvcpu.dp.rf.reg_file_arr[9][17] ),
    .A1(_13226_),
    .S(_13214_),
    .X(_13227_));
 sky130_fd_sc_hd__clkbuf_1 _14657_ (.A(_13227_),
    .X(_03189_));
 sky130_fd_sc_hd__mux4_2 _14658_ (.A0(\rvcpu.dp.plmw.ALUResultW[16] ),
    .A1(\rvcpu.dp.plmw.ReadDataW[16] ),
    .A2(\rvcpu.dp.plmw.PCPlus4W[16] ),
    .A3(\rvcpu.dp.plmw.lAuiPCW[16] ),
    .S0(_13192_),
    .S1(_13193_),
    .X(_13228_));
 sky130_fd_sc_hd__clkbuf_8 _14659_ (.A(_13228_),
    .X(_13229_));
 sky130_fd_sc_hd__mux2_1 _14660_ (.A0(\rvcpu.dp.rf.reg_file_arr[9][16] ),
    .A1(_13229_),
    .S(_13214_),
    .X(_13230_));
 sky130_fd_sc_hd__clkbuf_1 _14661_ (.A(_13230_),
    .X(_03188_));
 sky130_fd_sc_hd__mux4_2 _14662_ (.A0(\rvcpu.dp.plmw.ALUResultW[15] ),
    .A1(\rvcpu.dp.plmw.ReadDataW[15] ),
    .A2(\rvcpu.dp.plmw.PCPlus4W[15] ),
    .A3(\rvcpu.dp.plmw.lAuiPCW[15] ),
    .S0(_13168_),
    .S1(_13170_),
    .X(_13231_));
 sky130_fd_sc_hd__buf_4 _14663_ (.A(_13231_),
    .X(_13232_));
 sky130_fd_sc_hd__mux2_1 _14664_ (.A0(\rvcpu.dp.rf.reg_file_arr[9][15] ),
    .A1(_13232_),
    .S(_13214_),
    .X(_13233_));
 sky130_fd_sc_hd__clkbuf_1 _14665_ (.A(_13233_),
    .X(_03187_));
 sky130_fd_sc_hd__mux4_2 _14666_ (.A0(\rvcpu.dp.plmw.ALUResultW[14] ),
    .A1(\rvcpu.dp.plmw.ReadDataW[14] ),
    .A2(\rvcpu.dp.plmw.PCPlus4W[14] ),
    .A3(\rvcpu.dp.plmw.lAuiPCW[14] ),
    .S0(_13192_),
    .S1(_13193_),
    .X(_13234_));
 sky130_fd_sc_hd__buf_4 _14667_ (.A(_13234_),
    .X(_13235_));
 sky130_fd_sc_hd__mux2_1 _14668_ (.A0(\rvcpu.dp.rf.reg_file_arr[9][14] ),
    .A1(_13235_),
    .S(_13214_),
    .X(_13236_));
 sky130_fd_sc_hd__clkbuf_1 _14669_ (.A(_13236_),
    .X(_03186_));
 sky130_fd_sc_hd__mux4_2 _14670_ (.A0(\rvcpu.dp.plmw.ALUResultW[13] ),
    .A1(\rvcpu.dp.plmw.ReadDataW[13] ),
    .A2(\rvcpu.dp.plmw.PCPlus4W[13] ),
    .A3(\rvcpu.dp.plmw.lAuiPCW[13] ),
    .S0(_13169_),
    .S1(_13171_),
    .X(_13237_));
 sky130_fd_sc_hd__buf_4 _14671_ (.A(_13237_),
    .X(_13238_));
 sky130_fd_sc_hd__mux2_1 _14672_ (.A0(\rvcpu.dp.rf.reg_file_arr[9][13] ),
    .A1(_13238_),
    .S(_13214_),
    .X(_13239_));
 sky130_fd_sc_hd__clkbuf_1 _14673_ (.A(_13239_),
    .X(_03185_));
 sky130_fd_sc_hd__mux4_2 _14674_ (.A0(\rvcpu.dp.plmw.ALUResultW[12] ),
    .A1(\rvcpu.dp.plmw.ReadDataW[12] ),
    .A2(\rvcpu.dp.plmw.PCPlus4W[12] ),
    .A3(\rvcpu.dp.plmw.lAuiPCW[12] ),
    .S0(_13168_),
    .S1(_13170_),
    .X(_13240_));
 sky130_fd_sc_hd__buf_4 _14675_ (.A(_13240_),
    .X(_13241_));
 sky130_fd_sc_hd__mux2_1 _14676_ (.A0(\rvcpu.dp.rf.reg_file_arr[9][12] ),
    .A1(_13241_),
    .S(_13214_),
    .X(_13242_));
 sky130_fd_sc_hd__clkbuf_1 _14677_ (.A(_13242_),
    .X(_03184_));
 sky130_fd_sc_hd__mux4_2 _14678_ (.A0(\rvcpu.dp.plmw.ALUResultW[11] ),
    .A1(\rvcpu.dp.plmw.ReadDataW[11] ),
    .A2(\rvcpu.dp.plmw.PCPlus4W[11] ),
    .A3(\rvcpu.dp.plmw.lAuiPCW[11] ),
    .S0(_13168_),
    .S1(_13170_),
    .X(_13243_));
 sky130_fd_sc_hd__clkbuf_8 _14679_ (.A(_13243_),
    .X(_13244_));
 sky130_fd_sc_hd__buf_4 _14680_ (.A(_13180_),
    .X(_13245_));
 sky130_fd_sc_hd__mux2_1 _14681_ (.A0(\rvcpu.dp.rf.reg_file_arr[9][11] ),
    .A1(_13244_),
    .S(_13245_),
    .X(_13246_));
 sky130_fd_sc_hd__clkbuf_1 _14682_ (.A(_13246_),
    .X(_03183_));
 sky130_fd_sc_hd__mux4_2 _14683_ (.A0(\rvcpu.dp.plmw.ALUResultW[10] ),
    .A1(\rvcpu.dp.plmw.ReadDataW[10] ),
    .A2(\rvcpu.dp.plmw.PCPlus4W[10] ),
    .A3(\rvcpu.dp.plmw.lAuiPCW[10] ),
    .S0(_13169_),
    .S1(_13171_),
    .X(_13247_));
 sky130_fd_sc_hd__clkbuf_8 _14684_ (.A(_13247_),
    .X(_13248_));
 sky130_fd_sc_hd__mux2_1 _14685_ (.A0(\rvcpu.dp.rf.reg_file_arr[9][10] ),
    .A1(_13248_),
    .S(_13245_),
    .X(_13249_));
 sky130_fd_sc_hd__clkbuf_1 _14686_ (.A(_13249_),
    .X(_03182_));
 sky130_fd_sc_hd__mux4_2 _14687_ (.A0(\rvcpu.dp.plmw.ALUResultW[9] ),
    .A1(\rvcpu.dp.plmw.ReadDataW[9] ),
    .A2(\rvcpu.dp.plmw.PCPlus4W[9] ),
    .A3(\rvcpu.dp.plmw.lAuiPCW[9] ),
    .S0(_13168_),
    .S1(_13170_),
    .X(_13250_));
 sky130_fd_sc_hd__clkbuf_8 _14688_ (.A(_13250_),
    .X(_13251_));
 sky130_fd_sc_hd__mux2_1 _14689_ (.A0(\rvcpu.dp.rf.reg_file_arr[9][9] ),
    .A1(_13251_),
    .S(_13245_),
    .X(_13252_));
 sky130_fd_sc_hd__clkbuf_1 _14690_ (.A(_13252_),
    .X(_03181_));
 sky130_fd_sc_hd__mux4_2 _14691_ (.A0(\rvcpu.dp.plmw.ALUResultW[8] ),
    .A1(\rvcpu.dp.plmw.ReadDataW[8] ),
    .A2(\rvcpu.dp.plmw.PCPlus4W[8] ),
    .A3(\rvcpu.dp.plmw.lAuiPCW[8] ),
    .S0(_13169_),
    .S1(_13171_),
    .X(_13253_));
 sky130_fd_sc_hd__clkbuf_8 _14692_ (.A(_13253_),
    .X(_13254_));
 sky130_fd_sc_hd__mux2_1 _14693_ (.A0(\rvcpu.dp.rf.reg_file_arr[9][8] ),
    .A1(_13254_),
    .S(_13245_),
    .X(_13255_));
 sky130_fd_sc_hd__clkbuf_1 _14694_ (.A(_13255_),
    .X(_03180_));
 sky130_fd_sc_hd__mux4_2 _14695_ (.A0(\rvcpu.dp.plmw.ALUResultW[7] ),
    .A1(\rvcpu.dp.plmw.ReadDataW[7] ),
    .A2(\rvcpu.dp.plmw.PCPlus4W[7] ),
    .A3(\rvcpu.dp.plmw.lAuiPCW[7] ),
    .S0(_13192_),
    .S1(_13193_),
    .X(_13256_));
 sky130_fd_sc_hd__clkbuf_8 _14696_ (.A(_13256_),
    .X(_13257_));
 sky130_fd_sc_hd__mux2_1 _14697_ (.A0(\rvcpu.dp.rf.reg_file_arr[9][7] ),
    .A1(_13257_),
    .S(_13245_),
    .X(_13258_));
 sky130_fd_sc_hd__clkbuf_1 _14698_ (.A(_13258_),
    .X(_03179_));
 sky130_fd_sc_hd__mux4_2 _14699_ (.A0(\rvcpu.dp.plmw.ALUResultW[6] ),
    .A1(\rvcpu.dp.plmw.ReadDataW[6] ),
    .A2(\rvcpu.dp.plmw.PCPlus4W[6] ),
    .A3(\rvcpu.dp.plmw.lAuiPCW[6] ),
    .S0(_13192_),
    .S1(_13193_),
    .X(_13259_));
 sky130_fd_sc_hd__clkbuf_8 _14700_ (.A(_13259_),
    .X(_13260_));
 sky130_fd_sc_hd__mux2_1 _14701_ (.A0(\rvcpu.dp.rf.reg_file_arr[9][6] ),
    .A1(_13260_),
    .S(_13245_),
    .X(_13261_));
 sky130_fd_sc_hd__clkbuf_1 _14702_ (.A(_13261_),
    .X(_03178_));
 sky130_fd_sc_hd__mux4_2 _14703_ (.A0(\rvcpu.dp.plmw.ALUResultW[5] ),
    .A1(\rvcpu.dp.plmw.ReadDataW[5] ),
    .A2(\rvcpu.dp.plmw.PCPlus4W[5] ),
    .A3(\rvcpu.dp.plmw.lAuiPCW[5] ),
    .S0(_13192_),
    .S1(_13193_),
    .X(_13262_));
 sky130_fd_sc_hd__buf_4 _14704_ (.A(_13262_),
    .X(_13263_));
 sky130_fd_sc_hd__mux2_1 _14705_ (.A0(\rvcpu.dp.rf.reg_file_arr[9][5] ),
    .A1(_13263_),
    .S(_13245_),
    .X(_13264_));
 sky130_fd_sc_hd__clkbuf_1 _14706_ (.A(_13264_),
    .X(_03177_));
 sky130_fd_sc_hd__mux4_2 _14707_ (.A0(\rvcpu.dp.plmw.ALUResultW[4] ),
    .A1(\rvcpu.dp.plmw.ReadDataW[4] ),
    .A2(\rvcpu.dp.plmw.PCPlus4W[4] ),
    .A3(\rvcpu.dp.plmw.lAuiPCW[4] ),
    .S0(_13168_),
    .S1(_13170_),
    .X(_13265_));
 sky130_fd_sc_hd__clkbuf_8 _14708_ (.A(_13265_),
    .X(_13266_));
 sky130_fd_sc_hd__mux2_1 _14709_ (.A0(\rvcpu.dp.rf.reg_file_arr[9][4] ),
    .A1(_13266_),
    .S(_13245_),
    .X(_13267_));
 sky130_fd_sc_hd__clkbuf_1 _14710_ (.A(_13267_),
    .X(_03176_));
 sky130_fd_sc_hd__mux4_2 _14711_ (.A0(\rvcpu.dp.plmw.ALUResultW[3] ),
    .A1(\rvcpu.dp.plmw.ReadDataW[3] ),
    .A2(\rvcpu.dp.plmw.PCPlus4W[3] ),
    .A3(\rvcpu.dp.plmw.lAuiPCW[3] ),
    .S0(\rvcpu.dp.plmw.ResultSrcW[0] ),
    .S1(\rvcpu.dp.plmw.ResultSrcW[1] ),
    .X(_13268_));
 sky130_fd_sc_hd__clkbuf_8 _14712_ (.A(_13268_),
    .X(_13269_));
 sky130_fd_sc_hd__mux2_1 _14713_ (.A0(\rvcpu.dp.rf.reg_file_arr[9][3] ),
    .A1(_13269_),
    .S(_13245_),
    .X(_13270_));
 sky130_fd_sc_hd__clkbuf_1 _14714_ (.A(_13270_),
    .X(_03175_));
 sky130_fd_sc_hd__mux4_2 _14715_ (.A0(\rvcpu.dp.plmw.ALUResultW[2] ),
    .A1(\rvcpu.dp.plmw.ReadDataW[2] ),
    .A2(\rvcpu.dp.plmw.PCPlus4W[2] ),
    .A3(\rvcpu.dp.plmw.lAuiPCW[2] ),
    .S0(\rvcpu.dp.plmw.ResultSrcW[0] ),
    .S1(\rvcpu.dp.plmw.ResultSrcW[1] ),
    .X(_13271_));
 sky130_fd_sc_hd__buf_4 _14716_ (.A(_13271_),
    .X(_13272_));
 sky130_fd_sc_hd__mux2_1 _14717_ (.A0(\rvcpu.dp.rf.reg_file_arr[9][2] ),
    .A1(_13272_),
    .S(_13245_),
    .X(_13273_));
 sky130_fd_sc_hd__clkbuf_1 _14718_ (.A(_13273_),
    .X(_03174_));
 sky130_fd_sc_hd__mux4_2 _14719_ (.A0(\rvcpu.dp.plmw.ALUResultW[1] ),
    .A1(\rvcpu.dp.plmw.ReadDataW[1] ),
    .A2(\rvcpu.dp.plmw.PCPlus4W[1] ),
    .A3(\rvcpu.dp.plmw.lAuiPCW[1] ),
    .S0(\rvcpu.dp.plmw.ResultSrcW[0] ),
    .S1(\rvcpu.dp.plmw.ResultSrcW[1] ),
    .X(_13274_));
 sky130_fd_sc_hd__buf_4 _14720_ (.A(_13274_),
    .X(_13275_));
 sky130_fd_sc_hd__mux2_1 _14721_ (.A0(\rvcpu.dp.rf.reg_file_arr[9][1] ),
    .A1(_13275_),
    .S(_13180_),
    .X(_13276_));
 sky130_fd_sc_hd__clkbuf_1 _14722_ (.A(_13276_),
    .X(_03173_));
 sky130_fd_sc_hd__mux4_2 _14723_ (.A0(\rvcpu.dp.plmw.ALUResultW[0] ),
    .A1(\rvcpu.dp.plmw.ReadDataW[0] ),
    .A2(\rvcpu.dp.plmw.PCPlus4W[0] ),
    .A3(\rvcpu.dp.plmw.lAuiPCW[0] ),
    .S0(\rvcpu.dp.plmw.ResultSrcW[0] ),
    .S1(\rvcpu.dp.plmw.ResultSrcW[1] ),
    .X(_13277_));
 sky130_fd_sc_hd__buf_4 _14724_ (.A(_13277_),
    .X(_13278_));
 sky130_fd_sc_hd__mux2_1 _14725_ (.A0(\rvcpu.dp.rf.reg_file_arr[9][0] ),
    .A1(_13278_),
    .S(_13180_),
    .X(_13279_));
 sky130_fd_sc_hd__clkbuf_1 _14726_ (.A(_13279_),
    .X(_03172_));
 sky130_fd_sc_hd__clkbuf_4 _14727_ (.A(\rvcpu.dp.pcreg.q[2] ),
    .X(_13280_));
 sky130_fd_sc_hd__buf_4 _14728_ (.A(_13280_),
    .X(_13281_));
 sky130_fd_sc_hd__buf_2 _14729_ (.A(_13281_),
    .X(_13282_));
 sky130_fd_sc_hd__inv_2 _14730_ (.A(\rvcpu.dp.pcreg.q[6] ),
    .Y(_13283_));
 sky130_fd_sc_hd__buf_4 _14731_ (.A(\rvcpu.dp.pcreg.q[5] ),
    .X(_13284_));
 sky130_fd_sc_hd__nand2_1 _14732_ (.A(_13283_),
    .B(_13284_),
    .Y(_13285_));
 sky130_fd_sc_hd__buf_2 _14733_ (.A(\rvcpu.dp.pcreg.q[4] ),
    .X(_13286_));
 sky130_fd_sc_hd__buf_4 _14734_ (.A(_13286_),
    .X(_13287_));
 sky130_fd_sc_hd__clkbuf_4 _14735_ (.A(\rvcpu.dp.pcreg.q[3] ),
    .X(_13288_));
 sky130_fd_sc_hd__nand2b_4 _14736_ (.A_N(_13287_),
    .B(_13288_),
    .Y(_13289_));
 sky130_fd_sc_hd__or3_1 _14737_ (.A(_13282_),
    .B(_13285_),
    .C(_13289_),
    .X(_13290_));
 sky130_fd_sc_hd__clkbuf_4 _14738_ (.A(_13283_),
    .X(_13291_));
 sky130_fd_sc_hd__clkbuf_4 _14739_ (.A(_13291_),
    .X(_13292_));
 sky130_fd_sc_hd__and2_1 _14740_ (.A(\rvcpu.dp.pcreg.q[5] ),
    .B(_13281_),
    .X(_13293_));
 sky130_fd_sc_hd__clkbuf_4 _14741_ (.A(_13293_),
    .X(_13294_));
 sky130_fd_sc_hd__inv_2 _14742_ (.A(\rvcpu.dp.pcreg.q[5] ),
    .Y(_13295_));
 sky130_fd_sc_hd__buf_4 _14743_ (.A(_13295_),
    .X(_13296_));
 sky130_fd_sc_hd__clkbuf_4 _14744_ (.A(_13296_),
    .X(_13297_));
 sky130_fd_sc_hd__clkbuf_4 _14745_ (.A(_13297_),
    .X(_13298_));
 sky130_fd_sc_hd__and2_1 _14746_ (.A(_13286_),
    .B(\rvcpu.dp.pcreg.q[3] ),
    .X(_13299_));
 sky130_fd_sc_hd__buf_2 _14747_ (.A(_13299_),
    .X(_13300_));
 sky130_fd_sc_hd__clkbuf_4 _14748_ (.A(_13300_),
    .X(_13301_));
 sky130_fd_sc_hd__nor2_1 _14749_ (.A(_13298_),
    .B(_13301_),
    .Y(_13302_));
 sky130_fd_sc_hd__buf_4 _14750_ (.A(_13284_),
    .X(_13303_));
 sky130_fd_sc_hd__clkbuf_4 _14751_ (.A(_13303_),
    .X(_13304_));
 sky130_fd_sc_hd__buf_4 _14752_ (.A(_13288_),
    .X(_13305_));
 sky130_fd_sc_hd__or2_1 _14753_ (.A(\rvcpu.dp.pcreg.q[4] ),
    .B(\rvcpu.dp.pcreg.q[2] ),
    .X(_13306_));
 sky130_fd_sc_hd__buf_4 _14754_ (.A(_13306_),
    .X(_13307_));
 sky130_fd_sc_hd__nor2_4 _14755_ (.A(_13305_),
    .B(_13307_),
    .Y(_13308_));
 sky130_fd_sc_hd__nor2_2 _14756_ (.A(_13304_),
    .B(_13308_),
    .Y(_13309_));
 sky130_fd_sc_hd__or4_1 _14757_ (.A(_13292_),
    .B(_13294_),
    .C(_13302_),
    .D(_13309_),
    .X(_13310_));
 sky130_fd_sc_hd__inv_2 _14758_ (.A(\rvcpu.dp.pcreg.q[8] ),
    .Y(_13311_));
 sky130_fd_sc_hd__clkbuf_4 _14759_ (.A(_13311_),
    .X(_13312_));
 sky130_fd_sc_hd__clkbuf_4 _14760_ (.A(\rvcpu.dp.pcreg.q[7] ),
    .X(_13313_));
 sky130_fd_sc_hd__clkbuf_4 _14761_ (.A(_13313_),
    .X(_13314_));
 sky130_fd_sc_hd__nand2_2 _14762_ (.A(_13312_),
    .B(_13314_),
    .Y(_13315_));
 sky130_fd_sc_hd__a21oi_1 _14763_ (.A1(_13290_),
    .A2(_13310_),
    .B1(_13315_),
    .Y(_13316_));
 sky130_fd_sc_hd__nor2_2 _14764_ (.A(\rvcpu.dp.pcreg.q[6] ),
    .B(\rvcpu.dp.pcreg.q[5] ),
    .Y(_13317_));
 sky130_fd_sc_hd__and2_1 _14765_ (.A(\rvcpu.dp.pcreg.q[8] ),
    .B(_13313_),
    .X(_13318_));
 sky130_fd_sc_hd__clkbuf_4 _14766_ (.A(_13318_),
    .X(_13319_));
 sky130_fd_sc_hd__clkbuf_4 _14767_ (.A(_13305_),
    .X(_13320_));
 sky130_fd_sc_hd__nor2b_4 _14768_ (.A(_13280_),
    .B_N(_13286_),
    .Y(_13321_));
 sky130_fd_sc_hd__nor2b_4 _14769_ (.A(_13286_),
    .B_N(_13280_),
    .Y(_13322_));
 sky130_fd_sc_hd__nor2_4 _14770_ (.A(_13321_),
    .B(_13322_),
    .Y(_13323_));
 sky130_fd_sc_hd__nor2_4 _14771_ (.A(_13320_),
    .B(_13323_),
    .Y(_13324_));
 sky130_fd_sc_hd__a31o_1 _14772_ (.A1(_13317_),
    .A2(_13319_),
    .A3(_13324_),
    .B1(\rvcpu.dp.pcreg.q[9] ),
    .X(_13325_));
 sky130_fd_sc_hd__nor2_2 _14773_ (.A(_13312_),
    .B(_13314_),
    .Y(_13326_));
 sky130_fd_sc_hd__clkbuf_4 _14774_ (.A(_13326_),
    .X(_13327_));
 sky130_fd_sc_hd__clkbuf_4 _14775_ (.A(_13282_),
    .X(_13328_));
 sky130_fd_sc_hd__nand2_1 _14776_ (.A(_13296_),
    .B(_13300_),
    .Y(_13329_));
 sky130_fd_sc_hd__or2_2 _14777_ (.A(_13283_),
    .B(_13329_),
    .X(_13330_));
 sky130_fd_sc_hd__clkbuf_4 _14778_ (.A(\rvcpu.dp.pcreg.q[6] ),
    .X(_13331_));
 sky130_fd_sc_hd__clkbuf_4 _14779_ (.A(_13331_),
    .X(_13332_));
 sky130_fd_sc_hd__clkbuf_4 _14780_ (.A(_13332_),
    .X(_13333_));
 sky130_fd_sc_hd__or2b_1 _14781_ (.A(_13288_),
    .B_N(_13286_),
    .X(_13334_));
 sky130_fd_sc_hd__clkbuf_4 _14782_ (.A(_13334_),
    .X(_13335_));
 sky130_fd_sc_hd__nand2_8 _14783_ (.A(\rvcpu.dp.pcreg.q[5] ),
    .B(\rvcpu.dp.pcreg.q[2] ),
    .Y(_13336_));
 sky130_fd_sc_hd__nor2_2 _14784_ (.A(_13335_),
    .B(_13336_),
    .Y(_13337_));
 sky130_fd_sc_hd__nand2_1 _14785_ (.A(_13333_),
    .B(_13337_),
    .Y(_13338_));
 sky130_fd_sc_hd__o21ai_1 _14786_ (.A1(_13328_),
    .A2(_13330_),
    .B1(_13338_),
    .Y(_13339_));
 sky130_fd_sc_hd__and2b_1 _14787_ (.A_N(_13288_),
    .B(_13286_),
    .X(_13340_));
 sky130_fd_sc_hd__clkbuf_4 _14788_ (.A(_13340_),
    .X(_13341_));
 sky130_fd_sc_hd__and2_1 _14789_ (.A(_13296_),
    .B(_13281_),
    .X(_13342_));
 sky130_fd_sc_hd__buf_2 _14790_ (.A(_13342_),
    .X(_13343_));
 sky130_fd_sc_hd__nand2_2 _14791_ (.A(_13341_),
    .B(_13343_),
    .Y(_13344_));
 sky130_fd_sc_hd__or2b_1 _14792_ (.A(_13280_),
    .B_N(_13286_),
    .X(_13345_));
 sky130_fd_sc_hd__clkbuf_4 _14793_ (.A(_13345_),
    .X(_13346_));
 sky130_fd_sc_hd__or2b_1 _14794_ (.A(_13286_),
    .B_N(_13280_),
    .X(_13347_));
 sky130_fd_sc_hd__buf_4 _14795_ (.A(_13347_),
    .X(_13348_));
 sky130_fd_sc_hd__nand2_2 _14796_ (.A(_13346_),
    .B(_13348_),
    .Y(_13349_));
 sky130_fd_sc_hd__nand2_4 _14797_ (.A(_13284_),
    .B(_13305_),
    .Y(_13350_));
 sky130_fd_sc_hd__or2_1 _14798_ (.A(_13349_),
    .B(_13350_),
    .X(_13351_));
 sky130_fd_sc_hd__nor2_1 _14799_ (.A(_13314_),
    .B(_13331_),
    .Y(_13352_));
 sky130_fd_sc_hd__buf_2 _14800_ (.A(_13352_),
    .X(_13353_));
 sky130_fd_sc_hd__nand2_1 _14801_ (.A(_13312_),
    .B(_13353_),
    .Y(_13354_));
 sky130_fd_sc_hd__a21oi_1 _14802_ (.A1(_13344_),
    .A2(_13351_),
    .B1(_13354_),
    .Y(_13355_));
 sky130_fd_sc_hd__or2_1 _14803_ (.A(\rvcpu.dp.pcreg.q[8] ),
    .B(_13313_),
    .X(_13356_));
 sky130_fd_sc_hd__clkbuf_4 _14804_ (.A(_13356_),
    .X(_13357_));
 sky130_fd_sc_hd__clkbuf_4 _14805_ (.A(_13331_),
    .X(_13358_));
 sky130_fd_sc_hd__nor2_2 _14806_ (.A(_13289_),
    .B(_13336_),
    .Y(_13359_));
 sky130_fd_sc_hd__nand2_2 _14807_ (.A(_13358_),
    .B(_13359_),
    .Y(_13360_));
 sky130_fd_sc_hd__nor2_1 _14808_ (.A(_13357_),
    .B(_13360_),
    .Y(_13361_));
 sky130_fd_sc_hd__a211o_1 _14809_ (.A1(_13327_),
    .A2(_13339_),
    .B1(_13355_),
    .C1(_13361_),
    .X(_13362_));
 sky130_fd_sc_hd__nand2_2 _14810_ (.A(_13303_),
    .B(_13308_),
    .Y(_13363_));
 sky130_fd_sc_hd__nand2_2 _14811_ (.A(_13296_),
    .B(_13341_),
    .Y(_13364_));
 sky130_fd_sc_hd__and2_1 _14812_ (.A(_13313_),
    .B(\rvcpu.dp.pcreg.q[6] ),
    .X(_13365_));
 sky130_fd_sc_hd__nand2_4 _14813_ (.A(_13312_),
    .B(_13365_),
    .Y(_13366_));
 sky130_fd_sc_hd__a21oi_1 _14814_ (.A1(_13363_),
    .A2(_13364_),
    .B1(_13366_),
    .Y(_13367_));
 sky130_fd_sc_hd__buf_4 _14815_ (.A(_13312_),
    .X(_13368_));
 sky130_fd_sc_hd__nand2_4 _14816_ (.A(_13296_),
    .B(_13281_),
    .Y(_13369_));
 sky130_fd_sc_hd__clkbuf_4 _14817_ (.A(_13369_),
    .X(_13370_));
 sky130_fd_sc_hd__nor2_1 _14818_ (.A(_13286_),
    .B(_13288_),
    .Y(_13371_));
 sky130_fd_sc_hd__nor2_2 _14819_ (.A(_13371_),
    .B(_13300_),
    .Y(_13372_));
 sky130_fd_sc_hd__nand2_1 _14820_ (.A(_13314_),
    .B(_13291_),
    .Y(_13373_));
 sky130_fd_sc_hd__clkbuf_4 _14821_ (.A(_13373_),
    .X(_13374_));
 sky130_fd_sc_hd__nand2_1 _14822_ (.A(_13305_),
    .B(_13321_),
    .Y(_13375_));
 sky130_fd_sc_hd__nor2_1 _14823_ (.A(_13375_),
    .B(_13285_),
    .Y(_13376_));
 sky130_fd_sc_hd__or2_1 _14824_ (.A(_13288_),
    .B(_13306_),
    .X(_13377_));
 sky130_fd_sc_hd__buf_2 _14825_ (.A(_13377_),
    .X(_13378_));
 sky130_fd_sc_hd__nor2_1 _14826_ (.A(_13296_),
    .B(_13378_),
    .Y(_13379_));
 sky130_fd_sc_hd__or2_1 _14827_ (.A(_13286_),
    .B(_13288_),
    .X(_13380_));
 sky130_fd_sc_hd__nor2_2 _14828_ (.A(_13380_),
    .B(_13369_),
    .Y(_13381_));
 sky130_fd_sc_hd__o21a_1 _14829_ (.A1(_13379_),
    .A2(_13381_),
    .B1(_13331_),
    .X(_13382_));
 sky130_fd_sc_hd__nor2_1 _14830_ (.A(_13282_),
    .B(_13330_),
    .Y(_13383_));
 sky130_fd_sc_hd__or2_1 _14831_ (.A(_13382_),
    .B(_13383_),
    .X(_13384_));
 sky130_fd_sc_hd__clkbuf_4 _14832_ (.A(_13314_),
    .X(_13385_));
 sky130_fd_sc_hd__o21ai_1 _14833_ (.A1(_13376_),
    .A2(_13384_),
    .B1(_13385_),
    .Y(_13386_));
 sky130_fd_sc_hd__clkbuf_4 _14834_ (.A(_13287_),
    .X(_13387_));
 sky130_fd_sc_hd__or2_1 _14835_ (.A(\rvcpu.dp.pcreg.q[3] ),
    .B(_13280_),
    .X(_13388_));
 sky130_fd_sc_hd__buf_4 _14836_ (.A(_13388_),
    .X(_13389_));
 sky130_fd_sc_hd__nand2_4 _14837_ (.A(_13288_),
    .B(_13280_),
    .Y(_13390_));
 sky130_fd_sc_hd__nand2_4 _14838_ (.A(_13389_),
    .B(_13390_),
    .Y(_13391_));
 sky130_fd_sc_hd__nand2_2 _14839_ (.A(_13387_),
    .B(_13391_),
    .Y(_13392_));
 sky130_fd_sc_hd__nand2b_4 _14840_ (.A_N(_13281_),
    .B(_13288_),
    .Y(_13393_));
 sky130_fd_sc_hd__and3_1 _14841_ (.A(_13291_),
    .B(_13346_),
    .C(_13393_),
    .X(_13394_));
 sky130_fd_sc_hd__a2111o_1 _14842_ (.A1(_13332_),
    .A2(_13392_),
    .B1(_13394_),
    .C1(_13304_),
    .D1(_13314_),
    .X(_13395_));
 sky130_fd_sc_hd__o311a_1 _14843_ (.A1(_13370_),
    .A2(_13372_),
    .A3(_13374_),
    .B1(_13386_),
    .C1(_13395_),
    .X(_13396_));
 sky130_fd_sc_hd__buf_4 _14844_ (.A(_13296_),
    .X(_13397_));
 sky130_fd_sc_hd__nand2_4 _14845_ (.A(_13331_),
    .B(_13397_),
    .Y(_13398_));
 sky130_fd_sc_hd__nor2_2 _14846_ (.A(\rvcpu.dp.pcreg.q[3] ),
    .B(_13280_),
    .Y(_13399_));
 sky130_fd_sc_hd__and2_1 _14847_ (.A(\rvcpu.dp.pcreg.q[3] ),
    .B(\rvcpu.dp.pcreg.q[2] ),
    .X(_13400_));
 sky130_fd_sc_hd__buf_4 _14848_ (.A(_13400_),
    .X(_13401_));
 sky130_fd_sc_hd__nor2_4 _14849_ (.A(_13399_),
    .B(_13401_),
    .Y(_13402_));
 sky130_fd_sc_hd__nand2_4 _14850_ (.A(_13287_),
    .B(_13402_),
    .Y(_13403_));
 sky130_fd_sc_hd__o31a_1 _14851_ (.A1(_13398_),
    .A2(_13357_),
    .A3(_13403_),
    .B1(\rvcpu.dp.pcreg.q[9] ),
    .X(_13404_));
 sky130_fd_sc_hd__o21ai_1 _14852_ (.A1(_13368_),
    .A2(_13396_),
    .B1(_13404_),
    .Y(_13405_));
 sky130_fd_sc_hd__or2_1 _14853_ (.A(_13367_),
    .B(_13405_),
    .X(_13406_));
 sky130_fd_sc_hd__o31a_1 _14854_ (.A1(_13316_),
    .A2(_13325_),
    .A3(_13362_),
    .B1(_13406_),
    .X(net26));
 sky130_fd_sc_hd__nand2_1 _14855_ (.A(_13341_),
    .B(_13294_),
    .Y(_13407_));
 sky130_fd_sc_hd__and2_1 _14856_ (.A(_13312_),
    .B(_13313_),
    .X(_13408_));
 sky130_fd_sc_hd__clkbuf_4 _14857_ (.A(_13408_),
    .X(_13409_));
 sky130_fd_sc_hd__nand2_4 _14858_ (.A(_13291_),
    .B(_13409_),
    .Y(_13410_));
 sky130_fd_sc_hd__nor2_1 _14859_ (.A(_13407_),
    .B(_13410_),
    .Y(_13411_));
 sky130_fd_sc_hd__clkbuf_4 _14860_ (.A(\rvcpu.dp.pcreg.q[8] ),
    .X(_13412_));
 sky130_fd_sc_hd__nor2_2 _14861_ (.A(_13412_),
    .B(_13385_),
    .Y(_13413_));
 sky130_fd_sc_hd__nand2_8 _14862_ (.A(\rvcpu.dp.pcreg.q[4] ),
    .B(\rvcpu.dp.pcreg.q[3] ),
    .Y(_13414_));
 sky130_fd_sc_hd__nand2_2 _14863_ (.A(_13380_),
    .B(_13414_),
    .Y(_13415_));
 sky130_fd_sc_hd__nor2_2 _14864_ (.A(_13369_),
    .B(_13415_),
    .Y(_13416_));
 sky130_fd_sc_hd__or2_1 _14865_ (.A(_13332_),
    .B(_13416_),
    .X(_13417_));
 sky130_fd_sc_hd__or2b_1 _14866_ (.A(_13417_),
    .B_N(_13351_),
    .X(_13418_));
 sky130_fd_sc_hd__clkbuf_4 _14867_ (.A(_13371_),
    .X(_13419_));
 sky130_fd_sc_hd__nand2_4 _14868_ (.A(_13419_),
    .B(_13293_),
    .Y(_13420_));
 sky130_fd_sc_hd__nand2_1 _14869_ (.A(_13358_),
    .B(_13420_),
    .Y(_13421_));
 sky130_fd_sc_hd__or2_2 _14870_ (.A(_13313_),
    .B(_13331_),
    .X(_13422_));
 sky130_fd_sc_hd__clkbuf_4 _14871_ (.A(_13422_),
    .X(_13423_));
 sky130_fd_sc_hd__nor2_1 _14872_ (.A(_13281_),
    .B(_13414_),
    .Y(_13424_));
 sky130_fd_sc_hd__buf_4 _14873_ (.A(_13380_),
    .X(_13425_));
 sky130_fd_sc_hd__nor2_1 _14874_ (.A(_13425_),
    .B(_13336_),
    .Y(_13426_));
 sky130_fd_sc_hd__nor2_1 _14875_ (.A(_13424_),
    .B(_13426_),
    .Y(_13427_));
 sky130_fd_sc_hd__nor2_2 _14876_ (.A(_13313_),
    .B(_13283_),
    .Y(_13428_));
 sky130_fd_sc_hd__clkbuf_4 _14877_ (.A(_13428_),
    .X(_13429_));
 sky130_fd_sc_hd__clkbuf_4 _14878_ (.A(_13303_),
    .X(_13430_));
 sky130_fd_sc_hd__clkbuf_4 _14879_ (.A(_13430_),
    .X(_13431_));
 sky130_fd_sc_hd__nor2b_4 _14880_ (.A(\rvcpu.dp.pcreg.q[3] ),
    .B_N(_13280_),
    .Y(_13432_));
 sky130_fd_sc_hd__or2_1 _14881_ (.A(\rvcpu.dp.pcreg.q[5] ),
    .B(_13280_),
    .X(_13433_));
 sky130_fd_sc_hd__clkbuf_4 _14882_ (.A(_13433_),
    .X(_13434_));
 sky130_fd_sc_hd__nor2_2 _14883_ (.A(_13289_),
    .B(_13434_),
    .Y(_13435_));
 sky130_fd_sc_hd__a21o_1 _14884_ (.A1(_13431_),
    .A2(_13432_),
    .B1(_13435_),
    .X(_13436_));
 sky130_fd_sc_hd__a2bb2o_1 _14885_ (.A1_N(_13423_),
    .A2_N(_13427_),
    .B1(_13429_),
    .B2(_13436_),
    .X(_13437_));
 sky130_fd_sc_hd__clkbuf_4 _14886_ (.A(\rvcpu.dp.pcreg.q[8] ),
    .X(_13438_));
 sky130_fd_sc_hd__clkbuf_4 _14887_ (.A(_13438_),
    .X(_13439_));
 sky130_fd_sc_hd__a32o_1 _14888_ (.A1(_13413_),
    .A2(_13418_),
    .A3(_13421_),
    .B1(_13437_),
    .B2(_13439_),
    .X(_13440_));
 sky130_fd_sc_hd__o31a_1 _14889_ (.A1(_13325_),
    .A2(_13411_),
    .A3(_13440_),
    .B1(_13406_),
    .X(net25));
 sky130_fd_sc_hd__or2_2 _14890_ (.A(_13312_),
    .B(_13313_),
    .X(_13441_));
 sky130_fd_sc_hd__clkbuf_4 _14891_ (.A(_13441_),
    .X(_13442_));
 sky130_fd_sc_hd__or2_1 _14892_ (.A(_13337_),
    .B(_13435_),
    .X(_13443_));
 sky130_fd_sc_hd__nand2_1 _14893_ (.A(_13358_),
    .B(_13443_),
    .Y(_13444_));
 sky130_fd_sc_hd__nor2_1 _14894_ (.A(_13442_),
    .B(_13444_),
    .Y(_13445_));
 sky130_fd_sc_hd__and2b_1 _14895_ (.A_N(_13287_),
    .B(_13288_),
    .X(_13446_));
 sky130_fd_sc_hd__clkbuf_4 _14896_ (.A(_13446_),
    .X(_13447_));
 sky130_fd_sc_hd__nand2_1 _14897_ (.A(_13343_),
    .B(_13447_),
    .Y(_13448_));
 sky130_fd_sc_hd__and2_2 _14898_ (.A(_13397_),
    .B(_13387_),
    .X(_13449_));
 sky130_fd_sc_hd__nand2_1 _14899_ (.A(_13449_),
    .B(_13402_),
    .Y(_13450_));
 sky130_fd_sc_hd__nand2_4 _14900_ (.A(_13430_),
    .B(_13323_),
    .Y(_13451_));
 sky130_fd_sc_hd__a31o_1 _14901_ (.A1(_13448_),
    .A2(_13450_),
    .A3(_13451_),
    .B1(_13333_),
    .X(_13452_));
 sky130_fd_sc_hd__o21ai_1 _14902_ (.A1(_13378_),
    .A2(_13398_),
    .B1(_13452_),
    .Y(_13453_));
 sky130_fd_sc_hd__nor2_1 _14903_ (.A(_13287_),
    .B(_13390_),
    .Y(_13454_));
 sky130_fd_sc_hd__nand2_1 _14904_ (.A(_13317_),
    .B(_13454_),
    .Y(_13455_));
 sky130_fd_sc_hd__nor2_1 _14905_ (.A(_13315_),
    .B(_13455_),
    .Y(_13456_));
 sky130_fd_sc_hd__a211o_1 _14906_ (.A1(_13413_),
    .A2(_13453_),
    .B1(_13456_),
    .C1(_13325_),
    .X(_13457_));
 sky130_fd_sc_hd__o21a_1 _14907_ (.A1(_13445_),
    .A2(_13457_),
    .B1(_13406_),
    .X(net23));
 sky130_fd_sc_hd__nand2_4 _14908_ (.A(\rvcpu.dp.pcreg.q[8] ),
    .B(_13313_),
    .Y(_13458_));
 sky130_fd_sc_hd__nor2_1 _14909_ (.A(_13291_),
    .B(_13304_),
    .Y(_13459_));
 sky130_fd_sc_hd__a21o_1 _14910_ (.A1(_13321_),
    .A2(_13459_),
    .B1(_13337_),
    .X(_13460_));
 sky130_fd_sc_hd__a2bb2o_1 _14911_ (.A1_N(_13458_),
    .A2_N(_13360_),
    .B1(_13327_),
    .B2(_13460_),
    .X(_13461_));
 sky130_fd_sc_hd__nor2_1 _14912_ (.A(_13335_),
    .B(_13434_),
    .Y(_13462_));
 sky130_fd_sc_hd__clkbuf_4 _14913_ (.A(_13365_),
    .X(_13463_));
 sky130_fd_sc_hd__o21ai_1 _14914_ (.A1(_13379_),
    .A2(_13462_),
    .B1(_13463_),
    .Y(_13464_));
 sky130_fd_sc_hd__nor2_4 _14915_ (.A(_13425_),
    .B(_13434_),
    .Y(_13465_));
 sky130_fd_sc_hd__clkbuf_4 _14916_ (.A(_13412_),
    .X(_13466_));
 sky130_fd_sc_hd__nor2_1 _14917_ (.A(_13466_),
    .B(_13423_),
    .Y(_13467_));
 sky130_fd_sc_hd__a2bb2o_1 _14918_ (.A1_N(_13439_),
    .A2_N(_13464_),
    .B1(_13465_),
    .B2(_13467_),
    .X(_13468_));
 sky130_fd_sc_hd__o22a_1 _14919_ (.A1(_13457_),
    .A2(_13461_),
    .B1(_13468_),
    .B2(_13405_),
    .X(net22));
 sky130_fd_sc_hd__nand2_4 _14920_ (.A(\rvcpu.dp.pcreg.q[9] ),
    .B(_13368_),
    .Y(_13469_));
 sky130_fd_sc_hd__nor2_1 _14921_ (.A(_13341_),
    .B(_13336_),
    .Y(_13470_));
 sky130_fd_sc_hd__or2_1 _14922_ (.A(_13332_),
    .B(_13462_),
    .X(_13471_));
 sky130_fd_sc_hd__nand2_4 _14923_ (.A(_13303_),
    .B(_13414_),
    .Y(_13472_));
 sky130_fd_sc_hd__nor2_2 _14924_ (.A(_13402_),
    .B(_13472_),
    .Y(_13473_));
 sky130_fd_sc_hd__nand2_2 _14925_ (.A(_13333_),
    .B(_13364_),
    .Y(_13474_));
 sky130_fd_sc_hd__clkbuf_4 _14926_ (.A(_13314_),
    .X(_13475_));
 sky130_fd_sc_hd__o221a_1 _14927_ (.A1(_13470_),
    .A2(_13471_),
    .B1(_13473_),
    .B2(_13474_),
    .C1(_13475_),
    .X(_13476_));
 sky130_fd_sc_hd__nand2_1 _14928_ (.A(_13284_),
    .B(_13346_),
    .Y(_13477_));
 sky130_fd_sc_hd__or3_1 _14929_ (.A(_13432_),
    .B(_13422_),
    .C(_13477_),
    .X(_13478_));
 sky130_fd_sc_hd__or2_1 _14930_ (.A(_13322_),
    .B(_13478_),
    .X(_13479_));
 sky130_fd_sc_hd__or2_1 _14931_ (.A(_13329_),
    .B(_13422_),
    .X(_13480_));
 sky130_fd_sc_hd__nand2_1 _14932_ (.A(_13328_),
    .B(_13425_),
    .Y(_13481_));
 sky130_fd_sc_hd__or2_1 _14933_ (.A(_13313_),
    .B(_13283_),
    .X(_13482_));
 sky130_fd_sc_hd__clkbuf_4 _14934_ (.A(_13482_),
    .X(_13483_));
 sky130_fd_sc_hd__nand2_4 _14935_ (.A(_13284_),
    .B(_13287_),
    .Y(_13484_));
 sky130_fd_sc_hd__or3b_1 _14936_ (.A(_13481_),
    .B(_13483_),
    .C_N(_13484_),
    .X(_13485_));
 sky130_fd_sc_hd__and4b_1 _14937_ (.A_N(_13476_),
    .B(_13479_),
    .C(_13480_),
    .D(_13485_),
    .X(_13486_));
 sky130_fd_sc_hd__and2_1 _14938_ (.A(_13287_),
    .B(_13281_),
    .X(_13487_));
 sky130_fd_sc_hd__clkbuf_4 _14939_ (.A(_13487_),
    .X(_13488_));
 sky130_fd_sc_hd__nand2_4 _14940_ (.A(_13303_),
    .B(_13393_),
    .Y(_13489_));
 sky130_fd_sc_hd__nor2_1 _14941_ (.A(_13488_),
    .B(_13489_),
    .Y(_13490_));
 sky130_fd_sc_hd__o21ai_1 _14942_ (.A1(_13449_),
    .A2(_13490_),
    .B1(_13429_),
    .Y(_13491_));
 sky130_fd_sc_hd__or2_2 _14943_ (.A(_13295_),
    .B(_13432_),
    .X(_13492_));
 sky130_fd_sc_hd__nor2_1 _14944_ (.A(_13415_),
    .B(_13492_),
    .Y(_13493_));
 sky130_fd_sc_hd__nand2_1 _14945_ (.A(_13297_),
    .B(_13348_),
    .Y(_13494_));
 sky130_fd_sc_hd__nor2_1 _14946_ (.A(_13401_),
    .B(_13494_),
    .Y(_13495_));
 sky130_fd_sc_hd__clkbuf_4 _14947_ (.A(_13353_),
    .X(_13496_));
 sky130_fd_sc_hd__o21ai_1 _14948_ (.A1(_13493_),
    .A2(_13495_),
    .B1(_13496_),
    .Y(_13497_));
 sky130_fd_sc_hd__or3_1 _14949_ (.A(_13370_),
    .B(_13373_),
    .C(_13447_),
    .X(_13498_));
 sky130_fd_sc_hd__nand2_2 _14950_ (.A(\rvcpu.dp.pcreg.q[9] ),
    .B(_13438_),
    .Y(_13499_));
 sky130_fd_sc_hd__a41o_1 _14951_ (.A1(_13386_),
    .A2(_13491_),
    .A3(_13497_),
    .A4(_13498_),
    .B1(_13499_),
    .X(_13500_));
 sky130_fd_sc_hd__clkbuf_4 _14952_ (.A(_13357_),
    .X(_13501_));
 sky130_fd_sc_hd__a21o_1 _14953_ (.A1(_13330_),
    .A2(_13452_),
    .B1(_13501_),
    .X(_13502_));
 sky130_fd_sc_hd__nor2_1 _14954_ (.A(_13331_),
    .B(_13458_),
    .Y(_13503_));
 sky130_fd_sc_hd__clkbuf_4 _14955_ (.A(_13503_),
    .X(_13504_));
 sky130_fd_sc_hd__nor2_4 _14956_ (.A(_13284_),
    .B(_13300_),
    .Y(_13505_));
 sky130_fd_sc_hd__nor2_4 _14957_ (.A(_13287_),
    .B(_13281_),
    .Y(_13506_));
 sky130_fd_sc_hd__nor2_2 _14958_ (.A(_13296_),
    .B(_13506_),
    .Y(_13507_));
 sky130_fd_sc_hd__a22o_1 _14959_ (.A1(_13307_),
    .A2(_13505_),
    .B1(_13507_),
    .B2(_13402_),
    .X(_13508_));
 sky130_fd_sc_hd__clkbuf_4 _14960_ (.A(_13415_),
    .X(_13509_));
 sky130_fd_sc_hd__nand2_4 _14961_ (.A(_13397_),
    .B(_13307_),
    .Y(_13510_));
 sky130_fd_sc_hd__nor2_1 _14962_ (.A(_13509_),
    .B(_13510_),
    .Y(_13511_));
 sky130_fd_sc_hd__and3_1 _14963_ (.A(_13304_),
    .B(_13335_),
    .C(_13348_),
    .X(_13512_));
 sky130_fd_sc_hd__nand2_4 _14964_ (.A(\rvcpu.dp.pcreg.q[7] ),
    .B(\rvcpu.dp.pcreg.q[6] ),
    .Y(_13513_));
 sky130_fd_sc_hd__nor2_4 _14965_ (.A(_13311_),
    .B(_13513_),
    .Y(_13514_));
 sky130_fd_sc_hd__o21a_1 _14966_ (.A1(_13511_),
    .A2(_13512_),
    .B1(_13514_),
    .X(_13515_));
 sky130_fd_sc_hd__a211oi_1 _14967_ (.A1(_13504_),
    .A2(_13508_),
    .B1(_13515_),
    .C1(_13456_),
    .Y(_13516_));
 sky130_fd_sc_hd__clkbuf_4 _14968_ (.A(_13292_),
    .X(_13517_));
 sky130_fd_sc_hd__nand2_1 _14969_ (.A(_13517_),
    .B(_13337_),
    .Y(_13518_));
 sky130_fd_sc_hd__a211o_1 _14970_ (.A1(_13370_),
    .A2(_13472_),
    .B1(_13292_),
    .C1(_13419_),
    .X(_13519_));
 sky130_fd_sc_hd__a21o_1 _14971_ (.A1(_13518_),
    .A2(_13519_),
    .B1(_13442_),
    .X(_13520_));
 sky130_fd_sc_hd__clkbuf_4 _14972_ (.A(\rvcpu.dp.pcreg.q[9] ),
    .X(_13521_));
 sky130_fd_sc_hd__a31o_1 _14973_ (.A1(_13502_),
    .A2(_13516_),
    .A3(_13520_),
    .B1(_13521_),
    .X(_13522_));
 sky130_fd_sc_hd__o211ai_2 _14974_ (.A1(_13469_),
    .A2(_13486_),
    .B1(_13500_),
    .C1(_13522_),
    .Y(net21));
 sky130_fd_sc_hd__nor2_4 _14975_ (.A(\rvcpu.dp.pcreg.q[5] ),
    .B(_13322_),
    .Y(_13523_));
 sky130_fd_sc_hd__nand2_1 _14976_ (.A(_13335_),
    .B(_13523_),
    .Y(_13524_));
 sky130_fd_sc_hd__or2_1 _14977_ (.A(_13446_),
    .B(_13524_),
    .X(_13525_));
 sky130_fd_sc_hd__nand2_4 _14978_ (.A(_13287_),
    .B(_13281_),
    .Y(_13526_));
 sky130_fd_sc_hd__a311o_1 _14979_ (.A1(_13414_),
    .A2(_13526_),
    .A3(_13390_),
    .B1(_13483_),
    .C1(_13304_),
    .X(_13527_));
 sky130_fd_sc_hd__nor2_4 _14980_ (.A(_13335_),
    .B(_13369_),
    .Y(_13528_));
 sky130_fd_sc_hd__o21ai_1 _14981_ (.A1(_13528_),
    .A2(_13473_),
    .B1(_13463_),
    .Y(_13529_));
 sky130_fd_sc_hd__o211a_1 _14982_ (.A1(_13423_),
    .A2(_13525_),
    .B1(_13527_),
    .C1(_13529_),
    .X(_13530_));
 sky130_fd_sc_hd__nor2_2 _14983_ (.A(_13301_),
    .B(_13434_),
    .Y(_13531_));
 sky130_fd_sc_hd__a21oi_1 _14984_ (.A1(_13425_),
    .A2(_13531_),
    .B1(_13470_),
    .Y(_13532_));
 sky130_fd_sc_hd__clkbuf_4 _14985_ (.A(_13374_),
    .X(_13533_));
 sky130_fd_sc_hd__o22a_1 _14986_ (.A1(_13475_),
    .A2(_13360_),
    .B1(_13532_),
    .B2(_13533_),
    .X(_13534_));
 sky130_fd_sc_hd__a31oi_1 _14987_ (.A1(_13479_),
    .A2(_13530_),
    .A3(_13534_),
    .B1(_13439_),
    .Y(_13535_));
 sky130_fd_sc_hd__nor2_1 _14988_ (.A(_13393_),
    .B(_13484_),
    .Y(_13536_));
 sky130_fd_sc_hd__o21a_1 _14989_ (.A1(_13528_),
    .A2(_13536_),
    .B1(_13503_),
    .X(_13537_));
 sky130_fd_sc_hd__inv_2 _14990_ (.A(\rvcpu.dp.pcreg.q[9] ),
    .Y(_13538_));
 sky130_fd_sc_hd__clkbuf_4 _14991_ (.A(_13538_),
    .X(_13539_));
 sky130_fd_sc_hd__a211o_1 _14992_ (.A1(_13384_),
    .A2(_13319_),
    .B1(_13537_),
    .C1(_13539_),
    .X(_13540_));
 sky130_fd_sc_hd__nor2_2 _14993_ (.A(_13397_),
    .B(_13371_),
    .Y(_13541_));
 sky130_fd_sc_hd__clkbuf_4 _14994_ (.A(_13358_),
    .X(_13542_));
 sky130_fd_sc_hd__a211o_1 _14995_ (.A1(_13414_),
    .A2(_13541_),
    .B1(_13523_),
    .C1(_13542_),
    .X(_13543_));
 sky130_fd_sc_hd__o211a_1 _14996_ (.A1(_13474_),
    .A2(_13490_),
    .B1(_13543_),
    .C1(_13327_),
    .X(_13544_));
 sky130_fd_sc_hd__nand2_1 _14997_ (.A(_13303_),
    .B(_13322_),
    .Y(_13545_));
 sky130_fd_sc_hd__nor2_4 _14998_ (.A(_13287_),
    .B(_13391_),
    .Y(_13546_));
 sky130_fd_sc_hd__o31a_1 _14999_ (.A1(_13303_),
    .A2(_13321_),
    .A3(_13546_),
    .B1(_13331_),
    .X(_13547_));
 sky130_fd_sc_hd__or2_1 _15000_ (.A(_13391_),
    .B(_13484_),
    .X(_13548_));
 sky130_fd_sc_hd__and3_1 _15001_ (.A(_13545_),
    .B(_13547_),
    .C(_13548_),
    .X(_13549_));
 sky130_fd_sc_hd__nor2_1 _15002_ (.A(_13320_),
    .B(_13510_),
    .Y(_13550_));
 sky130_fd_sc_hd__a21o_1 _15003_ (.A1(_13509_),
    .A2(_13507_),
    .B1(_13550_),
    .X(_13551_));
 sky130_fd_sc_hd__inv_2 _15004_ (.A(_13364_),
    .Y(_13552_));
 sky130_fd_sc_hd__nor2_2 _15005_ (.A(_13341_),
    .B(_13492_),
    .Y(_13553_));
 sky130_fd_sc_hd__o21a_1 _15006_ (.A1(_13552_),
    .A2(_13553_),
    .B1(_13514_),
    .X(_13554_));
 sky130_fd_sc_hd__a311o_1 _15007_ (.A1(_13333_),
    .A2(_13326_),
    .A3(_13337_),
    .B1(_13554_),
    .C1(\rvcpu.dp.pcreg.q[9] ),
    .X(_13555_));
 sky130_fd_sc_hd__a21oi_1 _15008_ (.A1(_13344_),
    .A2(_13420_),
    .B1(_13410_),
    .Y(_13556_));
 sky130_fd_sc_hd__a211o_1 _15009_ (.A1(_13504_),
    .A2(_13551_),
    .B1(_13555_),
    .C1(_13556_),
    .X(_13557_));
 sky130_fd_sc_hd__or2_1 _15010_ (.A(_13305_),
    .B(_13346_),
    .X(_13558_));
 sky130_fd_sc_hd__buf_2 _15011_ (.A(_13558_),
    .X(_13559_));
 sky130_fd_sc_hd__nand2_1 _15012_ (.A(_13305_),
    .B(_13323_),
    .Y(_13560_));
 sky130_fd_sc_hd__and2_2 _15013_ (.A(_13303_),
    .B(_13560_),
    .X(_13561_));
 sky130_fd_sc_hd__nor2_2 _15014_ (.A(\rvcpu.dp.pcreg.q[5] ),
    .B(_13281_),
    .Y(_13562_));
 sky130_fd_sc_hd__a21oi_1 _15015_ (.A1(_13559_),
    .A2(_13561_),
    .B1(_13562_),
    .Y(_13563_));
 sky130_fd_sc_hd__or2_1 _15016_ (.A(_13333_),
    .B(_13563_),
    .X(_13564_));
 sky130_fd_sc_hd__nand2_2 _15017_ (.A(_13397_),
    .B(_13390_),
    .Y(_13565_));
 sky130_fd_sc_hd__o21ai_1 _15018_ (.A1(_13387_),
    .A2(_13565_),
    .B1(_13542_),
    .Y(_13566_));
 sky130_fd_sc_hd__a21o_1 _15019_ (.A1(_13403_),
    .A2(_13523_),
    .B1(_13561_),
    .X(_13567_));
 sky130_fd_sc_hd__a31o_1 _15020_ (.A1(_13333_),
    .A2(_13420_),
    .A3(_13525_),
    .B1(_13357_),
    .X(_13568_));
 sky130_fd_sc_hd__a21oi_1 _15021_ (.A1(_13517_),
    .A2(_13567_),
    .B1(_13568_),
    .Y(_13569_));
 sky130_fd_sc_hd__a31o_1 _15022_ (.A1(_13327_),
    .A2(_13564_),
    .A3(_13566_),
    .B1(_13569_),
    .X(_13570_));
 sky130_fd_sc_hd__a211o_1 _15023_ (.A1(_13409_),
    .A2(_13549_),
    .B1(_13557_),
    .C1(_13570_),
    .X(_13571_));
 sky130_fd_sc_hd__o31a_1 _15024_ (.A1(_13535_),
    .A2(_13540_),
    .A3(_13544_),
    .B1(_13571_),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_4 _15025_ (.A(_13521_),
    .X(_13572_));
 sky130_fd_sc_hd__clkbuf_4 _15026_ (.A(_13513_),
    .X(_13573_));
 sky130_fd_sc_hd__nand2_1 _15027_ (.A(_13397_),
    .B(_13414_),
    .Y(_13574_));
 sky130_fd_sc_hd__or2_1 _15028_ (.A(_13574_),
    .B(_13546_),
    .X(_13575_));
 sky130_fd_sc_hd__and2b_1 _15029_ (.A_N(_13553_),
    .B(_13575_),
    .X(_13576_));
 sky130_fd_sc_hd__or2_1 _15030_ (.A(_13322_),
    .B(_13492_),
    .X(_13577_));
 sky130_fd_sc_hd__nor2_1 _15031_ (.A(_13424_),
    .B(_13577_),
    .Y(_13578_));
 sky130_fd_sc_hd__nor2_1 _15032_ (.A(_13343_),
    .B(_13578_),
    .Y(_13579_));
 sky130_fd_sc_hd__o221a_1 _15033_ (.A1(_13573_),
    .A2(_13576_),
    .B1(_13579_),
    .B2(_13423_),
    .C1(_13466_),
    .X(_13580_));
 sky130_fd_sc_hd__clkbuf_4 _15034_ (.A(_13483_),
    .X(_13581_));
 sky130_fd_sc_hd__o21ba_1 _15035_ (.A1(_13324_),
    .A2(_13489_),
    .B1_N(_13381_),
    .X(_13582_));
 sky130_fd_sc_hd__a21oi_1 _15036_ (.A1(_13559_),
    .A2(_13561_),
    .B1(_13550_),
    .Y(_13583_));
 sky130_fd_sc_hd__o22a_1 _15037_ (.A1(_13581_),
    .A2(_13582_),
    .B1(_13583_),
    .B2(_13533_),
    .X(_13584_));
 sky130_fd_sc_hd__or3_1 _15038_ (.A(_13332_),
    .B(_13562_),
    .C(_13427_),
    .X(_13585_));
 sky130_fd_sc_hd__nor2_1 _15039_ (.A(_13282_),
    .B(_13415_),
    .Y(_13586_));
 sky130_fd_sc_hd__or3_1 _15040_ (.A(_13398_),
    .B(_13322_),
    .C(_13586_),
    .X(_13587_));
 sky130_fd_sc_hd__a31o_1 _15041_ (.A1(_13338_),
    .A2(_13585_),
    .A3(_13587_),
    .B1(_13385_),
    .X(_13588_));
 sky130_fd_sc_hd__nor2_2 _15042_ (.A(_13387_),
    .B(_13402_),
    .Y(_13589_));
 sky130_fd_sc_hd__a21oi_2 _15043_ (.A1(_13336_),
    .A2(_13472_),
    .B1(_13589_),
    .Y(_13590_));
 sky130_fd_sc_hd__or4_1 _15044_ (.A(_13374_),
    .B(_13416_),
    .C(_13465_),
    .D(_13590_),
    .X(_13591_));
 sky130_fd_sc_hd__nand2_1 _15045_ (.A(_13282_),
    .B(_13415_),
    .Y(_13592_));
 sky130_fd_sc_hd__and2_1 _15046_ (.A(_13297_),
    .B(_13592_),
    .X(_13593_));
 sky130_fd_sc_hd__a21oi_1 _15047_ (.A1(_13353_),
    .A2(_13593_),
    .B1(_13438_),
    .Y(_13594_));
 sky130_fd_sc_hd__and3_1 _15048_ (.A(_13588_),
    .B(_13591_),
    .C(_13594_),
    .X(_13595_));
 sky130_fd_sc_hd__a21oi_1 _15049_ (.A1(_13580_),
    .A2(_13584_),
    .B1(_13595_),
    .Y(_13596_));
 sky130_fd_sc_hd__nand2_1 _15050_ (.A(_13333_),
    .B(_13370_),
    .Y(_13597_));
 sky130_fd_sc_hd__nand2_2 _15051_ (.A(_13297_),
    .B(_13526_),
    .Y(_13598_));
 sky130_fd_sc_hd__clkbuf_4 _15052_ (.A(_13358_),
    .X(_13599_));
 sky130_fd_sc_hd__nor2_1 _15053_ (.A(_13599_),
    .B(_13473_),
    .Y(_13600_));
 sky130_fd_sc_hd__o21ai_1 _15054_ (.A1(_13598_),
    .A2(_13546_),
    .B1(_13600_),
    .Y(_13601_));
 sky130_fd_sc_hd__o311a_1 _15055_ (.A1(_13449_),
    .A2(_13490_),
    .A3(_13597_),
    .B1(_13601_),
    .C1(_13327_),
    .X(_13602_));
 sky130_fd_sc_hd__nand2_1 _15056_ (.A(_13291_),
    .B(_13578_),
    .Y(_13603_));
 sky130_fd_sc_hd__nand2_2 _15057_ (.A(_13328_),
    .B(_13447_),
    .Y(_13604_));
 sky130_fd_sc_hd__o21a_1 _15058_ (.A1(_13292_),
    .A2(_13604_),
    .B1(_13329_),
    .X(_13605_));
 sky130_fd_sc_hd__a21oi_1 _15059_ (.A1(_13603_),
    .A2(_13605_),
    .B1(_13501_),
    .Y(_13606_));
 sky130_fd_sc_hd__and3_2 _15060_ (.A(_13397_),
    .B(_13387_),
    .C(_13390_),
    .X(_13607_));
 sky130_fd_sc_hd__nor2_2 _15061_ (.A(\rvcpu.dp.pcreg.q[8] ),
    .B(_13513_),
    .Y(_13608_));
 sky130_fd_sc_hd__o21a_1 _15062_ (.A1(_13607_),
    .A2(_13473_),
    .B1(_13608_),
    .X(_13609_));
 sky130_fd_sc_hd__nand2_1 _15063_ (.A(_13335_),
    .B(_13294_),
    .Y(_13610_));
 sky130_fd_sc_hd__a21oi_1 _15064_ (.A1(_13364_),
    .A2(_13610_),
    .B1(_13410_),
    .Y(_13611_));
 sky130_fd_sc_hd__or4_1 _15065_ (.A(_13540_),
    .B(_13606_),
    .C(_13609_),
    .D(_13611_),
    .X(_13612_));
 sky130_fd_sc_hd__o22a_1 _15066_ (.A1(_13572_),
    .A2(_13596_),
    .B1(_13602_),
    .B2(_13612_),
    .X(net19));
 sky130_fd_sc_hd__nor2_1 _15067_ (.A(_13284_),
    .B(_13372_),
    .Y(_13613_));
 sky130_fd_sc_hd__or3_1 _15068_ (.A(_13331_),
    .B(_13562_),
    .C(_13613_),
    .X(_13614_));
 sky130_fd_sc_hd__or2_1 _15069_ (.A(_13397_),
    .B(_13282_),
    .X(_13615_));
 sky130_fd_sc_hd__nor2_1 _15070_ (.A(_13615_),
    .B(_13447_),
    .Y(_13616_));
 sky130_fd_sc_hd__or3_1 _15071_ (.A(_13470_),
    .B(_13614_),
    .C(_13616_),
    .X(_13617_));
 sky130_fd_sc_hd__a21oi_1 _15072_ (.A1(_13338_),
    .A2(_13617_),
    .B1(_13501_),
    .Y(_13618_));
 sky130_fd_sc_hd__a21o_1 _15073_ (.A1(_13289_),
    .A2(_13507_),
    .B1(_13511_),
    .X(_13619_));
 sky130_fd_sc_hd__a211o_1 _15074_ (.A1(_13504_),
    .A2(_13619_),
    .B1(_13515_),
    .C1(_13521_),
    .X(_13620_));
 sky130_fd_sc_hd__a21o_1 _15075_ (.A1(_13301_),
    .A2(_13562_),
    .B1(_13359_),
    .X(_13621_));
 sky130_fd_sc_hd__nor2_1 _15076_ (.A(_13509_),
    .B(_13489_),
    .Y(_13622_));
 sky130_fd_sc_hd__a22o_1 _15077_ (.A1(_13496_),
    .A2(_13621_),
    .B1(_13622_),
    .B2(_13429_),
    .X(_13623_));
 sky130_fd_sc_hd__a2bb2o_1 _15078_ (.A1_N(_13410_),
    .A2_N(_13420_),
    .B1(_13623_),
    .B2(_13466_),
    .X(_13624_));
 sky130_fd_sc_hd__a21boi_1 _15079_ (.A1(_13450_),
    .A2(_13489_),
    .B1_N(_13484_),
    .Y(_13625_));
 sky130_fd_sc_hd__or4_1 _15080_ (.A(_13358_),
    .B(_13607_),
    .C(_13465_),
    .D(_13493_),
    .X(_13626_));
 sky130_fd_sc_hd__o211a_1 _15081_ (.A1(_13517_),
    .A2(_13625_),
    .B1(_13626_),
    .C1(_13326_),
    .X(_13627_));
 sky130_fd_sc_hd__nor2_2 _15082_ (.A(_13320_),
    .B(_13346_),
    .Y(_13628_));
 sky130_fd_sc_hd__o21a_1 _15083_ (.A1(_13628_),
    .A2(_13359_),
    .B1(_13608_),
    .X(_13629_));
 sky130_fd_sc_hd__nand2_1 _15084_ (.A(_13282_),
    .B(_13317_),
    .Y(_13630_));
 sky130_fd_sc_hd__nor2_1 _15085_ (.A(_13447_),
    .B(_13630_),
    .Y(_13631_));
 sky130_fd_sc_hd__o31a_1 _15086_ (.A1(_13376_),
    .A2(_13383_),
    .A3(_13631_),
    .B1(_13319_),
    .X(_13632_));
 sky130_fd_sc_hd__or4_1 _15087_ (.A(_13538_),
    .B(_13611_),
    .C(_13629_),
    .D(_13632_),
    .X(_13633_));
 sky130_fd_sc_hd__nor2_2 _15088_ (.A(_13389_),
    .B(_13484_),
    .Y(_13634_));
 sky130_fd_sc_hd__nand2_1 _15089_ (.A(_13428_),
    .B(_13634_),
    .Y(_13635_));
 sky130_fd_sc_hd__a41o_1 _15090_ (.A1(_13478_),
    .A2(_13480_),
    .A3(_13527_),
    .A4(_13635_),
    .B1(_13438_),
    .X(_13636_));
 sky130_fd_sc_hd__or3b_1 _15091_ (.A(_13627_),
    .B(_13633_),
    .C_N(_13636_),
    .X(_13637_));
 sky130_fd_sc_hd__o31a_1 _15092_ (.A1(_13618_),
    .A2(_13620_),
    .A3(_13624_),
    .B1(_13637_),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_4 _15093_ (.A(_13521_),
    .X(_13638_));
 sky130_fd_sc_hd__nor2_2 _15094_ (.A(_13401_),
    .B(_13484_),
    .Y(_13639_));
 sky130_fd_sc_hd__and2_1 _15095_ (.A(_13304_),
    .B(_13589_),
    .X(_13640_));
 sky130_fd_sc_hd__a211o_1 _15096_ (.A1(_13403_),
    .A2(_13523_),
    .B1(_13639_),
    .C1(_13640_),
    .X(_13641_));
 sky130_fd_sc_hd__or2_1 _15097_ (.A(_13454_),
    .B(_13477_),
    .X(_13642_));
 sky130_fd_sc_hd__or2_1 _15098_ (.A(_13399_),
    .B(_13642_),
    .X(_13643_));
 sky130_fd_sc_hd__nand2_1 _15099_ (.A(_13524_),
    .B(_13643_),
    .Y(_13644_));
 sky130_fd_sc_hd__a21o_1 _15100_ (.A1(_13393_),
    .A2(_13523_),
    .B1(_13470_),
    .X(_13645_));
 sky130_fd_sc_hd__and2_2 _15101_ (.A(_13314_),
    .B(_13292_),
    .X(_13646_));
 sky130_fd_sc_hd__a221o_1 _15102_ (.A1(_13353_),
    .A2(_13644_),
    .B1(_13645_),
    .B2(_13646_),
    .C1(_13412_),
    .X(_13647_));
 sky130_fd_sc_hd__nor2_1 _15103_ (.A(_13488_),
    .B(_13492_),
    .Y(_13648_));
 sky130_fd_sc_hd__nand2_2 _15104_ (.A(_13297_),
    .B(_13560_),
    .Y(_13649_));
 sky130_fd_sc_hd__nor2_1 _15105_ (.A(_13324_),
    .B(_13649_),
    .Y(_13650_));
 sky130_fd_sc_hd__o21a_1 _15106_ (.A1(_13648_),
    .A2(_13650_),
    .B1(_13429_),
    .X(_13651_));
 sky130_fd_sc_hd__a211o_1 _15107_ (.A1(_13463_),
    .A2(_13641_),
    .B1(_13647_),
    .C1(_13651_),
    .X(_13652_));
 sky130_fd_sc_hd__a21o_1 _15108_ (.A1(_13392_),
    .A2(_13523_),
    .B1(_13536_),
    .X(_13653_));
 sky130_fd_sc_hd__and3_1 _15109_ (.A(_13387_),
    .B(_13389_),
    .C(_13390_),
    .X(_13654_));
 sky130_fd_sc_hd__a31o_1 _15110_ (.A1(_13298_),
    .A2(_13463_),
    .A3(_13654_),
    .B1(_13368_),
    .X(_13655_));
 sky130_fd_sc_hd__nor2_1 _15111_ (.A(_13303_),
    .B(_13432_),
    .Y(_13656_));
 sky130_fd_sc_hd__and2_1 _15112_ (.A(_13348_),
    .B(_13656_),
    .X(_13657_));
 sky130_fd_sc_hd__and2b_1 _15113_ (.A_N(_13282_),
    .B(_13305_),
    .X(_13658_));
 sky130_fd_sc_hd__nor2_2 _15114_ (.A(_13658_),
    .B(_13484_),
    .Y(_13659_));
 sky130_fd_sc_hd__o21a_1 _15115_ (.A1(_13657_),
    .A2(_13659_),
    .B1(_13353_),
    .X(_13660_));
 sky130_fd_sc_hd__a41o_1 _15116_ (.A1(_13307_),
    .A2(_13393_),
    .A3(_13598_),
    .A4(_13429_),
    .B1(_13660_),
    .X(_13661_));
 sky130_fd_sc_hd__a211o_1 _15117_ (.A1(_13646_),
    .A2(_13653_),
    .B1(_13655_),
    .C1(_13661_),
    .X(_13662_));
 sky130_fd_sc_hd__nor2_1 _15118_ (.A(_13417_),
    .B(_13590_),
    .Y(_13663_));
 sky130_fd_sc_hd__o31a_1 _15119_ (.A1(_13412_),
    .A2(_13549_),
    .A3(_13663_),
    .B1(_13357_),
    .X(_13664_));
 sky130_fd_sc_hd__clkbuf_4 _15120_ (.A(_13320_),
    .X(_13665_));
 sky130_fd_sc_hd__nand2_1 _15121_ (.A(_13665_),
    .B(_13294_),
    .Y(_13666_));
 sky130_fd_sc_hd__and4_1 _15122_ (.A(_13425_),
    .B(_13428_),
    .C(_13494_),
    .D(_13666_),
    .X(_13667_));
 sky130_fd_sc_hd__nand2_2 _15123_ (.A(_13298_),
    .B(_13349_),
    .Y(_13668_));
 sky130_fd_sc_hd__a211o_1 _15124_ (.A1(_13668_),
    .A2(_13451_),
    .B1(_13423_),
    .C1(_13324_),
    .X(_13669_));
 sky130_fd_sc_hd__or3b_1 _15125_ (.A(_13664_),
    .B(_13667_),
    .C_N(_13669_),
    .X(_13670_));
 sky130_fd_sc_hd__nor2_2 _15126_ (.A(_13296_),
    .B(_13347_),
    .Y(_13671_));
 sky130_fd_sc_hd__nand2_2 _15127_ (.A(\rvcpu.dp.pcreg.q[6] ),
    .B(_13389_),
    .Y(_13672_));
 sky130_fd_sc_hd__or3_1 _15128_ (.A(_13671_),
    .B(_13562_),
    .C(_13672_),
    .X(_13673_));
 sky130_fd_sc_hd__and3_1 _15129_ (.A(_13346_),
    .B(_13389_),
    .C(_13317_),
    .X(_13674_));
 sky130_fd_sc_hd__inv_2 _15130_ (.A(_13674_),
    .Y(_13675_));
 sky130_fd_sc_hd__a41o_1 _15131_ (.A1(_13330_),
    .A2(_13603_),
    .A3(_13673_),
    .A4(_13675_),
    .B1(_13475_),
    .X(_13676_));
 sky130_fd_sc_hd__o22a_1 _15132_ (.A1(_13372_),
    .A2(_13336_),
    .B1(_13510_),
    .B2(_13401_),
    .X(_13677_));
 sky130_fd_sc_hd__nor2_1 _15133_ (.A(_13607_),
    .B(_13553_),
    .Y(_13678_));
 sky130_fd_sc_hd__o221a_1 _15134_ (.A1(_13533_),
    .A2(_13677_),
    .B1(_13678_),
    .B2(_13573_),
    .C1(_13438_),
    .X(_13679_));
 sky130_fd_sc_hd__a21oi_1 _15135_ (.A1(_13676_),
    .A2(_13679_),
    .B1(_13638_),
    .Y(_13680_));
 sky130_fd_sc_hd__a32o_1 _15136_ (.A1(_13638_),
    .A2(_13652_),
    .A3(_13662_),
    .B1(_13670_),
    .B2(_13680_),
    .X(net17));
 sky130_fd_sc_hd__inv_2 _15137_ (.A(_13546_),
    .Y(_13681_));
 sky130_fd_sc_hd__clkbuf_4 _15138_ (.A(_13304_),
    .X(_13682_));
 sky130_fd_sc_hd__a311o_1 _15139_ (.A1(_13335_),
    .A2(_13526_),
    .A3(_13681_),
    .B1(_13573_),
    .C1(_13682_),
    .X(_13683_));
 sky130_fd_sc_hd__or3_1 _15140_ (.A(_13573_),
    .B(_13472_),
    .C(_13546_),
    .X(_13684_));
 sky130_fd_sc_hd__nor2_1 _15141_ (.A(_13328_),
    .B(_13289_),
    .Y(_13685_));
 sky130_fd_sc_hd__o41a_1 _15142_ (.A1(_13488_),
    .A2(_13685_),
    .A3(_13581_),
    .A4(_13492_),
    .B1(_13527_),
    .X(_13686_));
 sky130_fd_sc_hd__a21o_1 _15143_ (.A1(_13524_),
    .A2(_13642_),
    .B1(_13423_),
    .X(_13687_));
 sky130_fd_sc_hd__a41o_1 _15144_ (.A1(_13683_),
    .A2(_13684_),
    .A3(_13686_),
    .A4(_13687_),
    .B1(_13439_),
    .X(_13688_));
 sky130_fd_sc_hd__nor2_2 _15145_ (.A(_13430_),
    .B(_13447_),
    .Y(_13689_));
 sky130_fd_sc_hd__and2_1 _15146_ (.A(_13403_),
    .B(_13507_),
    .X(_13690_));
 sky130_fd_sc_hd__a21oi_1 _15147_ (.A1(_13375_),
    .A2(_13689_),
    .B1(_13690_),
    .Y(_13691_));
 sky130_fd_sc_hd__nand2_1 _15148_ (.A(_13297_),
    .B(_13419_),
    .Y(_13692_));
 sky130_fd_sc_hd__nand2_1 _15149_ (.A(_13297_),
    .B(_13506_),
    .Y(_13693_));
 sky130_fd_sc_hd__nand2_1 _15150_ (.A(_13291_),
    .B(_13319_),
    .Y(_13694_));
 sky130_fd_sc_hd__a31o_1 _15151_ (.A1(_13692_),
    .A2(_13403_),
    .A3(_13693_),
    .B1(_13694_),
    .X(_13695_));
 sky130_fd_sc_hd__nor2_1 _15152_ (.A(_13447_),
    .B(_13434_),
    .Y(_13696_));
 sky130_fd_sc_hd__nand2_1 _15153_ (.A(_13333_),
    .B(_13344_),
    .Y(_13697_));
 sky130_fd_sc_hd__nor2_1 _15154_ (.A(_13506_),
    .B(_13472_),
    .Y(_13698_));
 sky130_fd_sc_hd__o32a_1 _15155_ (.A1(_13599_),
    .A2(_13659_),
    .A3(_13696_),
    .B1(_13697_),
    .B2(_13698_),
    .X(_13699_));
 sky130_fd_sc_hd__nand2_1 _15156_ (.A(_13327_),
    .B(_13699_),
    .Y(_13700_));
 sky130_fd_sc_hd__o211a_1 _15157_ (.A1(_13410_),
    .A2(_13691_),
    .B1(_13695_),
    .C1(_13700_),
    .X(_13701_));
 sky130_fd_sc_hd__o311a_1 _15158_ (.A1(_13328_),
    .A2(_13330_),
    .A3(_13458_),
    .B1(_13701_),
    .C1(_13572_),
    .X(_13702_));
 sky130_fd_sc_hd__or2_2 _15159_ (.A(_13305_),
    .B(_13526_),
    .X(_13703_));
 sky130_fd_sc_hd__nor2_1 _15160_ (.A(_13475_),
    .B(_13290_),
    .Y(_13704_));
 sky130_fd_sc_hd__a311o_1 _15161_ (.A1(_13429_),
    .A2(_13703_),
    .A3(_13541_),
    .B1(_13664_),
    .C1(_13704_),
    .X(_13705_));
 sky130_fd_sc_hd__clkbuf_4 _15162_ (.A(_13475_),
    .X(_13706_));
 sky130_fd_sc_hd__o21ai_1 _15163_ (.A1(_13419_),
    .A2(_13603_),
    .B1(_13673_),
    .Y(_13707_));
 sky130_fd_sc_hd__nor2_1 _15164_ (.A(_13674_),
    .B(_13707_),
    .Y(_13708_));
 sky130_fd_sc_hd__o2bb2a_1 _15165_ (.A1_N(_13509_),
    .A2_N(_13507_),
    .B1(_13565_),
    .B2(_13506_),
    .X(_13709_));
 sky130_fd_sc_hd__o21a_1 _15166_ (.A1(_13308_),
    .A2(_13565_),
    .B1(_13577_),
    .X(_13710_));
 sky130_fd_sc_hd__o221a_1 _15167_ (.A1(_13533_),
    .A2(_13709_),
    .B1(_13710_),
    .B2(_13573_),
    .C1(_13466_),
    .X(_13711_));
 sky130_fd_sc_hd__o21ai_1 _15168_ (.A1(_13706_),
    .A2(_13708_),
    .B1(_13711_),
    .Y(_13712_));
 sky130_fd_sc_hd__a21oi_1 _15169_ (.A1(_13705_),
    .A2(_13712_),
    .B1(_13572_),
    .Y(_13713_));
 sky130_fd_sc_hd__a21oi_4 _15170_ (.A1(_13688_),
    .A2(_13702_),
    .B1(_13713_),
    .Y(net16));
 sky130_fd_sc_hd__a21o_1 _15171_ (.A1(_13307_),
    .A2(_13317_),
    .B1(_13707_),
    .X(_13714_));
 sky130_fd_sc_hd__a21o_1 _15172_ (.A1(_13509_),
    .A2(_13294_),
    .B1(_13607_),
    .X(_13715_));
 sky130_fd_sc_hd__a22o_1 _15173_ (.A1(_13326_),
    .A2(_13714_),
    .B1(_13715_),
    .B2(_13504_),
    .X(_13716_));
 sky130_fd_sc_hd__nand2_2 _15174_ (.A(_13320_),
    .B(_13349_),
    .Y(_13717_));
 sky130_fd_sc_hd__o21a_1 _15175_ (.A1(_13320_),
    .A2(_13349_),
    .B1(_13430_),
    .X(_13718_));
 sky130_fd_sc_hd__a211o_1 _15176_ (.A1(_13717_),
    .A2(_13718_),
    .B1(_13374_),
    .C1(_13416_),
    .X(_13719_));
 sky130_fd_sc_hd__a211o_1 _15177_ (.A1(_13346_),
    .A2(_13391_),
    .B1(_13483_),
    .C1(_13298_),
    .X(_13720_));
 sky130_fd_sc_hd__nor2_2 _15178_ (.A(_13397_),
    .B(_13341_),
    .Y(_13721_));
 sky130_fd_sc_hd__o32a_1 _15179_ (.A1(_13401_),
    .A2(_13323_),
    .A3(_13721_),
    .B1(_13492_),
    .B2(_13321_),
    .X(_13722_));
 sky130_fd_sc_hd__or2_1 _15180_ (.A(_13513_),
    .B(_13722_),
    .X(_13723_));
 sky130_fd_sc_hd__a31o_1 _15181_ (.A1(_13719_),
    .A2(_13720_),
    .A3(_13723_),
    .B1(_13412_),
    .X(_13724_));
 sky130_fd_sc_hd__or3b_1 _15182_ (.A(_13554_),
    .B(_13716_),
    .C_N(_13724_),
    .X(_13725_));
 sky130_fd_sc_hd__o2111a_1 _15183_ (.A1(_13431_),
    .A2(_13289_),
    .B1(_13403_),
    .C1(_13307_),
    .D1(_13646_),
    .X(_13726_));
 sky130_fd_sc_hd__o221a_1 _15184_ (.A1(_13324_),
    .A2(_13489_),
    .B1(_13589_),
    .B2(_13431_),
    .C1(_13429_),
    .X(_13727_));
 sky130_fd_sc_hd__nand2_1 _15185_ (.A(_13320_),
    .B(_13523_),
    .Y(_13728_));
 sky130_fd_sc_hd__nand2_1 _15186_ (.A(_13451_),
    .B(_13728_),
    .Y(_13729_));
 sky130_fd_sc_hd__a31o_1 _15187_ (.A1(_13389_),
    .A2(_13353_),
    .A3(_13729_),
    .B1(_13412_),
    .X(_13730_));
 sky130_fd_sc_hd__o31a_1 _15188_ (.A1(_13465_),
    .A2(_13639_),
    .A3(_13640_),
    .B1(_13463_),
    .X(_13731_));
 sky130_fd_sc_hd__or4_1 _15189_ (.A(_13726_),
    .B(_13727_),
    .C(_13730_),
    .D(_13731_),
    .X(_13732_));
 sky130_fd_sc_hd__a21oi_1 _15190_ (.A1(_13344_),
    .A2(_13548_),
    .B1(_13533_),
    .Y(_13733_));
 sky130_fd_sc_hd__a21oi_1 _15191_ (.A1(_13336_),
    .A2(_13703_),
    .B1(_13581_),
    .Y(_13734_));
 sky130_fd_sc_hd__a21oi_1 _15192_ (.A1(_13392_),
    .A2(_13434_),
    .B1(_13423_),
    .Y(_13735_));
 sky130_fd_sc_hd__o41a_1 _15193_ (.A1(_13655_),
    .A2(_13733_),
    .A3(_13734_),
    .A4(_13735_),
    .B1(_13638_),
    .X(_13736_));
 sky130_fd_sc_hd__a22o_1 _15194_ (.A1(_13539_),
    .A2(_13725_),
    .B1(_13732_),
    .B2(_13736_),
    .X(net15));
 sky130_fd_sc_hd__or2_2 _15195_ (.A(_13282_),
    .B(_13415_),
    .X(_13737_));
 sky130_fd_sc_hd__o31a_1 _15196_ (.A1(_13301_),
    .A2(_13488_),
    .A3(_13550_),
    .B1(_13646_),
    .X(_13738_));
 sky130_fd_sc_hd__a41o_1 _15197_ (.A1(_13706_),
    .A2(_13459_),
    .A3(_13348_),
    .A4(_13737_),
    .B1(_13738_),
    .X(_13739_));
 sky130_fd_sc_hd__o21a_1 _15198_ (.A1(_13639_),
    .A2(_13657_),
    .B1(_13496_),
    .X(_13740_));
 sky130_fd_sc_hd__and3_1 _15199_ (.A(_13430_),
    .B(_13387_),
    .C(_13320_),
    .X(_13741_));
 sky130_fd_sc_hd__or4b_1 _15200_ (.A(_13385_),
    .B(_13672_),
    .C(_13741_),
    .D_N(_13598_),
    .X(_13742_));
 sky130_fd_sc_hd__or3b_1 _15201_ (.A(_13740_),
    .B(_13499_),
    .C_N(_13742_),
    .X(_13743_));
 sky130_fd_sc_hd__nand2_1 _15202_ (.A(_13526_),
    .B(_13541_),
    .Y(_13744_));
 sky130_fd_sc_hd__a21oi_1 _15203_ (.A1(_13575_),
    .A2(_13744_),
    .B1(_13581_),
    .Y(_13745_));
 sky130_fd_sc_hd__a21oi_1 _15204_ (.A1(_13298_),
    .A2(_13589_),
    .B1(_13616_),
    .Y(_13746_));
 sky130_fd_sc_hd__nand2_1 _15205_ (.A(_13350_),
    .B(_13545_),
    .Y(_13747_));
 sky130_fd_sc_hd__a21o_1 _15206_ (.A1(_13391_),
    .A2(_13523_),
    .B1(_13747_),
    .X(_13748_));
 sky130_fd_sc_hd__a32o_1 _15207_ (.A1(_13364_),
    .A2(_13353_),
    .A3(_13746_),
    .B1(_13748_),
    .B2(_13646_),
    .X(_13749_));
 sky130_fd_sc_hd__nand2_1 _15208_ (.A(_13296_),
    .B(_13393_),
    .Y(_13750_));
 sky130_fd_sc_hd__inv_2 _15209_ (.A(_13493_),
    .Y(_13751_));
 sky130_fd_sc_hd__a21oi_1 _15210_ (.A1(_13750_),
    .A2(_13751_),
    .B1(_13573_),
    .Y(_13752_));
 sky130_fd_sc_hd__or4_1 _15211_ (.A(_13469_),
    .B(_13745_),
    .C(_13749_),
    .D(_13752_),
    .X(_13753_));
 sky130_fd_sc_hd__a211o_1 _15212_ (.A1(_13304_),
    .A2(_13546_),
    .B1(_13465_),
    .C1(_13607_),
    .X(_13754_));
 sky130_fd_sc_hd__nand2_1 _15213_ (.A(_13290_),
    .B(_13444_),
    .Y(_13755_));
 sky130_fd_sc_hd__a22o_1 _15214_ (.A1(_13504_),
    .A2(_13754_),
    .B1(_13755_),
    .B2(_13409_),
    .X(_13756_));
 sky130_fd_sc_hd__or4_1 _15215_ (.A(_13361_),
    .B(_13456_),
    .C(_13555_),
    .D(_13756_),
    .X(_13757_));
 sky130_fd_sc_hd__o211a_1 _15216_ (.A1(_13739_),
    .A2(_13743_),
    .B1(_13753_),
    .C1(_13757_),
    .X(net14));
 sky130_fd_sc_hd__nand2_2 _15217_ (.A(_13343_),
    .B(_13300_),
    .Y(_13758_));
 sky130_fd_sc_hd__nor2_1 _15218_ (.A(_13314_),
    .B(_13758_),
    .Y(_13759_));
 sky130_fd_sc_hd__or2_1 _15219_ (.A(_13372_),
    .B(_13630_),
    .X(_13760_));
 sky130_fd_sc_hd__mux2_1 _15220_ (.A0(_13385_),
    .A1(_13759_),
    .S(_13760_),
    .X(_13761_));
 sky130_fd_sc_hd__and2_1 _15221_ (.A(_13466_),
    .B(_13761_),
    .X(_13762_));
 sky130_fd_sc_hd__nor2_1 _15222_ (.A(_13397_),
    .B(_13282_),
    .Y(_13763_));
 sky130_fd_sc_hd__or3_2 _15223_ (.A(_13332_),
    .B(_13763_),
    .C(_13721_),
    .X(_13764_));
 sky130_fd_sc_hd__a211oi_1 _15224_ (.A1(_13298_),
    .A2(_13717_),
    .B1(_13764_),
    .C1(_13315_),
    .Y(_13765_));
 sky130_fd_sc_hd__o21a_1 _15225_ (.A1(_13402_),
    .A2(_13484_),
    .B1(_13692_),
    .X(_13766_));
 sky130_fd_sc_hd__clkbuf_4 _15226_ (.A(_13285_),
    .X(_13767_));
 sky130_fd_sc_hd__or4_1 _15227_ (.A(_13506_),
    .B(_13767_),
    .C(_13432_),
    .D(_13357_),
    .X(_13768_));
 sky130_fd_sc_hd__o311a_1 _15228_ (.A1(_13682_),
    .A2(_13366_),
    .A3(_13526_),
    .B1(_13768_),
    .C1(_13521_),
    .X(_13769_));
 sky130_fd_sc_hd__o31ai_1 _15229_ (.A1(_13439_),
    .A2(_13581_),
    .A3(_13766_),
    .B1(_13769_),
    .Y(_13770_));
 sky130_fd_sc_hd__or2_1 _15230_ (.A(_13767_),
    .B(_13559_),
    .X(_13771_));
 sky130_fd_sc_hd__a21o_1 _15231_ (.A1(_13360_),
    .A2(_13771_),
    .B1(_13315_),
    .X(_13772_));
 sky130_fd_sc_hd__or2_1 _15232_ (.A(_13331_),
    .B(_13284_),
    .X(_13773_));
 sky130_fd_sc_hd__or3_1 _15233_ (.A(_13378_),
    .B(_13773_),
    .C(_13442_),
    .X(_13774_));
 sky130_fd_sc_hd__nand2_1 _15234_ (.A(_13772_),
    .B(_13774_),
    .Y(_13775_));
 sky130_fd_sc_hd__o32a_1 _15235_ (.A1(_13762_),
    .A2(_13765_),
    .A3(_13770_),
    .B1(_13775_),
    .B2(_13572_),
    .X(net12));
 sky130_fd_sc_hd__a31o_2 _15236_ (.A1(_13346_),
    .A2(_13393_),
    .A3(_13592_),
    .B1(_13285_),
    .X(_13776_));
 sky130_fd_sc_hd__inv_2 _15237_ (.A(_13776_),
    .Y(_13777_));
 sky130_fd_sc_hd__a221o_1 _15238_ (.A1(_13542_),
    .A2(_13525_),
    .B1(_13717_),
    .B2(_13317_),
    .C1(_13438_),
    .X(_13778_));
 sky130_fd_sc_hd__or3_1 _15239_ (.A(_13419_),
    .B(_13323_),
    .C(_13750_),
    .X(_13779_));
 sky130_fd_sc_hd__nand2_4 _15240_ (.A(_13305_),
    .B(_13346_),
    .Y(_13780_));
 sky130_fd_sc_hd__nand2_1 _15241_ (.A(_13721_),
    .B(_13780_),
    .Y(_13781_));
 sky130_fd_sc_hd__a31o_1 _15242_ (.A1(_13428_),
    .A2(_13703_),
    .A3(_13574_),
    .B1(_13312_),
    .X(_13782_));
 sky130_fd_sc_hd__a31o_1 _15243_ (.A1(_13352_),
    .A2(_13779_),
    .A3(_13781_),
    .B1(_13782_),
    .X(_13783_));
 sky130_fd_sc_hd__o211a_1 _15244_ (.A1(_13777_),
    .A2(_13778_),
    .B1(_13783_),
    .C1(_13501_),
    .X(_13784_));
 sky130_fd_sc_hd__nand2_1 _15245_ (.A(_13599_),
    .B(_13379_),
    .Y(_13785_));
 sky130_fd_sc_hd__o32a_1 _15246_ (.A1(_13358_),
    .A2(_13432_),
    .A3(_13488_),
    .B1(_13685_),
    .B2(_13598_),
    .X(_13786_));
 sky130_fd_sc_hd__a31o_1 _15247_ (.A1(_13785_),
    .A2(_13773_),
    .A3(_13786_),
    .B1(_13458_),
    .X(_13787_));
 sky130_fd_sc_hd__or4_1 _15248_ (.A(_13343_),
    .B(_13321_),
    .C(_13401_),
    .D(_13354_),
    .X(_13788_));
 sky130_fd_sc_hd__o311a_1 _15249_ (.A1(_13501_),
    .A2(_13566_),
    .A3(_13659_),
    .B1(_13787_),
    .C1(_13788_),
    .X(_13789_));
 sky130_fd_sc_hd__nand2_1 _15250_ (.A(_13638_),
    .B(_13789_),
    .Y(_13790_));
 sky130_fd_sc_hd__a211o_1 _15251_ (.A1(_13329_),
    .A2(_13744_),
    .B1(_13483_),
    .C1(\rvcpu.dp.pcreg.q[8] ),
    .X(_13791_));
 sky130_fd_sc_hd__nand2_1 _15252_ (.A(_13539_),
    .B(_13791_),
    .Y(_13792_));
 sky130_fd_sc_hd__and4_1 _15253_ (.A(_13284_),
    .B(_13307_),
    .C(_13289_),
    .D(_13403_),
    .X(_13793_));
 sky130_fd_sc_hd__or3_1 _15254_ (.A(_13373_),
    .B(_13416_),
    .C(_13793_),
    .X(_13794_));
 sky130_fd_sc_hd__nor2_1 _15255_ (.A(_13438_),
    .B(_13794_),
    .Y(_13795_));
 sky130_fd_sc_hd__nand2_2 _15256_ (.A(_13284_),
    .B(_13425_),
    .Y(_13796_));
 sky130_fd_sc_hd__nand2_1 _15257_ (.A(_13369_),
    .B(_13796_),
    .Y(_13797_));
 sky130_fd_sc_hd__or3b_1 _15258_ (.A(_13291_),
    .B(_13337_),
    .C_N(_13797_),
    .X(_13798_));
 sky130_fd_sc_hd__a31o_1 _15259_ (.A1(_13675_),
    .A2(_13776_),
    .A3(_13798_),
    .B1(_13441_),
    .X(_13799_));
 sky130_fd_sc_hd__or2_1 _15260_ (.A(_13320_),
    .B(_13434_),
    .X(_13800_));
 sky130_fd_sc_hd__o21ai_1 _15261_ (.A1(_13430_),
    .A2(_13628_),
    .B1(_13484_),
    .Y(_13801_));
 sky130_fd_sc_hd__a32oi_2 _15262_ (.A1(_13420_),
    .A2(_13514_),
    .A3(_13800_),
    .B1(_13801_),
    .B2(_13503_),
    .Y(_13802_));
 sky130_fd_sc_hd__o311a_1 _15263_ (.A1(_13366_),
    .A2(_13416_),
    .A3(_13671_),
    .B1(_13799_),
    .C1(_13802_),
    .X(_13803_));
 sky130_fd_sc_hd__or4b_1 _15264_ (.A(_13355_),
    .B(_13792_),
    .C(_13795_),
    .D_N(_13803_),
    .X(_13804_));
 sky130_fd_sc_hd__o21a_1 _15265_ (.A1(_13784_),
    .A2(_13790_),
    .B1(_13804_),
    .X(net11));
 sky130_fd_sc_hd__nand2_1 _15266_ (.A(_13431_),
    .B(_13589_),
    .Y(_13805_));
 sky130_fd_sc_hd__a21oi_1 _15267_ (.A1(_13805_),
    .A2(_13758_),
    .B1(_13533_),
    .Y(_13806_));
 sky130_fd_sc_hd__or3_1 _15268_ (.A(_13449_),
    .B(_13658_),
    .C(_13671_),
    .X(_13807_));
 sky130_fd_sc_hd__a221o_1 _15269_ (.A1(_13463_),
    .A2(_13728_),
    .B1(_13807_),
    .B2(_13428_),
    .C1(_13412_),
    .X(_13808_));
 sky130_fd_sc_hd__nor2_1 _15270_ (.A(_13401_),
    .B(_13451_),
    .Y(_13809_));
 sky130_fd_sc_hd__o21a_1 _15271_ (.A1(_13435_),
    .A2(_13809_),
    .B1(_13353_),
    .X(_13810_));
 sky130_fd_sc_hd__nand2_1 _15272_ (.A(_13332_),
    .B(_13363_),
    .Y(_13811_));
 sky130_fd_sc_hd__a21o_1 _15273_ (.A1(_13307_),
    .A2(_13689_),
    .B1(_13811_),
    .X(_13812_));
 sky130_fd_sc_hd__or4_1 _15274_ (.A(_13300_),
    .B(_13767_),
    .C(_13488_),
    .D(_13401_),
    .X(_13813_));
 sky130_fd_sc_hd__a31o_1 _15275_ (.A1(_13385_),
    .A2(_13812_),
    .A3(_13813_),
    .B1(_13783_),
    .X(_13814_));
 sky130_fd_sc_hd__o31a_1 _15276_ (.A1(_13806_),
    .A2(_13808_),
    .A3(_13810_),
    .B1(_13814_),
    .X(_13815_));
 sky130_fd_sc_hd__a31o_1 _15277_ (.A1(_13630_),
    .A2(_13776_),
    .A3(_13798_),
    .B1(_13441_),
    .X(_13816_));
 sky130_fd_sc_hd__a21o_1 _15278_ (.A1(_13599_),
    .A2(_13536_),
    .B1(_13802_),
    .X(_13817_));
 sky130_fd_sc_hd__a31o_1 _15279_ (.A1(_13328_),
    .A2(_13692_),
    .A3(_13414_),
    .B1(_13366_),
    .X(_13818_));
 sky130_fd_sc_hd__o211a_1 _15280_ (.A1(_13412_),
    .A2(_13794_),
    .B1(_13818_),
    .C1(_13791_),
    .X(_13819_));
 sky130_fd_sc_hd__a31o_1 _15281_ (.A1(_13816_),
    .A2(_13817_),
    .A3(_13819_),
    .B1(_13521_),
    .X(_13820_));
 sky130_fd_sc_hd__a21bo_1 _15282_ (.A1(_13638_),
    .A2(_13815_),
    .B1_N(_13820_),
    .X(_13821_));
 sky130_fd_sc_hd__buf_1 _15283_ (.A(_13821_),
    .X(net10));
 sky130_fd_sc_hd__a31o_1 _15284_ (.A1(_13419_),
    .A2(_13370_),
    .A3(_13496_),
    .B1(_13469_),
    .X(_13822_));
 sky130_fd_sc_hd__clkbuf_4 _15285_ (.A(_13599_),
    .X(_13823_));
 sky130_fd_sc_hd__nand2_1 _15286_ (.A(_13392_),
    .B(_13523_),
    .Y(_13824_));
 sky130_fd_sc_hd__nand3_1 _15287_ (.A(_13823_),
    .B(_13350_),
    .C(_13824_),
    .Y(_13825_));
 sky130_fd_sc_hd__a21o_1 _15288_ (.A1(_13604_),
    .A2(_13505_),
    .B1(_13764_),
    .X(_13826_));
 sky130_fd_sc_hd__o21ai_1 _15289_ (.A1(_13682_),
    .A2(_13780_),
    .B1(_13805_),
    .Y(_13827_));
 sky130_fd_sc_hd__a32o_1 _15290_ (.A1(_13706_),
    .A2(_13825_),
    .A3(_13826_),
    .B1(_13827_),
    .B2(_13429_),
    .X(_13828_));
 sky130_fd_sc_hd__or4_1 _15291_ (.A(_13430_),
    .B(_13506_),
    .C(_13447_),
    .D(_13654_),
    .X(_13829_));
 sky130_fd_sc_hd__a21oi_1 _15292_ (.A1(_13643_),
    .A2(_13829_),
    .B1(_13581_),
    .Y(_13830_));
 sky130_fd_sc_hd__or2_1 _15293_ (.A(_13415_),
    .B(_13510_),
    .X(_13831_));
 sky130_fd_sc_hd__or3_1 _15294_ (.A(_13298_),
    .B(_13488_),
    .C(_13447_),
    .X(_13832_));
 sky130_fd_sc_hd__a31o_1 _15295_ (.A1(_13430_),
    .A2(_13375_),
    .A3(_13348_),
    .B1(_13614_),
    .X(_13833_));
 sky130_fd_sc_hd__and3b_1 _15296_ (.A_N(_13547_),
    .B(_13833_),
    .C(_13385_),
    .X(_13834_));
 sky130_fd_sc_hd__a31o_1 _15297_ (.A1(_13496_),
    .A2(_13831_),
    .A3(_13832_),
    .B1(_13834_),
    .X(_13835_));
 sky130_fd_sc_hd__o311a_1 _15298_ (.A1(_13432_),
    .A2(_13322_),
    .A3(_13796_),
    .B1(_13776_),
    .C1(_13370_),
    .X(_13836_));
 sky130_fd_sc_hd__a21oi_1 _15299_ (.A1(_13559_),
    .A2(_13689_),
    .B1(_13639_),
    .Y(_13837_));
 sky130_fd_sc_hd__a22o_1 _15300_ (.A1(_13449_),
    .A2(_13389_),
    .B1(_13509_),
    .B2(_13763_),
    .X(_13838_));
 sky130_fd_sc_hd__nand2_1 _15301_ (.A(_13463_),
    .B(_13838_),
    .Y(_13839_));
 sky130_fd_sc_hd__o221a_1 _15302_ (.A1(_13385_),
    .A2(_13836_),
    .B1(_13837_),
    .B2(_13374_),
    .C1(_13839_),
    .X(_13840_));
 sky130_fd_sc_hd__or4_1 _15303_ (.A(_13419_),
    .B(_13293_),
    .C(_13482_),
    .D(_13505_),
    .X(_13841_));
 sky130_fd_sc_hd__a21o_1 _15304_ (.A1(_13487_),
    .A2(_13350_),
    .B1(_13513_),
    .X(_13842_));
 sky130_fd_sc_hd__and3_1 _15305_ (.A(_13312_),
    .B(_13841_),
    .C(_13842_),
    .X(_13843_));
 sky130_fd_sc_hd__o311a_1 _15306_ (.A1(_13423_),
    .A2(_13561_),
    .A3(_13657_),
    .B1(_13794_),
    .C1(_13843_),
    .X(_13844_));
 sky130_fd_sc_hd__a21oi_1 _15307_ (.A1(_13466_),
    .A2(_13840_),
    .B1(_13844_),
    .Y(_13845_));
 sky130_fd_sc_hd__o32a_1 _15308_ (.A1(_13499_),
    .A2(_13830_),
    .A3(_13835_),
    .B1(_13845_),
    .B2(_13638_),
    .X(_13846_));
 sky130_fd_sc_hd__o21a_1 _15309_ (.A1(_13822_),
    .A2(_13828_),
    .B1(_13846_),
    .X(net9));
 sky130_fd_sc_hd__nand2_1 _15310_ (.A(_13414_),
    .B(_13562_),
    .Y(_13847_));
 sky130_fd_sc_hd__o221ai_1 _15311_ (.A1(_13767_),
    .A2(_13324_),
    .B1(_13847_),
    .B2(_13823_),
    .C1(_13319_),
    .Y(_13848_));
 sky130_fd_sc_hd__a31o_1 _15312_ (.A1(_13823_),
    .A2(_13420_),
    .A3(_13693_),
    .B1(_13848_),
    .X(_13849_));
 sky130_fd_sc_hd__inv_2 _15313_ (.A(_13392_),
    .Y(_13850_));
 sky130_fd_sc_hd__o32a_1 _15314_ (.A1(_13850_),
    .A2(_13447_),
    .A3(_13309_),
    .B1(_13598_),
    .B2(_13509_),
    .X(_13851_));
 sky130_fd_sc_hd__nor2_1 _15315_ (.A(_13542_),
    .B(_13851_),
    .Y(_13852_));
 sky130_fd_sc_hd__nor2_1 _15316_ (.A(_13494_),
    .B(_13780_),
    .Y(_13853_));
 sky130_fd_sc_hd__a21oi_1 _15317_ (.A1(_13398_),
    .A2(_13672_),
    .B1(_13853_),
    .Y(_13854_));
 sky130_fd_sc_hd__or3_1 _15318_ (.A(_13366_),
    .B(_13301_),
    .C(_13426_),
    .X(_13855_));
 sky130_fd_sc_hd__o311a_1 _15319_ (.A1(_13359_),
    .A2(_13410_),
    .A3(_13465_),
    .B1(_13855_),
    .C1(\rvcpu.dp.pcreg.q[9] ),
    .X(_13856_));
 sky130_fd_sc_hd__a21o_1 _15320_ (.A1(_13548_),
    .A2(_13847_),
    .B1(_13599_),
    .X(_13857_));
 sky130_fd_sc_hd__or2_2 _15321_ (.A(_13307_),
    .B(_13350_),
    .X(_13858_));
 sky130_fd_sc_hd__or3_1 _15322_ (.A(_13292_),
    .B(_13301_),
    .C(_13510_),
    .X(_13859_));
 sky130_fd_sc_hd__a31o_1 _15323_ (.A1(_13857_),
    .A2(_13858_),
    .A3(_13859_),
    .B1(_13501_),
    .X(_13860_));
 sky130_fd_sc_hd__o311a_1 _15324_ (.A1(_13442_),
    .A2(_13852_),
    .A3(_13854_),
    .B1(_13856_),
    .C1(_13860_),
    .X(_13861_));
 sky130_fd_sc_hd__nand2_1 _15325_ (.A(_13517_),
    .B(_13563_),
    .Y(_13862_));
 sky130_fd_sc_hd__a21o_1 _15326_ (.A1(_13798_),
    .A2(_13862_),
    .B1(_13442_),
    .X(_13863_));
 sky130_fd_sc_hd__nand2_1 _15327_ (.A(_13608_),
    .B(_13578_),
    .Y(_13864_));
 sky130_fd_sc_hd__nand2_1 _15328_ (.A(_13615_),
    .B(_13472_),
    .Y(_13865_));
 sky130_fd_sc_hd__o32a_1 _15329_ (.A1(_13449_),
    .A2(_13694_),
    .A3(_13865_),
    .B1(_13455_),
    .B2(_13357_),
    .X(_13866_));
 sky130_fd_sc_hd__nor2_1 _15330_ (.A(_13430_),
    .B(_13399_),
    .Y(_13867_));
 sky130_fd_sc_hd__o21ai_1 _15331_ (.A1(_13867_),
    .A2(_13639_),
    .B1(_13514_),
    .Y(_13868_));
 sky130_fd_sc_hd__o31a_1 _15332_ (.A1(_13366_),
    .A2(_13308_),
    .A3(_13598_),
    .B1(_13868_),
    .X(_13869_));
 sky130_fd_sc_hd__and4b_1 _15333_ (.A_N(_13792_),
    .B(_13864_),
    .C(_13866_),
    .D(_13869_),
    .X(_13870_));
 sky130_fd_sc_hd__o311a_1 _15334_ (.A1(_13410_),
    .A2(_13416_),
    .A3(_13590_),
    .B1(_13863_),
    .C1(_13870_),
    .X(_13871_));
 sky130_fd_sc_hd__a21oi_1 _15335_ (.A1(_13849_),
    .A2(_13861_),
    .B1(_13871_),
    .Y(net8));
 sky130_fd_sc_hd__or2_1 _15336_ (.A(_13509_),
    .B(_13565_),
    .X(_13872_));
 sky130_fd_sc_hd__a221o_1 _15337_ (.A1(_13692_),
    .A2(_13322_),
    .B1(_13872_),
    .B2(_13517_),
    .C1(_13458_),
    .X(_13873_));
 sky130_fd_sc_hd__nor2_1 _15338_ (.A(_13696_),
    .B(_13873_),
    .Y(_13874_));
 sky130_fd_sc_hd__a31o_1 _15339_ (.A1(_13409_),
    .A2(_13459_),
    .A3(_13488_),
    .B1(_13521_),
    .X(_13875_));
 sky130_fd_sc_hd__nor2_2 _15340_ (.A(_13414_),
    .B(_13336_),
    .Y(_13876_));
 sky130_fd_sc_hd__and3_1 _15341_ (.A(_13368_),
    .B(_13646_),
    .C(_13876_),
    .X(_13877_));
 sky130_fd_sc_hd__a21o_1 _15342_ (.A1(_13608_),
    .A2(_13528_),
    .B1(_13539_),
    .X(_13878_));
 sky130_fd_sc_hd__a21oi_1 _15343_ (.A1(_13668_),
    .A2(_13489_),
    .B1(_13374_),
    .Y(_13879_));
 sky130_fd_sc_hd__nor2_1 _15344_ (.A(_13387_),
    .B(_13750_),
    .Y(_13880_));
 sky130_fd_sc_hd__a211o_1 _15345_ (.A1(_13332_),
    .A2(_13307_),
    .B1(_13350_),
    .C1(_13314_),
    .X(_13881_));
 sky130_fd_sc_hd__a21bo_1 _15346_ (.A1(_13428_),
    .A2(_13880_),
    .B1_N(_13881_),
    .X(_13882_));
 sky130_fd_sc_hd__a211o_1 _15347_ (.A1(_13291_),
    .A2(_13343_),
    .B1(_13352_),
    .C1(_13759_),
    .X(_13883_));
 sky130_fd_sc_hd__o31a_1 _15348_ (.A1(_13422_),
    .A2(_13465_),
    .A3(_13622_),
    .B1(_13883_),
    .X(_13884_));
 sky130_fd_sc_hd__a41o_1 _15349_ (.A1(_13431_),
    .A2(_13526_),
    .A3(_13428_),
    .A4(_13737_),
    .B1(_13312_),
    .X(_13885_));
 sky130_fd_sc_hd__o32a_1 _15350_ (.A1(_13438_),
    .A2(_13879_),
    .A3(_13882_),
    .B1(_13884_),
    .B2(_13885_),
    .X(_13886_));
 sky130_fd_sc_hd__a211o_1 _15351_ (.A1(_13608_),
    .A2(_13690_),
    .B1(_13878_),
    .C1(_13886_),
    .X(_13887_));
 sky130_fd_sc_hd__o31a_1 _15352_ (.A1(_13874_),
    .A2(_13875_),
    .A3(_13877_),
    .B1(_13887_),
    .X(net7));
 sky130_fd_sc_hd__a211o_1 _15353_ (.A1(_13693_),
    .A2(_13780_),
    .B1(_13435_),
    .C1(_13581_),
    .X(_13888_));
 sky130_fd_sc_hd__o31ai_1 _15354_ (.A1(_13528_),
    .A2(_13359_),
    .A3(_13634_),
    .B1(_13463_),
    .Y(_13889_));
 sky130_fd_sc_hd__o21a_1 _15355_ (.A1(_13665_),
    .A2(_13668_),
    .B1(_13610_),
    .X(_13890_));
 sky130_fd_sc_hd__o21a_1 _15356_ (.A1(_13533_),
    .A2(_13890_),
    .B1(_13478_),
    .X(_13891_));
 sky130_fd_sc_hd__a31o_1 _15357_ (.A1(_13888_),
    .A2(_13889_),
    .A3(_13891_),
    .B1(_13439_),
    .X(_13892_));
 sky130_fd_sc_hd__nor2_2 _15358_ (.A(_13332_),
    .B(_13634_),
    .Y(_13893_));
 sky130_fd_sc_hd__a311o_1 _15359_ (.A1(_13358_),
    .A2(_13545_),
    .A3(_13758_),
    .B1(_13893_),
    .C1(_13441_),
    .X(_13894_));
 sky130_fd_sc_hd__o211a_1 _15360_ (.A1(_13368_),
    .A2(_13498_),
    .B1(_13894_),
    .C1(\rvcpu.dp.pcreg.q[9] ),
    .X(_13895_));
 sky130_fd_sc_hd__a31o_1 _15361_ (.A1(_13370_),
    .A2(_13862_),
    .A3(_13858_),
    .B1(_13442_),
    .X(_13896_));
 sky130_fd_sc_hd__or2_1 _15362_ (.A(_13466_),
    .B(_13841_),
    .X(_13897_));
 sky130_fd_sc_hd__o21ai_1 _15363_ (.A1(_13528_),
    .A2(_13512_),
    .B1(_13514_),
    .Y(_13898_));
 sky130_fd_sc_hd__nor2_1 _15364_ (.A(_13638_),
    .B(_13537_),
    .Y(_13899_));
 sky130_fd_sc_hd__o21ba_1 _15365_ (.A1(_13472_),
    .A2(_13589_),
    .B1_N(_13417_),
    .X(_13900_));
 sky130_fd_sc_hd__o21ai_1 _15366_ (.A1(_13549_),
    .A2(_13900_),
    .B1(_13409_),
    .Y(_13901_));
 sky130_fd_sc_hd__o2111a_1 _15367_ (.A1(_13343_),
    .A2(_13897_),
    .B1(_13898_),
    .C1(_13899_),
    .D1(_13901_),
    .X(_13902_));
 sky130_fd_sc_hd__a32o_1 _15368_ (.A1(_13774_),
    .A2(_13892_),
    .A3(_13895_),
    .B1(_13896_),
    .B2(_13902_),
    .X(_13903_));
 sky130_fd_sc_hd__inv_2 _15369_ (.A(_13903_),
    .Y(net6));
 sky130_fd_sc_hd__a31oi_1 _15370_ (.A1(_13368_),
    .A2(_13646_),
    .A3(_13793_),
    .B1(_13521_),
    .Y(_13904_));
 sky130_fd_sc_hd__o21ai_1 _15371_ (.A1(_13528_),
    .A2(_13553_),
    .B1(_13514_),
    .Y(_13905_));
 sky130_fd_sc_hd__or3_1 _15372_ (.A(_13694_),
    .B(_13656_),
    .C(_13865_),
    .X(_13906_));
 sky130_fd_sc_hd__a21o_1 _15373_ (.A1(_13407_),
    .A2(_13448_),
    .B1(_13366_),
    .X(_13907_));
 sky130_fd_sc_hd__o2111a_1 _15374_ (.A1(_13785_),
    .A2(_13501_),
    .B1(_13905_),
    .C1(_13906_),
    .D1(_13907_),
    .X(_13908_));
 sky130_fd_sc_hd__nor2_1 _15375_ (.A(_13304_),
    .B(_13425_),
    .Y(_13909_));
 sky130_fd_sc_hd__or3_1 _15376_ (.A(_13909_),
    .B(_13471_),
    .C(_13690_),
    .X(_13910_));
 sky130_fd_sc_hd__o311a_1 _15377_ (.A1(_13359_),
    .A2(_13474_),
    .A3(_13634_),
    .B1(_13910_),
    .C1(_13409_),
    .X(_13911_));
 sky130_fd_sc_hd__a21oi_1 _15378_ (.A1(_13419_),
    .A2(_13370_),
    .B1(_13416_),
    .Y(_13912_));
 sky130_fd_sc_hd__or4_1 _15379_ (.A(_13308_),
    .B(_13767_),
    .C(_13357_),
    .D(_13654_),
    .X(_13913_));
 sky130_fd_sc_hd__or3_1 _15380_ (.A(_13432_),
    .B(_13773_),
    .C(_13441_),
    .X(_13914_));
 sky130_fd_sc_hd__o2bb2a_1 _15381_ (.A1_N(_13382_),
    .A2_N(_13319_),
    .B1(_13349_),
    .B2(_13914_),
    .X(_13915_));
 sky130_fd_sc_hd__o311a_1 _15382_ (.A1(_13412_),
    .A2(_13483_),
    .A3(_13912_),
    .B1(_13913_),
    .C1(_13915_),
    .X(_13916_));
 sky130_fd_sc_hd__and3b_1 _15383_ (.A_N(_13911_),
    .B(_13916_),
    .C(_13895_),
    .X(_13917_));
 sky130_fd_sc_hd__a21oi_1 _15384_ (.A1(_13904_),
    .A2(_13908_),
    .B1(_13917_),
    .Y(net5));
 sky130_fd_sc_hd__o21a_1 _15385_ (.A1(_13528_),
    .A2(_13634_),
    .B1(_13646_),
    .X(_13918_));
 sky130_fd_sc_hd__a211oi_1 _15386_ (.A1(_13706_),
    .A2(_13339_),
    .B1(_13918_),
    .C1(_13439_),
    .Y(_13919_));
 sky130_fd_sc_hd__or3b_1 _15387_ (.A(_13309_),
    .B(_13581_),
    .C_N(_13451_),
    .X(_13920_));
 sky130_fd_sc_hd__or3_1 _15388_ (.A(_13297_),
    .B(_13422_),
    .C(_13586_),
    .X(_13921_));
 sky130_fd_sc_hd__nand2_1 _15389_ (.A(_13496_),
    .B(_13443_),
    .Y(_13922_));
 sky130_fd_sc_hd__o311a_1 _15390_ (.A1(_13298_),
    .A2(_13374_),
    .A3(_13604_),
    .B1(_13635_),
    .C1(_13438_),
    .X(_13923_));
 sky130_fd_sc_hd__and3_1 _15391_ (.A(_13464_),
    .B(_13922_),
    .C(_13923_),
    .X(_13924_));
 sky130_fd_sc_hd__a31o_1 _15392_ (.A1(_13919_),
    .A2(_13920_),
    .A3(_13921_),
    .B1(_13924_),
    .X(_13925_));
 sky130_fd_sc_hd__a2bb2o_1 _15393_ (.A1_N(_13419_),
    .A2_N(_13603_),
    .B1(_13381_),
    .B2(_13599_),
    .X(_13926_));
 sky130_fd_sc_hd__o21ai_1 _15394_ (.A1(_13665_),
    .A2(_13323_),
    .B1(_13666_),
    .Y(_13927_));
 sky130_fd_sc_hd__a221o_1 _15395_ (.A1(_13327_),
    .A2(_13926_),
    .B1(_13927_),
    .B2(_13504_),
    .C1(_13521_),
    .X(_13928_));
 sky130_fd_sc_hd__nand2_1 _15396_ (.A(_13434_),
    .B(_13574_),
    .Y(_13929_));
 sky130_fd_sc_hd__a211o_1 _15397_ (.A1(_13378_),
    .A2(_13929_),
    .B1(_13590_),
    .C1(_13410_),
    .X(_13930_));
 sky130_fd_sc_hd__and4b_1 _15398_ (.A_N(_13928_),
    .B(_13930_),
    .C(_13897_),
    .D(_13864_),
    .X(_13931_));
 sky130_fd_sc_hd__a21o_1 _15399_ (.A1(_13572_),
    .A2(_13925_),
    .B1(_13931_),
    .X(_13932_));
 sky130_fd_sc_hd__inv_2 _15400_ (.A(_13932_),
    .Y(net4));
 sky130_fd_sc_hd__a21oi_1 _15401_ (.A1(_13496_),
    .A2(_13523_),
    .B1(_13368_),
    .Y(_13933_));
 sky130_fd_sc_hd__o211ai_1 _15402_ (.A1(_13593_),
    .A2(_13764_),
    .B1(_13385_),
    .C1(_13360_),
    .Y(_13934_));
 sky130_fd_sc_hd__o311a_1 _15403_ (.A1(_13483_),
    .A2(_13416_),
    .A3(_13741_),
    .B1(_13921_),
    .C1(_13934_),
    .X(_13935_));
 sky130_fd_sc_hd__a22o_1 _15404_ (.A1(_13402_),
    .A2(_13505_),
    .B1(_13737_),
    .B2(_13431_),
    .X(_13936_));
 sky130_fd_sc_hd__or2_1 _15405_ (.A(_13449_),
    .B(_13718_),
    .X(_13937_));
 sky130_fd_sc_hd__a22o_1 _15406_ (.A1(_13429_),
    .A2(_13936_),
    .B1(_13937_),
    .B2(_13353_),
    .X(_13938_));
 sky130_fd_sc_hd__o2bb2a_1 _15407_ (.A1_N(_13933_),
    .A2_N(_13935_),
    .B1(_13938_),
    .B2(_13466_),
    .X(_13939_));
 sky130_fd_sc_hd__inv_2 _15408_ (.A(_13649_),
    .Y(_13940_));
 sky130_fd_sc_hd__o21a_1 _15409_ (.A1(_13665_),
    .A2(_13348_),
    .B1(_13940_),
    .X(_13941_));
 sky130_fd_sc_hd__a21oi_1 _15410_ (.A1(_13682_),
    .A2(_13378_),
    .B1(_13941_),
    .Y(_13942_));
 sky130_fd_sc_hd__a21o_1 _15411_ (.A1(_13298_),
    .A2(_13681_),
    .B1(_13507_),
    .X(_13943_));
 sky130_fd_sc_hd__a2bb2o_1 _15412_ (.A1_N(_13410_),
    .A2_N(_13942_),
    .B1(_13943_),
    .B2(_13608_),
    .X(_13944_));
 sky130_fd_sc_hd__a31o_1 _15413_ (.A1(_13392_),
    .A2(_13348_),
    .A3(_13796_),
    .B1(_13513_),
    .X(_13945_));
 sky130_fd_sc_hd__o21ai_1 _15414_ (.A1(_13309_),
    .A2(_13809_),
    .B1(_13428_),
    .Y(_13946_));
 sky130_fd_sc_hd__o311a_1 _15415_ (.A1(_13431_),
    .A2(_13628_),
    .A3(_13423_),
    .B1(_13945_),
    .C1(_13946_),
    .X(_13947_));
 sky130_fd_sc_hd__o31ai_1 _15416_ (.A1(_13533_),
    .A2(_13640_),
    .A3(_13853_),
    .B1(_13947_),
    .Y(_13948_));
 sky130_fd_sc_hd__and2_1 _15417_ (.A(_13305_),
    .B(_13349_),
    .X(_13949_));
 sky130_fd_sc_hd__and3_1 _15418_ (.A(_13425_),
    .B(_13390_),
    .C(_13317_),
    .X(_13950_));
 sky130_fd_sc_hd__a31o_1 _15419_ (.A1(_13459_),
    .A2(_13526_),
    .A3(_13509_),
    .B1(_13950_),
    .X(_13951_));
 sky130_fd_sc_hd__a221o_1 _15420_ (.A1(_13504_),
    .A2(_13949_),
    .B1(_13951_),
    .B2(_13319_),
    .C1(_13539_),
    .X(_13952_));
 sky130_fd_sc_hd__o211a_1 _15421_ (.A1(_13298_),
    .A2(_13341_),
    .B1(_13336_),
    .C1(_13333_),
    .X(_13953_));
 sky130_fd_sc_hd__o21ai_1 _15422_ (.A1(_13324_),
    .A2(_13649_),
    .B1(_13953_),
    .Y(_13954_));
 sky130_fd_sc_hd__o211a_1 _15423_ (.A1(_13940_),
    .A2(_13764_),
    .B1(_13954_),
    .C1(_13327_),
    .X(_13955_));
 sky130_fd_sc_hd__a211o_1 _15424_ (.A1(_13368_),
    .A2(_13948_),
    .B1(_13952_),
    .C1(_13955_),
    .X(_13956_));
 sky130_fd_sc_hd__o31a_1 _15425_ (.A1(_13572_),
    .A2(_13939_),
    .A3(_13944_),
    .B1(_13956_),
    .X(net3));
 sky130_fd_sc_hd__or4_1 _15426_ (.A(_13292_),
    .B(_13401_),
    .C(_13628_),
    .D(_13718_),
    .X(_13957_));
 sky130_fd_sc_hd__o311a_1 _15427_ (.A1(_13542_),
    .A2(_13473_),
    .A3(_13853_),
    .B1(_13957_),
    .C1(_13475_),
    .X(_13958_));
 sky130_fd_sc_hd__or3_1 _15428_ (.A(_13303_),
    .B(_13321_),
    .C(_13454_),
    .X(_13959_));
 sky130_fd_sc_hd__a21oi_1 _15429_ (.A1(_13858_),
    .A2(_13959_),
    .B1(_13423_),
    .Y(_13960_));
 sky130_fd_sc_hd__nor2_1 _15430_ (.A(_13958_),
    .B(_13960_),
    .Y(_13961_));
 sky130_fd_sc_hd__a211o_1 _15431_ (.A1(_13431_),
    .A2(_13432_),
    .B1(_13613_),
    .C1(_13333_),
    .X(_13962_));
 sky130_fd_sc_hd__or3b_1 _15432_ (.A(_13506_),
    .B(_13398_),
    .C_N(_13703_),
    .X(_13963_));
 sky130_fd_sc_hd__a31o_1 _15433_ (.A1(_13785_),
    .A2(_13962_),
    .A3(_13963_),
    .B1(_13458_),
    .X(_13964_));
 sky130_fd_sc_hd__nor2_1 _15434_ (.A(_13509_),
    .B(_13565_),
    .Y(_13965_));
 sky130_fd_sc_hd__a221o_1 _15435_ (.A1(_13517_),
    .A2(_13965_),
    .B1(_13953_),
    .B2(_13448_),
    .C1(_13442_),
    .X(_13966_));
 sky130_fd_sc_hd__a311o_1 _15436_ (.A1(_13451_),
    .A2(_13666_),
    .A3(_13872_),
    .B1(_13483_),
    .C1(_13438_),
    .X(_13967_));
 sky130_fd_sc_hd__a31o_1 _15437_ (.A1(_13964_),
    .A2(_13966_),
    .A3(_13967_),
    .B1(_13539_),
    .X(_13968_));
 sky130_fd_sc_hd__or3b_1 _15438_ (.A(_13533_),
    .B(_13359_),
    .C_N(_13829_),
    .X(_13969_));
 sky130_fd_sc_hd__a21oi_1 _15439_ (.A1(_13692_),
    .A2(_13389_),
    .B1(_13465_),
    .Y(_13970_));
 sky130_fd_sc_hd__a32o_1 _15440_ (.A1(_13358_),
    .A2(_13450_),
    .A3(_13489_),
    .B1(_13758_),
    .B2(_13893_),
    .X(_13971_));
 sky130_fd_sc_hd__o221a_1 _15441_ (.A1(_13573_),
    .A2(_13970_),
    .B1(_13971_),
    .B2(_13475_),
    .C1(_13368_),
    .X(_13972_));
 sky130_fd_sc_hd__o21a_1 _15442_ (.A1(_13431_),
    .A2(_13628_),
    .B1(_13642_),
    .X(_13973_));
 sky130_fd_sc_hd__a21bo_1 _15443_ (.A1(_13328_),
    .A2(_13301_),
    .B1_N(_13858_),
    .X(_13974_));
 sky130_fd_sc_hd__a21o_1 _15444_ (.A1(_13472_),
    .A2(_13565_),
    .B1(_13482_),
    .X(_13975_));
 sky130_fd_sc_hd__o211a_1 _15445_ (.A1(_13374_),
    .A2(_13974_),
    .B1(_13975_),
    .C1(_13412_),
    .X(_13976_));
 sky130_fd_sc_hd__o21ai_1 _15446_ (.A1(_13561_),
    .A2(_13656_),
    .B1(_13353_),
    .Y(_13977_));
 sky130_fd_sc_hd__o211a_1 _15447_ (.A1(_13573_),
    .A2(_13973_),
    .B1(_13976_),
    .C1(_13977_),
    .X(_13978_));
 sky130_fd_sc_hd__a211o_1 _15448_ (.A1(_13969_),
    .A2(_13972_),
    .B1(_13521_),
    .C1(_13978_),
    .X(_13979_));
 sky130_fd_sc_hd__o211ai_2 _15449_ (.A1(_13469_),
    .A2(_13961_),
    .B1(_13968_),
    .C1(_13979_),
    .Y(net33));
 sky130_fd_sc_hd__o21a_1 _15450_ (.A1(_13553_),
    .A2(_13597_),
    .B1(_13564_),
    .X(_13980_));
 sky130_fd_sc_hd__o21ai_1 _15451_ (.A1(_13308_),
    .A2(_13565_),
    .B1(_13832_),
    .Y(_13981_));
 sky130_fd_sc_hd__o31a_1 _15452_ (.A1(_13506_),
    .A2(_13399_),
    .A3(_13593_),
    .B1(_13504_),
    .X(_13982_));
 sky130_fd_sc_hd__a21oi_1 _15453_ (.A1(_13514_),
    .A2(_13981_),
    .B1(_13982_),
    .Y(_13983_));
 sky130_fd_sc_hd__o211a_1 _15454_ (.A1(_13706_),
    .A2(_13980_),
    .B1(_13983_),
    .C1(_13664_),
    .X(_13984_));
 sky130_fd_sc_hd__a211o_1 _15455_ (.A1(_13402_),
    .A2(_13505_),
    .B1(_13294_),
    .C1(_13292_),
    .X(_13985_));
 sky130_fd_sc_hd__or3_1 _15456_ (.A(_13823_),
    .B(_13747_),
    .C(_13929_),
    .X(_13986_));
 sky130_fd_sc_hd__a21oi_1 _15457_ (.A1(_13985_),
    .A2(_13986_),
    .B1(_13501_),
    .Y(_13987_));
 sky130_fd_sc_hd__or4_1 _15458_ (.A(_13682_),
    .B(_13573_),
    .C(_13321_),
    .D(_13402_),
    .X(_13988_));
 sky130_fd_sc_hd__a311o_1 _15459_ (.A1(_13665_),
    .A2(_13346_),
    .A3(_13484_),
    .B1(_13639_),
    .C1(_13581_),
    .X(_13989_));
 sky130_fd_sc_hd__or3b_1 _15460_ (.A(_13607_),
    .B(_13465_),
    .C_N(_13781_),
    .X(_13990_));
 sky130_fd_sc_hd__a21oi_1 _15461_ (.A1(_13559_),
    .A2(_13351_),
    .B1(_13533_),
    .Y(_13991_));
 sky130_fd_sc_hd__a21oi_1 _15462_ (.A1(_13496_),
    .A2(_13990_),
    .B1(_13991_),
    .Y(_13992_));
 sky130_fd_sc_hd__a31o_1 _15463_ (.A1(_13988_),
    .A2(_13989_),
    .A3(_13992_),
    .B1(_13499_),
    .X(_13993_));
 sky130_fd_sc_hd__nor2_1 _15464_ (.A(_13528_),
    .B(_13435_),
    .Y(_13994_));
 sky130_fd_sc_hd__nand2_1 _15465_ (.A(_13893_),
    .B(_13994_),
    .Y(_13995_));
 sky130_fd_sc_hd__nand2_1 _15466_ (.A(_13350_),
    .B(_13995_),
    .Y(_13996_));
 sky130_fd_sc_hd__o21ai_1 _15467_ (.A1(_13381_),
    .A2(_13996_),
    .B1(_13706_),
    .Y(_13997_));
 sky130_fd_sc_hd__or4b_1 _15468_ (.A(_13341_),
    .B(_13302_),
    .C(_13581_),
    .D_N(_13328_),
    .X(_13998_));
 sky130_fd_sc_hd__o21ai_1 _15469_ (.A1(_13341_),
    .A2(_13668_),
    .B1(_13858_),
    .Y(_13999_));
 sky130_fd_sc_hd__nand2_1 _15470_ (.A(_13496_),
    .B(_13999_),
    .Y(_14000_));
 sky130_fd_sc_hd__a31o_1 _15471_ (.A1(_13997_),
    .A2(_13998_),
    .A3(_14000_),
    .B1(_13469_),
    .X(_14001_));
 sky130_fd_sc_hd__o311a_1 _15472_ (.A1(_13572_),
    .A2(_13984_),
    .A3(_13987_),
    .B1(_13993_),
    .C1(_14001_),
    .X(_14002_));
 sky130_fd_sc_hd__inv_2 _15473_ (.A(_14002_),
    .Y(net32));
 sky130_fd_sc_hd__inv_2 _15474_ (.A(_13893_),
    .Y(_14003_));
 sky130_fd_sc_hd__and2_1 _15475_ (.A(_13372_),
    .B(_13867_),
    .X(_14004_));
 sky130_fd_sc_hd__o221a_1 _15476_ (.A1(_13909_),
    .A2(_13811_),
    .B1(_14003_),
    .B2(_14004_),
    .C1(_13319_),
    .X(_14005_));
 sky130_fd_sc_hd__o21ai_1 _15477_ (.A1(_13308_),
    .A2(_13598_),
    .B1(_13600_),
    .Y(_14006_));
 sky130_fd_sc_hd__a31o_1 _15478_ (.A1(_13327_),
    .A2(_13697_),
    .A3(_14006_),
    .B1(_13539_),
    .X(_14007_));
 sky130_fd_sc_hd__or3b_1 _15479_ (.A(_13690_),
    .B(_13292_),
    .C_N(_13693_),
    .X(_14008_));
 sky130_fd_sc_hd__or3_2 _15480_ (.A(_13320_),
    .B(_13285_),
    .C(_13349_),
    .X(_14009_));
 sky130_fd_sc_hd__o311a_1 _15481_ (.A1(_13599_),
    .A2(_13391_),
    .A3(_13510_),
    .B1(_14008_),
    .C1(_14009_),
    .X(_14010_));
 sky130_fd_sc_hd__or3_1 _15482_ (.A(_13297_),
    .B(_13322_),
    .C(_13586_),
    .X(_14011_));
 sky130_fd_sc_hd__a32o_1 _15483_ (.A1(_13542_),
    .A2(_13824_),
    .A3(_14011_),
    .B1(_13994_),
    .B2(_13600_),
    .X(_14012_));
 sky130_fd_sc_hd__a2bb2o_1 _15484_ (.A1_N(_14010_),
    .A2_N(_13501_),
    .B1(_13409_),
    .B2(_14012_),
    .X(_14013_));
 sky130_fd_sc_hd__a211o_1 _15485_ (.A1(_13541_),
    .A2(_13560_),
    .B1(_13880_),
    .C1(_13332_),
    .X(_14014_));
 sky130_fd_sc_hd__o311a_1 _15486_ (.A1(_13321_),
    .A2(_13421_),
    .A3(_13495_),
    .B1(_14014_),
    .C1(_13385_),
    .X(_14015_));
 sky130_fd_sc_hd__a31o_1 _15487_ (.A1(_13682_),
    .A2(_13399_),
    .A3(_13429_),
    .B1(_14015_),
    .X(_14016_));
 sky130_fd_sc_hd__or3b_1 _15488_ (.A(_13358_),
    .B(_13424_),
    .C_N(_13689_),
    .X(_14017_));
 sky130_fd_sc_hd__o311a_1 _15489_ (.A1(_13517_),
    .A2(_13308_),
    .A3(_14004_),
    .B1(_14017_),
    .C1(_13413_),
    .X(_14018_));
 sky130_fd_sc_hd__a221o_1 _15490_ (.A1(_13439_),
    .A2(_14016_),
    .B1(_14018_),
    .B2(_13776_),
    .C1(_13638_),
    .X(_14019_));
 sky130_fd_sc_hd__o31a_1 _15491_ (.A1(_14005_),
    .A2(_14007_),
    .A3(_14013_),
    .B1(_14019_),
    .X(net31));
 sky130_fd_sc_hd__nor2_1 _15492_ (.A(_13308_),
    .B(_13654_),
    .Y(_14020_));
 sky130_fd_sc_hd__o21ai_1 _15493_ (.A1(_13682_),
    .A2(_14020_),
    .B1(_13599_),
    .Y(_14021_));
 sky130_fd_sc_hd__a21oi_1 _15494_ (.A1(_13800_),
    .A2(_13893_),
    .B1(_13475_),
    .Y(_14022_));
 sky130_fd_sc_hd__o211a_1 _15495_ (.A1(_13337_),
    .A2(_13474_),
    .B1(_13995_),
    .C1(_13475_),
    .X(_14023_));
 sky130_fd_sc_hd__a21oi_1 _15496_ (.A1(_14021_),
    .A2(_14022_),
    .B1(_14023_),
    .Y(_14024_));
 sky130_fd_sc_hd__a21oi_1 _15497_ (.A1(_13517_),
    .A2(_13337_),
    .B1(_13853_),
    .Y(_14025_));
 sky130_fd_sc_hd__a211o_1 _15498_ (.A1(_13425_),
    .A2(_13847_),
    .B1(_13465_),
    .C1(_13513_),
    .X(_14026_));
 sky130_fd_sc_hd__a221o_1 _15499_ (.A1(_13370_),
    .A2(_13348_),
    .B1(_13505_),
    .B2(_13425_),
    .C1(_13374_),
    .X(_14027_));
 sky130_fd_sc_hd__o211a_1 _15500_ (.A1(_13475_),
    .A2(_14025_),
    .B1(_14026_),
    .C1(_14027_),
    .X(_14028_));
 sky130_fd_sc_hd__o31a_1 _15501_ (.A1(_13398_),
    .A2(_13488_),
    .A3(_13402_),
    .B1(_14009_),
    .X(_14029_));
 sky130_fd_sc_hd__o21ai_1 _15502_ (.A1(_13381_),
    .A2(_13876_),
    .B1(_13504_),
    .Y(_14030_));
 sky130_fd_sc_hd__o221a_1 _15503_ (.A1(_13458_),
    .A2(_13360_),
    .B1(_14029_),
    .B2(_13357_),
    .C1(_14030_),
    .X(_14031_));
 sky130_fd_sc_hd__o22a_1 _15504_ (.A1(_13499_),
    .A2(_14028_),
    .B1(_14031_),
    .B2(_13638_),
    .X(_14032_));
 sky130_fd_sc_hd__o21ai_2 _15505_ (.A1(_13469_),
    .A2(_14024_),
    .B1(_14032_),
    .Y(net30));
 sky130_fd_sc_hd__o21bai_1 _15506_ (.A1(_13454_),
    .A2(_13613_),
    .B1_N(_13597_),
    .Y(_14033_));
 sky130_fd_sc_hd__or3b_1 _15507_ (.A(_13322_),
    .B(_13492_),
    .C_N(_13394_),
    .X(_14034_));
 sky130_fd_sc_hd__o311a_1 _15508_ (.A1(_13542_),
    .A2(_13372_),
    .A3(_13510_),
    .B1(_14033_),
    .C1(_14034_),
    .X(_14035_));
 sky130_fd_sc_hd__nor2_1 _15509_ (.A(_13458_),
    .B(_14035_),
    .Y(_14036_));
 sky130_fd_sc_hd__nand2_1 _15510_ (.A(_13542_),
    .B(_13622_),
    .Y(_14037_));
 sky130_fd_sc_hd__a211o_1 _15511_ (.A1(_13297_),
    .A2(_13546_),
    .B1(_13294_),
    .C1(_13292_),
    .X(_14038_));
 sky130_fd_sc_hd__a21oi_1 _15512_ (.A1(_14009_),
    .A2(_14038_),
    .B1(_13357_),
    .Y(_14039_));
 sky130_fd_sc_hd__a31o_1 _15513_ (.A1(_13326_),
    .A2(_13585_),
    .A3(_14037_),
    .B1(_14039_),
    .X(_14040_));
 sky130_fd_sc_hd__a31o_1 _15514_ (.A1(_13409_),
    .A2(_13310_),
    .A3(_13617_),
    .B1(_14040_),
    .X(_14041_));
 sky130_fd_sc_hd__o32a_1 _15515_ (.A1(_13542_),
    .A2(_13531_),
    .A3(_13698_),
    .B1(_13648_),
    .B2(_14021_),
    .X(_14042_));
 sky130_fd_sc_hd__o22a_1 _15516_ (.A1(_13767_),
    .A2(_13389_),
    .B1(_13780_),
    .B2(_13430_),
    .X(_14043_));
 sky130_fd_sc_hd__or2b_1 _15517_ (.A(_13659_),
    .B_N(_14043_),
    .X(_14044_));
 sky130_fd_sc_hd__and3_1 _15518_ (.A(_13327_),
    .B(_13771_),
    .C(_14044_),
    .X(_14045_));
 sky130_fd_sc_hd__nand2_1 _15519_ (.A(_13737_),
    .B(_13656_),
    .Y(_14046_));
 sky130_fd_sc_hd__a31o_1 _15520_ (.A1(_13504_),
    .A2(_13831_),
    .A3(_13577_),
    .B1(_13538_),
    .X(_14047_));
 sky130_fd_sc_hd__mux2_1 _15521_ (.A0(_13949_),
    .A1(_14020_),
    .S(_13304_),
    .X(_14048_));
 sky130_fd_sc_hd__a21o_1 _15522_ (.A1(_13893_),
    .A2(_13959_),
    .B1(_13315_),
    .X(_14049_));
 sky130_fd_sc_hd__a21oi_1 _15523_ (.A1(_13599_),
    .A2(_14048_),
    .B1(_14049_),
    .Y(_14050_));
 sky130_fd_sc_hd__a311o_1 _15524_ (.A1(_13514_),
    .A2(_13796_),
    .A3(_14046_),
    .B1(_14047_),
    .C1(_14050_),
    .X(_14051_));
 sky130_fd_sc_hd__a211o_1 _15525_ (.A1(_13413_),
    .A2(_14042_),
    .B1(_14045_),
    .C1(_14051_),
    .X(_14052_));
 sky130_fd_sc_hd__o31a_1 _15526_ (.A1(_13572_),
    .A2(_14036_),
    .A3(_14041_),
    .B1(_14052_),
    .X(net29));
 sky130_fd_sc_hd__o21bai_1 _15527_ (.A1(_13665_),
    .A2(_13451_),
    .B1_N(_13985_),
    .Y(_14053_));
 sky130_fd_sc_hd__a21oi_1 _15528_ (.A1(_14009_),
    .A2(_14053_),
    .B1(_13706_),
    .Y(_14054_));
 sky130_fd_sc_hd__or2_1 _15529_ (.A(_13664_),
    .B(_14054_),
    .X(_14055_));
 sky130_fd_sc_hd__and3_1 _15530_ (.A(_13542_),
    .B(_13604_),
    .C(_13721_),
    .X(_14056_));
 sky130_fd_sc_hd__a211o_1 _15531_ (.A1(_13517_),
    .A2(_13302_),
    .B1(_13941_),
    .C1(_14056_),
    .X(_14057_));
 sky130_fd_sc_hd__a21oi_1 _15532_ (.A1(_13319_),
    .A2(_14057_),
    .B1(_13572_),
    .Y(_14058_));
 sky130_fd_sc_hd__a31o_1 _15533_ (.A1(_13682_),
    .A2(_13665_),
    .A3(_13348_),
    .B1(_13597_),
    .X(_14059_));
 sky130_fd_sc_hd__a21o_1 _15534_ (.A1(_13564_),
    .A2(_14059_),
    .B1(_13442_),
    .X(_14060_));
 sky130_fd_sc_hd__o21ai_1 _15535_ (.A1(_13398_),
    .A2(_13546_),
    .B1(_13872_),
    .Y(_14061_));
 sky130_fd_sc_hd__o21ai_1 _15536_ (.A1(_13512_),
    .A2(_13965_),
    .B1(_13823_),
    .Y(_14062_));
 sky130_fd_sc_hd__o211ai_1 _15537_ (.A1(_13512_),
    .A2(_14061_),
    .B1(_14062_),
    .C1(_13319_),
    .Y(_14063_));
 sky130_fd_sc_hd__or3_1 _15538_ (.A(_13422_),
    .B(_13531_),
    .C(_13616_),
    .X(_14064_));
 sky130_fd_sc_hd__a221o_1 _15539_ (.A1(_13665_),
    .A2(_13294_),
    .B1(_13559_),
    .B2(_13689_),
    .C1(_13483_),
    .X(_14065_));
 sky130_fd_sc_hd__a21oi_1 _15540_ (.A1(_13403_),
    .A2(_13689_),
    .B1(_13747_),
    .Y(_14066_));
 sky130_fd_sc_hd__o21a_1 _15541_ (.A1(_13341_),
    .A2(_13510_),
    .B1(_13744_),
    .X(_14067_));
 sky130_fd_sc_hd__o22a_1 _15542_ (.A1(_13374_),
    .A2(_14066_),
    .B1(_14067_),
    .B2(_13513_),
    .X(_14068_));
 sky130_fd_sc_hd__a31o_1 _15543_ (.A1(_14064_),
    .A2(_14065_),
    .A3(_14068_),
    .B1(_13466_),
    .X(_14069_));
 sky130_fd_sc_hd__o32a_1 _15544_ (.A1(_13767_),
    .A2(_13488_),
    .A3(_13401_),
    .B1(_13477_),
    .B2(_13672_),
    .X(_14070_));
 sky130_fd_sc_hd__a21o_1 _15545_ (.A1(_13649_),
    .A2(_14070_),
    .B1(_13442_),
    .X(_14071_));
 sky130_fd_sc_hd__and4_1 _15546_ (.A(_13638_),
    .B(_14063_),
    .C(_14069_),
    .D(_14071_),
    .X(_14072_));
 sky130_fd_sc_hd__a31oi_4 _15547_ (.A1(_14055_),
    .A2(_14058_),
    .A3(_14060_),
    .B1(_14072_),
    .Y(net28));
 sky130_fd_sc_hd__nor2_1 _15548_ (.A(_13501_),
    .B(_14029_),
    .Y(_14073_));
 sky130_fd_sc_hd__o22a_1 _15549_ (.A1(_13762_),
    .A2(_13878_),
    .B1(_14073_),
    .B2(_13572_),
    .X(net27));
 sky130_fd_sc_hd__nand2_1 _15550_ (.A(_13823_),
    .B(_13435_),
    .Y(_14074_));
 sky130_fd_sc_hd__a31o_1 _15551_ (.A1(_13760_),
    .A2(_13420_),
    .A3(_14074_),
    .B1(_13458_),
    .X(_14075_));
 sky130_fd_sc_hd__a21oi_1 _15552_ (.A1(_13467_),
    .A2(_13462_),
    .B1(_13878_),
    .Y(_14076_));
 sky130_fd_sc_hd__o22a_1 _15553_ (.A1(_13378_),
    .A2(_13767_),
    .B1(_13780_),
    .B2(_13398_),
    .X(_14077_));
 sky130_fd_sc_hd__a21o_1 _15554_ (.A1(_13455_),
    .A2(_14077_),
    .B1(_13442_),
    .X(_14078_));
 sky130_fd_sc_hd__a31o_1 _15555_ (.A1(_13431_),
    .A2(_13559_),
    .A3(_13780_),
    .B1(_13531_),
    .X(_14079_));
 sky130_fd_sc_hd__a21oi_1 _15556_ (.A1(_13363_),
    .A2(_13575_),
    .B1(_13483_),
    .Y(_14080_));
 sky130_fd_sc_hd__a21oi_1 _15557_ (.A1(_13496_),
    .A2(_14079_),
    .B1(_14080_),
    .Y(_14081_));
 sky130_fd_sc_hd__and3_1 _15558_ (.A(_13291_),
    .B(_13414_),
    .C(_13294_),
    .X(_14082_));
 sky130_fd_sc_hd__o32a_1 _15559_ (.A1(_13301_),
    .A2(_13767_),
    .A3(_13481_),
    .B1(_13797_),
    .B2(_14082_),
    .X(_14083_));
 sky130_fd_sc_hd__o22a_1 _15560_ (.A1(_13419_),
    .A2(_13370_),
    .B1(_13301_),
    .B2(_13336_),
    .X(_14084_));
 sky130_fd_sc_hd__a211o_1 _15561_ (.A1(_13398_),
    .A2(_13767_),
    .B1(_13458_),
    .C1(_13378_),
    .X(_14085_));
 sky130_fd_sc_hd__o221a_1 _15562_ (.A1(_13441_),
    .A2(_14083_),
    .B1(_14084_),
    .B2(_13366_),
    .C1(_14085_),
    .X(_14086_));
 sky130_fd_sc_hd__o211a_1 _15563_ (.A1(_13466_),
    .A2(_14081_),
    .B1(_14086_),
    .C1(_13904_),
    .X(_14087_));
 sky130_fd_sc_hd__a31oi_2 _15564_ (.A1(_14075_),
    .A2(_14076_),
    .A3(_14078_),
    .B1(_14087_),
    .Y(net24));
 sky130_fd_sc_hd__or3_1 _15565_ (.A(_13573_),
    .B(_13796_),
    .C(_13499_),
    .X(_14088_));
 sky130_fd_sc_hd__buf_1 _15566_ (.A(_14088_),
    .X(net13));
 sky130_fd_sc_hd__or3b_2 _15567_ (.A(_13174_),
    .B(\rvcpu.dp.plmw.RdW[3] ),
    .C_N(_13176_),
    .X(_14089_));
 sky130_fd_sc_hd__nand3_4 _15568_ (.A(\rvcpu.dp.plmw.RegWriteW ),
    .B(\rvcpu.dp.plmw.RdW[0] ),
    .C(\rvcpu.dp.plmw.RdW[1] ),
    .Y(_14090_));
 sky130_fd_sc_hd__nor2_2 _15569_ (.A(_14089_),
    .B(_14090_),
    .Y(_14091_));
 sky130_fd_sc_hd__buf_4 _15570_ (.A(_14091_),
    .X(_14092_));
 sky130_fd_sc_hd__mux2_1 _15571_ (.A0(\rvcpu.dp.rf.reg_file_arr[19][31] ),
    .A1(_13173_),
    .S(_14092_),
    .X(_14093_));
 sky130_fd_sc_hd__clkbuf_1 _15572_ (.A(_14093_),
    .X(_02219_));
 sky130_fd_sc_hd__mux2_1 _15573_ (.A0(\rvcpu.dp.rf.reg_file_arr[19][30] ),
    .A1(_13184_),
    .S(_14092_),
    .X(_14094_));
 sky130_fd_sc_hd__clkbuf_1 _15574_ (.A(_14094_),
    .X(_02218_));
 sky130_fd_sc_hd__mux2_1 _15575_ (.A0(\rvcpu.dp.rf.reg_file_arr[19][29] ),
    .A1(_13187_),
    .S(_14092_),
    .X(_14095_));
 sky130_fd_sc_hd__clkbuf_1 _15576_ (.A(_14095_),
    .X(_02217_));
 sky130_fd_sc_hd__mux2_1 _15577_ (.A0(\rvcpu.dp.rf.reg_file_arr[19][28] ),
    .A1(_13190_),
    .S(_14092_),
    .X(_14096_));
 sky130_fd_sc_hd__clkbuf_1 _15578_ (.A(_14096_),
    .X(_02216_));
 sky130_fd_sc_hd__mux2_1 _15579_ (.A0(\rvcpu.dp.rf.reg_file_arr[19][27] ),
    .A1(_13195_),
    .S(_14092_),
    .X(_14097_));
 sky130_fd_sc_hd__clkbuf_1 _15580_ (.A(_14097_),
    .X(_02215_));
 sky130_fd_sc_hd__mux2_1 _15581_ (.A0(\rvcpu.dp.rf.reg_file_arr[19][26] ),
    .A1(_13198_),
    .S(_14092_),
    .X(_14098_));
 sky130_fd_sc_hd__clkbuf_1 _15582_ (.A(_14098_),
    .X(_02214_));
 sky130_fd_sc_hd__mux2_1 _15583_ (.A0(\rvcpu.dp.rf.reg_file_arr[19][25] ),
    .A1(_13201_),
    .S(_14092_),
    .X(_14099_));
 sky130_fd_sc_hd__clkbuf_1 _15584_ (.A(_14099_),
    .X(_02213_));
 sky130_fd_sc_hd__mux2_1 _15585_ (.A0(\rvcpu.dp.rf.reg_file_arr[19][24] ),
    .A1(_13204_),
    .S(_14092_),
    .X(_14100_));
 sky130_fd_sc_hd__clkbuf_1 _15586_ (.A(_14100_),
    .X(_02212_));
 sky130_fd_sc_hd__mux2_1 _15587_ (.A0(\rvcpu.dp.rf.reg_file_arr[19][23] ),
    .A1(_13207_),
    .S(_14092_),
    .X(_14101_));
 sky130_fd_sc_hd__clkbuf_1 _15588_ (.A(_14101_),
    .X(_02211_));
 sky130_fd_sc_hd__mux2_1 _15589_ (.A0(\rvcpu.dp.rf.reg_file_arr[19][22] ),
    .A1(_13210_),
    .S(_14092_),
    .X(_14102_));
 sky130_fd_sc_hd__clkbuf_1 _15590_ (.A(_14102_),
    .X(_02210_));
 sky130_fd_sc_hd__clkbuf_4 _15591_ (.A(_14091_),
    .X(_14103_));
 sky130_fd_sc_hd__mux2_1 _15592_ (.A0(\rvcpu.dp.rf.reg_file_arr[19][21] ),
    .A1(_13213_),
    .S(_14103_),
    .X(_14104_));
 sky130_fd_sc_hd__clkbuf_1 _15593_ (.A(_14104_),
    .X(_02209_));
 sky130_fd_sc_hd__mux2_1 _15594_ (.A0(\rvcpu.dp.rf.reg_file_arr[19][20] ),
    .A1(_13217_),
    .S(_14103_),
    .X(_14105_));
 sky130_fd_sc_hd__clkbuf_1 _15595_ (.A(_14105_),
    .X(_02208_));
 sky130_fd_sc_hd__mux2_1 _15596_ (.A0(\rvcpu.dp.rf.reg_file_arr[19][19] ),
    .A1(_13220_),
    .S(_14103_),
    .X(_14106_));
 sky130_fd_sc_hd__clkbuf_1 _15597_ (.A(_14106_),
    .X(_02207_));
 sky130_fd_sc_hd__mux2_1 _15598_ (.A0(\rvcpu.dp.rf.reg_file_arr[19][18] ),
    .A1(_13223_),
    .S(_14103_),
    .X(_14107_));
 sky130_fd_sc_hd__clkbuf_1 _15599_ (.A(_14107_),
    .X(_02206_));
 sky130_fd_sc_hd__mux2_1 _15600_ (.A0(\rvcpu.dp.rf.reg_file_arr[19][17] ),
    .A1(_13226_),
    .S(_14103_),
    .X(_14108_));
 sky130_fd_sc_hd__clkbuf_1 _15601_ (.A(_14108_),
    .X(_02205_));
 sky130_fd_sc_hd__mux2_1 _15602_ (.A0(\rvcpu.dp.rf.reg_file_arr[19][16] ),
    .A1(_13229_),
    .S(_14103_),
    .X(_14109_));
 sky130_fd_sc_hd__clkbuf_1 _15603_ (.A(_14109_),
    .X(_02204_));
 sky130_fd_sc_hd__mux2_1 _15604_ (.A0(\rvcpu.dp.rf.reg_file_arr[19][15] ),
    .A1(_13232_),
    .S(_14103_),
    .X(_14110_));
 sky130_fd_sc_hd__clkbuf_1 _15605_ (.A(_14110_),
    .X(_02203_));
 sky130_fd_sc_hd__mux2_1 _15606_ (.A0(\rvcpu.dp.rf.reg_file_arr[19][14] ),
    .A1(_13235_),
    .S(_14103_),
    .X(_14111_));
 sky130_fd_sc_hd__clkbuf_1 _15607_ (.A(_14111_),
    .X(_02202_));
 sky130_fd_sc_hd__mux2_1 _15608_ (.A0(\rvcpu.dp.rf.reg_file_arr[19][13] ),
    .A1(_13238_),
    .S(_14103_),
    .X(_14112_));
 sky130_fd_sc_hd__clkbuf_1 _15609_ (.A(_14112_),
    .X(_02201_));
 sky130_fd_sc_hd__mux2_1 _15610_ (.A0(\rvcpu.dp.rf.reg_file_arr[19][12] ),
    .A1(_13241_),
    .S(_14103_),
    .X(_14113_));
 sky130_fd_sc_hd__clkbuf_1 _15611_ (.A(_14113_),
    .X(_02200_));
 sky130_fd_sc_hd__buf_4 _15612_ (.A(_14091_),
    .X(_14114_));
 sky130_fd_sc_hd__mux2_1 _15613_ (.A0(\rvcpu.dp.rf.reg_file_arr[19][11] ),
    .A1(_13244_),
    .S(_14114_),
    .X(_14115_));
 sky130_fd_sc_hd__clkbuf_1 _15614_ (.A(_14115_),
    .X(_02199_));
 sky130_fd_sc_hd__mux2_1 _15615_ (.A0(\rvcpu.dp.rf.reg_file_arr[19][10] ),
    .A1(_13248_),
    .S(_14114_),
    .X(_14116_));
 sky130_fd_sc_hd__clkbuf_1 _15616_ (.A(_14116_),
    .X(_02198_));
 sky130_fd_sc_hd__mux2_1 _15617_ (.A0(\rvcpu.dp.rf.reg_file_arr[19][9] ),
    .A1(_13251_),
    .S(_14114_),
    .X(_14117_));
 sky130_fd_sc_hd__clkbuf_1 _15618_ (.A(_14117_),
    .X(_02197_));
 sky130_fd_sc_hd__mux2_1 _15619_ (.A0(\rvcpu.dp.rf.reg_file_arr[19][8] ),
    .A1(_13254_),
    .S(_14114_),
    .X(_14118_));
 sky130_fd_sc_hd__clkbuf_1 _15620_ (.A(_14118_),
    .X(_02196_));
 sky130_fd_sc_hd__mux2_1 _15621_ (.A0(\rvcpu.dp.rf.reg_file_arr[19][7] ),
    .A1(_13257_),
    .S(_14114_),
    .X(_14119_));
 sky130_fd_sc_hd__clkbuf_1 _15622_ (.A(_14119_),
    .X(_02195_));
 sky130_fd_sc_hd__mux2_1 _15623_ (.A0(\rvcpu.dp.rf.reg_file_arr[19][6] ),
    .A1(_13260_),
    .S(_14114_),
    .X(_14120_));
 sky130_fd_sc_hd__clkbuf_1 _15624_ (.A(_14120_),
    .X(_02194_));
 sky130_fd_sc_hd__mux2_1 _15625_ (.A0(\rvcpu.dp.rf.reg_file_arr[19][5] ),
    .A1(_13263_),
    .S(_14114_),
    .X(_14121_));
 sky130_fd_sc_hd__clkbuf_1 _15626_ (.A(_14121_),
    .X(_02193_));
 sky130_fd_sc_hd__mux2_1 _15627_ (.A0(\rvcpu.dp.rf.reg_file_arr[19][4] ),
    .A1(_13266_),
    .S(_14114_),
    .X(_14122_));
 sky130_fd_sc_hd__clkbuf_1 _15628_ (.A(_14122_),
    .X(_02192_));
 sky130_fd_sc_hd__mux2_1 _15629_ (.A0(\rvcpu.dp.rf.reg_file_arr[19][3] ),
    .A1(_13269_),
    .S(_14114_),
    .X(_14123_));
 sky130_fd_sc_hd__clkbuf_1 _15630_ (.A(_14123_),
    .X(_02191_));
 sky130_fd_sc_hd__mux2_1 _15631_ (.A0(\rvcpu.dp.rf.reg_file_arr[19][2] ),
    .A1(_13272_),
    .S(_14114_),
    .X(_14124_));
 sky130_fd_sc_hd__clkbuf_1 _15632_ (.A(_14124_),
    .X(_02190_));
 sky130_fd_sc_hd__mux2_1 _15633_ (.A0(\rvcpu.dp.rf.reg_file_arr[19][1] ),
    .A1(_13275_),
    .S(_14091_),
    .X(_14125_));
 sky130_fd_sc_hd__clkbuf_1 _15634_ (.A(_14125_),
    .X(_02189_));
 sky130_fd_sc_hd__mux2_1 _15635_ (.A0(\rvcpu.dp.rf.reg_file_arr[19][0] ),
    .A1(_13278_),
    .S(_14091_),
    .X(_14126_));
 sky130_fd_sc_hd__clkbuf_1 _15636_ (.A(_14126_),
    .X(_02188_));
 sky130_fd_sc_hd__buf_4 _15637_ (.A(_13172_),
    .X(_14127_));
 sky130_fd_sc_hd__nor2_4 _15638_ (.A(\rvcpu.dp.plmw.RdW[1] ),
    .B(_13178_),
    .Y(_14128_));
 sky130_fd_sc_hd__and3_2 _15639_ (.A(_13174_),
    .B(\rvcpu.dp.plmw.RdW[3] ),
    .C(_13176_),
    .X(_14129_));
 sky130_fd_sc_hd__nand2_2 _15640_ (.A(_14128_),
    .B(_14129_),
    .Y(_14130_));
 sky130_fd_sc_hd__clkbuf_4 _15641_ (.A(_14130_),
    .X(_14131_));
 sky130_fd_sc_hd__mux2_1 _15642_ (.A0(_14127_),
    .A1(\rvcpu.dp.rf.reg_file_arr[29][31] ),
    .S(_14131_),
    .X(_14132_));
 sky130_fd_sc_hd__clkbuf_1 _15643_ (.A(_14132_),
    .X(_02187_));
 sky130_fd_sc_hd__buf_4 _15644_ (.A(_13183_),
    .X(_14133_));
 sky130_fd_sc_hd__mux2_1 _15645_ (.A0(_14133_),
    .A1(\rvcpu.dp.rf.reg_file_arr[29][30] ),
    .S(_14131_),
    .X(_14134_));
 sky130_fd_sc_hd__clkbuf_1 _15646_ (.A(_14134_),
    .X(_02186_));
 sky130_fd_sc_hd__buf_4 _15647_ (.A(_13186_),
    .X(_14135_));
 sky130_fd_sc_hd__mux2_1 _15648_ (.A0(_14135_),
    .A1(\rvcpu.dp.rf.reg_file_arr[29][29] ),
    .S(_14131_),
    .X(_14136_));
 sky130_fd_sc_hd__clkbuf_1 _15649_ (.A(_14136_),
    .X(_02185_));
 sky130_fd_sc_hd__buf_4 _15650_ (.A(_13189_),
    .X(_14137_));
 sky130_fd_sc_hd__mux2_1 _15651_ (.A0(_14137_),
    .A1(\rvcpu.dp.rf.reg_file_arr[29][28] ),
    .S(_14131_),
    .X(_14138_));
 sky130_fd_sc_hd__clkbuf_1 _15652_ (.A(_14138_),
    .X(_02184_));
 sky130_fd_sc_hd__buf_4 _15653_ (.A(_13194_),
    .X(_14139_));
 sky130_fd_sc_hd__mux2_1 _15654_ (.A0(_14139_),
    .A1(\rvcpu.dp.rf.reg_file_arr[29][27] ),
    .S(_14131_),
    .X(_14140_));
 sky130_fd_sc_hd__clkbuf_1 _15655_ (.A(_14140_),
    .X(_02183_));
 sky130_fd_sc_hd__buf_4 _15656_ (.A(_13197_),
    .X(_14141_));
 sky130_fd_sc_hd__mux2_1 _15657_ (.A0(_14141_),
    .A1(\rvcpu.dp.rf.reg_file_arr[29][26] ),
    .S(_14131_),
    .X(_14142_));
 sky130_fd_sc_hd__clkbuf_1 _15658_ (.A(_14142_),
    .X(_02182_));
 sky130_fd_sc_hd__clkbuf_8 _15659_ (.A(_13200_),
    .X(_14143_));
 sky130_fd_sc_hd__mux2_1 _15660_ (.A0(_14143_),
    .A1(\rvcpu.dp.rf.reg_file_arr[29][25] ),
    .S(_14131_),
    .X(_14144_));
 sky130_fd_sc_hd__clkbuf_1 _15661_ (.A(_14144_),
    .X(_02181_));
 sky130_fd_sc_hd__buf_4 _15662_ (.A(_13203_),
    .X(_14145_));
 sky130_fd_sc_hd__mux2_1 _15663_ (.A0(_14145_),
    .A1(\rvcpu.dp.rf.reg_file_arr[29][24] ),
    .S(_14131_),
    .X(_14146_));
 sky130_fd_sc_hd__clkbuf_1 _15664_ (.A(_14146_),
    .X(_02180_));
 sky130_fd_sc_hd__clkbuf_8 _15665_ (.A(_13206_),
    .X(_14147_));
 sky130_fd_sc_hd__mux2_1 _15666_ (.A0(_14147_),
    .A1(\rvcpu.dp.rf.reg_file_arr[29][23] ),
    .S(_14131_),
    .X(_14148_));
 sky130_fd_sc_hd__clkbuf_1 _15667_ (.A(_14148_),
    .X(_02179_));
 sky130_fd_sc_hd__buf_4 _15668_ (.A(_13209_),
    .X(_14149_));
 sky130_fd_sc_hd__mux2_1 _15669_ (.A0(_14149_),
    .A1(\rvcpu.dp.rf.reg_file_arr[29][22] ),
    .S(_14131_),
    .X(_14150_));
 sky130_fd_sc_hd__clkbuf_1 _15670_ (.A(_14150_),
    .X(_02178_));
 sky130_fd_sc_hd__buf_4 _15671_ (.A(_13212_),
    .X(_14151_));
 sky130_fd_sc_hd__clkbuf_4 _15672_ (.A(_14130_),
    .X(_14152_));
 sky130_fd_sc_hd__mux2_1 _15673_ (.A0(_14151_),
    .A1(\rvcpu.dp.rf.reg_file_arr[29][21] ),
    .S(_14152_),
    .X(_14153_));
 sky130_fd_sc_hd__clkbuf_1 _15674_ (.A(_14153_),
    .X(_02177_));
 sky130_fd_sc_hd__buf_4 _15675_ (.A(_13216_),
    .X(_14154_));
 sky130_fd_sc_hd__mux2_1 _15676_ (.A0(_14154_),
    .A1(\rvcpu.dp.rf.reg_file_arr[29][20] ),
    .S(_14152_),
    .X(_14155_));
 sky130_fd_sc_hd__clkbuf_1 _15677_ (.A(_14155_),
    .X(_02176_));
 sky130_fd_sc_hd__buf_4 _15678_ (.A(_13219_),
    .X(_14156_));
 sky130_fd_sc_hd__mux2_1 _15679_ (.A0(_14156_),
    .A1(\rvcpu.dp.rf.reg_file_arr[29][19] ),
    .S(_14152_),
    .X(_14157_));
 sky130_fd_sc_hd__clkbuf_1 _15680_ (.A(_14157_),
    .X(_02175_));
 sky130_fd_sc_hd__buf_4 _15681_ (.A(_13222_),
    .X(_14158_));
 sky130_fd_sc_hd__mux2_1 _15682_ (.A0(_14158_),
    .A1(\rvcpu.dp.rf.reg_file_arr[29][18] ),
    .S(_14152_),
    .X(_14159_));
 sky130_fd_sc_hd__clkbuf_1 _15683_ (.A(_14159_),
    .X(_02174_));
 sky130_fd_sc_hd__buf_4 _15684_ (.A(_13225_),
    .X(_14160_));
 sky130_fd_sc_hd__mux2_1 _15685_ (.A0(_14160_),
    .A1(\rvcpu.dp.rf.reg_file_arr[29][17] ),
    .S(_14152_),
    .X(_14161_));
 sky130_fd_sc_hd__clkbuf_1 _15686_ (.A(_14161_),
    .X(_02173_));
 sky130_fd_sc_hd__buf_4 _15687_ (.A(_13228_),
    .X(_14162_));
 sky130_fd_sc_hd__mux2_1 _15688_ (.A0(_14162_),
    .A1(\rvcpu.dp.rf.reg_file_arr[29][16] ),
    .S(_14152_),
    .X(_14163_));
 sky130_fd_sc_hd__clkbuf_1 _15689_ (.A(_14163_),
    .X(_02172_));
 sky130_fd_sc_hd__buf_4 _15690_ (.A(_13231_),
    .X(_14164_));
 sky130_fd_sc_hd__mux2_1 _15691_ (.A0(_14164_),
    .A1(\rvcpu.dp.rf.reg_file_arr[29][15] ),
    .S(_14152_),
    .X(_14165_));
 sky130_fd_sc_hd__clkbuf_1 _15692_ (.A(_14165_),
    .X(_02171_));
 sky130_fd_sc_hd__buf_4 _15693_ (.A(_13234_),
    .X(_14166_));
 sky130_fd_sc_hd__mux2_1 _15694_ (.A0(_14166_),
    .A1(\rvcpu.dp.rf.reg_file_arr[29][14] ),
    .S(_14152_),
    .X(_14167_));
 sky130_fd_sc_hd__clkbuf_1 _15695_ (.A(_14167_),
    .X(_02170_));
 sky130_fd_sc_hd__buf_4 _15696_ (.A(_13237_),
    .X(_14168_));
 sky130_fd_sc_hd__mux2_1 _15697_ (.A0(_14168_),
    .A1(\rvcpu.dp.rf.reg_file_arr[29][13] ),
    .S(_14152_),
    .X(_14169_));
 sky130_fd_sc_hd__clkbuf_1 _15698_ (.A(_14169_),
    .X(_02169_));
 sky130_fd_sc_hd__buf_4 _15699_ (.A(_13240_),
    .X(_14170_));
 sky130_fd_sc_hd__mux2_1 _15700_ (.A0(_14170_),
    .A1(\rvcpu.dp.rf.reg_file_arr[29][12] ),
    .S(_14152_),
    .X(_14171_));
 sky130_fd_sc_hd__clkbuf_1 _15701_ (.A(_14171_),
    .X(_02168_));
 sky130_fd_sc_hd__buf_4 _15702_ (.A(_13243_),
    .X(_14172_));
 sky130_fd_sc_hd__buf_4 _15703_ (.A(_14130_),
    .X(_14173_));
 sky130_fd_sc_hd__mux2_1 _15704_ (.A0(_14172_),
    .A1(\rvcpu.dp.rf.reg_file_arr[29][11] ),
    .S(_14173_),
    .X(_14174_));
 sky130_fd_sc_hd__clkbuf_1 _15705_ (.A(_14174_),
    .X(_02167_));
 sky130_fd_sc_hd__buf_4 _15706_ (.A(_13247_),
    .X(_14175_));
 sky130_fd_sc_hd__mux2_1 _15707_ (.A0(_14175_),
    .A1(\rvcpu.dp.rf.reg_file_arr[29][10] ),
    .S(_14173_),
    .X(_14176_));
 sky130_fd_sc_hd__clkbuf_1 _15708_ (.A(_14176_),
    .X(_02166_));
 sky130_fd_sc_hd__buf_4 _15709_ (.A(_13250_),
    .X(_14177_));
 sky130_fd_sc_hd__mux2_1 _15710_ (.A0(_14177_),
    .A1(\rvcpu.dp.rf.reg_file_arr[29][9] ),
    .S(_14173_),
    .X(_14178_));
 sky130_fd_sc_hd__clkbuf_1 _15711_ (.A(_14178_),
    .X(_02165_));
 sky130_fd_sc_hd__buf_4 _15712_ (.A(_13253_),
    .X(_14179_));
 sky130_fd_sc_hd__mux2_1 _15713_ (.A0(_14179_),
    .A1(\rvcpu.dp.rf.reg_file_arr[29][8] ),
    .S(_14173_),
    .X(_14180_));
 sky130_fd_sc_hd__clkbuf_1 _15714_ (.A(_14180_),
    .X(_02164_));
 sky130_fd_sc_hd__buf_4 _15715_ (.A(_13256_),
    .X(_14181_));
 sky130_fd_sc_hd__mux2_1 _15716_ (.A0(_14181_),
    .A1(\rvcpu.dp.rf.reg_file_arr[29][7] ),
    .S(_14173_),
    .X(_14182_));
 sky130_fd_sc_hd__clkbuf_1 _15717_ (.A(_14182_),
    .X(_02163_));
 sky130_fd_sc_hd__clkbuf_8 _15718_ (.A(_13259_),
    .X(_14183_));
 sky130_fd_sc_hd__mux2_1 _15719_ (.A0(_14183_),
    .A1(\rvcpu.dp.rf.reg_file_arr[29][6] ),
    .S(_14173_),
    .X(_14184_));
 sky130_fd_sc_hd__clkbuf_1 _15720_ (.A(_14184_),
    .X(_02162_));
 sky130_fd_sc_hd__buf_4 _15721_ (.A(_13262_),
    .X(_14185_));
 sky130_fd_sc_hd__mux2_1 _15722_ (.A0(_14185_),
    .A1(\rvcpu.dp.rf.reg_file_arr[29][5] ),
    .S(_14173_),
    .X(_14186_));
 sky130_fd_sc_hd__clkbuf_1 _15723_ (.A(_14186_),
    .X(_02161_));
 sky130_fd_sc_hd__clkbuf_8 _15724_ (.A(_13265_),
    .X(_14187_));
 sky130_fd_sc_hd__mux2_1 _15725_ (.A0(_14187_),
    .A1(\rvcpu.dp.rf.reg_file_arr[29][4] ),
    .S(_14173_),
    .X(_14188_));
 sky130_fd_sc_hd__clkbuf_1 _15726_ (.A(_14188_),
    .X(_02160_));
 sky130_fd_sc_hd__buf_4 _15727_ (.A(_13268_),
    .X(_14189_));
 sky130_fd_sc_hd__mux2_1 _15728_ (.A0(_14189_),
    .A1(\rvcpu.dp.rf.reg_file_arr[29][3] ),
    .S(_14173_),
    .X(_14190_));
 sky130_fd_sc_hd__clkbuf_1 _15729_ (.A(_14190_),
    .X(_02159_));
 sky130_fd_sc_hd__buf_4 _15730_ (.A(_13271_),
    .X(_14191_));
 sky130_fd_sc_hd__mux2_1 _15731_ (.A0(_14191_),
    .A1(\rvcpu.dp.rf.reg_file_arr[29][2] ),
    .S(_14173_),
    .X(_14192_));
 sky130_fd_sc_hd__clkbuf_1 _15732_ (.A(_14192_),
    .X(_02158_));
 sky130_fd_sc_hd__buf_4 _15733_ (.A(_13274_),
    .X(_14193_));
 sky130_fd_sc_hd__mux2_1 _15734_ (.A0(_14193_),
    .A1(\rvcpu.dp.rf.reg_file_arr[29][1] ),
    .S(_14130_),
    .X(_14194_));
 sky130_fd_sc_hd__clkbuf_1 _15735_ (.A(_14194_),
    .X(_02157_));
 sky130_fd_sc_hd__buf_4 _15736_ (.A(_13277_),
    .X(_14195_));
 sky130_fd_sc_hd__mux2_1 _15737_ (.A0(_14195_),
    .A1(\rvcpu.dp.rf.reg_file_arr[29][0] ),
    .S(_14130_),
    .X(_14196_));
 sky130_fd_sc_hd__clkbuf_1 _15738_ (.A(_14196_),
    .X(_02156_));
 sky130_fd_sc_hd__and3_4 _15739_ (.A(\rvcpu.dp.plmw.RegWriteW ),
    .B(\rvcpu.dp.plmw.RdW[0] ),
    .C(\rvcpu.dp.plmw.RdW[1] ),
    .X(_14197_));
 sky130_fd_sc_hd__nand2_2 _15740_ (.A(_14197_),
    .B(_14129_),
    .Y(_14198_));
 sky130_fd_sc_hd__clkbuf_4 _15741_ (.A(_14198_),
    .X(_14199_));
 sky130_fd_sc_hd__mux2_1 _15742_ (.A0(_14127_),
    .A1(\rvcpu.dp.rf.reg_file_arr[31][31] ),
    .S(_14199_),
    .X(_14200_));
 sky130_fd_sc_hd__clkbuf_1 _15743_ (.A(_14200_),
    .X(_02155_));
 sky130_fd_sc_hd__mux2_1 _15744_ (.A0(_14133_),
    .A1(\rvcpu.dp.rf.reg_file_arr[31][30] ),
    .S(_14199_),
    .X(_14201_));
 sky130_fd_sc_hd__clkbuf_1 _15745_ (.A(_14201_),
    .X(_02154_));
 sky130_fd_sc_hd__mux2_1 _15746_ (.A0(_14135_),
    .A1(\rvcpu.dp.rf.reg_file_arr[31][29] ),
    .S(_14199_),
    .X(_14202_));
 sky130_fd_sc_hd__clkbuf_1 _15747_ (.A(_14202_),
    .X(_02153_));
 sky130_fd_sc_hd__mux2_1 _15748_ (.A0(_14137_),
    .A1(\rvcpu.dp.rf.reg_file_arr[31][28] ),
    .S(_14199_),
    .X(_14203_));
 sky130_fd_sc_hd__clkbuf_1 _15749_ (.A(_14203_),
    .X(_02152_));
 sky130_fd_sc_hd__mux2_1 _15750_ (.A0(_14139_),
    .A1(\rvcpu.dp.rf.reg_file_arr[31][27] ),
    .S(_14199_),
    .X(_14204_));
 sky130_fd_sc_hd__clkbuf_1 _15751_ (.A(_14204_),
    .X(_02151_));
 sky130_fd_sc_hd__mux2_1 _15752_ (.A0(_14141_),
    .A1(\rvcpu.dp.rf.reg_file_arr[31][26] ),
    .S(_14199_),
    .X(_14205_));
 sky130_fd_sc_hd__clkbuf_1 _15753_ (.A(_14205_),
    .X(_02150_));
 sky130_fd_sc_hd__mux2_1 _15754_ (.A0(_14143_),
    .A1(\rvcpu.dp.rf.reg_file_arr[31][25] ),
    .S(_14199_),
    .X(_14206_));
 sky130_fd_sc_hd__clkbuf_1 _15755_ (.A(_14206_),
    .X(_02149_));
 sky130_fd_sc_hd__mux2_1 _15756_ (.A0(_14145_),
    .A1(\rvcpu.dp.rf.reg_file_arr[31][24] ),
    .S(_14199_),
    .X(_14207_));
 sky130_fd_sc_hd__clkbuf_1 _15757_ (.A(_14207_),
    .X(_02148_));
 sky130_fd_sc_hd__mux2_1 _15758_ (.A0(_14147_),
    .A1(\rvcpu.dp.rf.reg_file_arr[31][23] ),
    .S(_14199_),
    .X(_14208_));
 sky130_fd_sc_hd__clkbuf_1 _15759_ (.A(_14208_),
    .X(_02147_));
 sky130_fd_sc_hd__mux2_1 _15760_ (.A0(_14149_),
    .A1(\rvcpu.dp.rf.reg_file_arr[31][22] ),
    .S(_14199_),
    .X(_14209_));
 sky130_fd_sc_hd__clkbuf_1 _15761_ (.A(_14209_),
    .X(_02146_));
 sky130_fd_sc_hd__clkbuf_4 _15762_ (.A(_14198_),
    .X(_14210_));
 sky130_fd_sc_hd__mux2_1 _15763_ (.A0(_14151_),
    .A1(\rvcpu.dp.rf.reg_file_arr[31][21] ),
    .S(_14210_),
    .X(_14211_));
 sky130_fd_sc_hd__clkbuf_1 _15764_ (.A(_14211_),
    .X(_02145_));
 sky130_fd_sc_hd__mux2_1 _15765_ (.A0(_14154_),
    .A1(\rvcpu.dp.rf.reg_file_arr[31][20] ),
    .S(_14210_),
    .X(_14212_));
 sky130_fd_sc_hd__clkbuf_1 _15766_ (.A(_14212_),
    .X(_02144_));
 sky130_fd_sc_hd__mux2_1 _15767_ (.A0(_14156_),
    .A1(\rvcpu.dp.rf.reg_file_arr[31][19] ),
    .S(_14210_),
    .X(_14213_));
 sky130_fd_sc_hd__clkbuf_1 _15768_ (.A(_14213_),
    .X(_02143_));
 sky130_fd_sc_hd__mux2_1 _15769_ (.A0(_14158_),
    .A1(\rvcpu.dp.rf.reg_file_arr[31][18] ),
    .S(_14210_),
    .X(_14214_));
 sky130_fd_sc_hd__clkbuf_1 _15770_ (.A(_14214_),
    .X(_02142_));
 sky130_fd_sc_hd__mux2_1 _15771_ (.A0(_14160_),
    .A1(\rvcpu.dp.rf.reg_file_arr[31][17] ),
    .S(_14210_),
    .X(_14215_));
 sky130_fd_sc_hd__clkbuf_1 _15772_ (.A(_14215_),
    .X(_02141_));
 sky130_fd_sc_hd__mux2_1 _15773_ (.A0(_14162_),
    .A1(\rvcpu.dp.rf.reg_file_arr[31][16] ),
    .S(_14210_),
    .X(_14216_));
 sky130_fd_sc_hd__clkbuf_1 _15774_ (.A(_14216_),
    .X(_02140_));
 sky130_fd_sc_hd__mux2_1 _15775_ (.A0(_14164_),
    .A1(\rvcpu.dp.rf.reg_file_arr[31][15] ),
    .S(_14210_),
    .X(_14217_));
 sky130_fd_sc_hd__clkbuf_1 _15776_ (.A(_14217_),
    .X(_02139_));
 sky130_fd_sc_hd__mux2_1 _15777_ (.A0(_14166_),
    .A1(\rvcpu.dp.rf.reg_file_arr[31][14] ),
    .S(_14210_),
    .X(_14218_));
 sky130_fd_sc_hd__clkbuf_1 _15778_ (.A(_14218_),
    .X(_02138_));
 sky130_fd_sc_hd__mux2_1 _15779_ (.A0(_14168_),
    .A1(\rvcpu.dp.rf.reg_file_arr[31][13] ),
    .S(_14210_),
    .X(_14219_));
 sky130_fd_sc_hd__clkbuf_1 _15780_ (.A(_14219_),
    .X(_02137_));
 sky130_fd_sc_hd__mux2_1 _15781_ (.A0(_14170_),
    .A1(\rvcpu.dp.rf.reg_file_arr[31][12] ),
    .S(_14210_),
    .X(_14220_));
 sky130_fd_sc_hd__clkbuf_1 _15782_ (.A(_14220_),
    .X(_02136_));
 sky130_fd_sc_hd__buf_4 _15783_ (.A(_14198_),
    .X(_14221_));
 sky130_fd_sc_hd__mux2_1 _15784_ (.A0(_14172_),
    .A1(\rvcpu.dp.rf.reg_file_arr[31][11] ),
    .S(_14221_),
    .X(_14222_));
 sky130_fd_sc_hd__clkbuf_1 _15785_ (.A(_14222_),
    .X(_02135_));
 sky130_fd_sc_hd__mux2_1 _15786_ (.A0(_14175_),
    .A1(\rvcpu.dp.rf.reg_file_arr[31][10] ),
    .S(_14221_),
    .X(_14223_));
 sky130_fd_sc_hd__clkbuf_1 _15787_ (.A(_14223_),
    .X(_02134_));
 sky130_fd_sc_hd__mux2_1 _15788_ (.A0(_14177_),
    .A1(\rvcpu.dp.rf.reg_file_arr[31][9] ),
    .S(_14221_),
    .X(_14224_));
 sky130_fd_sc_hd__clkbuf_1 _15789_ (.A(_14224_),
    .X(_02133_));
 sky130_fd_sc_hd__mux2_1 _15790_ (.A0(_14179_),
    .A1(\rvcpu.dp.rf.reg_file_arr[31][8] ),
    .S(_14221_),
    .X(_14225_));
 sky130_fd_sc_hd__clkbuf_1 _15791_ (.A(_14225_),
    .X(_02132_));
 sky130_fd_sc_hd__mux2_1 _15792_ (.A0(_14181_),
    .A1(\rvcpu.dp.rf.reg_file_arr[31][7] ),
    .S(_14221_),
    .X(_14226_));
 sky130_fd_sc_hd__clkbuf_1 _15793_ (.A(_14226_),
    .X(_02131_));
 sky130_fd_sc_hd__mux2_1 _15794_ (.A0(_14183_),
    .A1(\rvcpu.dp.rf.reg_file_arr[31][6] ),
    .S(_14221_),
    .X(_14227_));
 sky130_fd_sc_hd__clkbuf_1 _15795_ (.A(_14227_),
    .X(_02130_));
 sky130_fd_sc_hd__mux2_1 _15796_ (.A0(_14185_),
    .A1(\rvcpu.dp.rf.reg_file_arr[31][5] ),
    .S(_14221_),
    .X(_14228_));
 sky130_fd_sc_hd__clkbuf_1 _15797_ (.A(_14228_),
    .X(_02129_));
 sky130_fd_sc_hd__mux2_1 _15798_ (.A0(_14187_),
    .A1(\rvcpu.dp.rf.reg_file_arr[31][4] ),
    .S(_14221_),
    .X(_14229_));
 sky130_fd_sc_hd__clkbuf_1 _15799_ (.A(_14229_),
    .X(_02128_));
 sky130_fd_sc_hd__mux2_1 _15800_ (.A0(_14189_),
    .A1(\rvcpu.dp.rf.reg_file_arr[31][3] ),
    .S(_14221_),
    .X(_14230_));
 sky130_fd_sc_hd__clkbuf_1 _15801_ (.A(_14230_),
    .X(_02127_));
 sky130_fd_sc_hd__mux2_1 _15802_ (.A0(_14191_),
    .A1(\rvcpu.dp.rf.reg_file_arr[31][2] ),
    .S(_14221_),
    .X(_14231_));
 sky130_fd_sc_hd__clkbuf_1 _15803_ (.A(_14231_),
    .X(_02126_));
 sky130_fd_sc_hd__mux2_1 _15804_ (.A0(_14193_),
    .A1(\rvcpu.dp.rf.reg_file_arr[31][1] ),
    .S(_14198_),
    .X(_14232_));
 sky130_fd_sc_hd__clkbuf_1 _15805_ (.A(_14232_),
    .X(_02125_));
 sky130_fd_sc_hd__mux2_1 _15806_ (.A0(_14195_),
    .A1(\rvcpu.dp.rf.reg_file_arr[31][0] ),
    .S(_14198_),
    .X(_14233_));
 sky130_fd_sc_hd__clkbuf_1 _15807_ (.A(_14233_),
    .X(_02124_));
 sky130_fd_sc_hd__or3_4 _15808_ (.A(_13174_),
    .B(\rvcpu.dp.plmw.RdW[3] ),
    .C(_13176_),
    .X(_14234_));
 sky130_fd_sc_hd__nor2_2 _15809_ (.A(_14090_),
    .B(_14234_),
    .Y(_14235_));
 sky130_fd_sc_hd__buf_4 _15810_ (.A(_14235_),
    .X(_14236_));
 sky130_fd_sc_hd__mux2_1 _15811_ (.A0(\rvcpu.dp.rf.reg_file_arr[3][31] ),
    .A1(_13173_),
    .S(_14236_),
    .X(_14237_));
 sky130_fd_sc_hd__clkbuf_1 _15812_ (.A(_14237_),
    .X(_02115_));
 sky130_fd_sc_hd__mux2_1 _15813_ (.A0(\rvcpu.dp.rf.reg_file_arr[3][30] ),
    .A1(_13184_),
    .S(_14236_),
    .X(_14238_));
 sky130_fd_sc_hd__clkbuf_1 _15814_ (.A(_14238_),
    .X(_02114_));
 sky130_fd_sc_hd__mux2_1 _15815_ (.A0(\rvcpu.dp.rf.reg_file_arr[3][29] ),
    .A1(_13187_),
    .S(_14236_),
    .X(_14239_));
 sky130_fd_sc_hd__clkbuf_1 _15816_ (.A(_14239_),
    .X(_02113_));
 sky130_fd_sc_hd__mux2_1 _15817_ (.A0(\rvcpu.dp.rf.reg_file_arr[3][28] ),
    .A1(_13190_),
    .S(_14236_),
    .X(_14240_));
 sky130_fd_sc_hd__clkbuf_1 _15818_ (.A(_14240_),
    .X(_02112_));
 sky130_fd_sc_hd__mux2_1 _15819_ (.A0(\rvcpu.dp.rf.reg_file_arr[3][27] ),
    .A1(_13195_),
    .S(_14236_),
    .X(_14241_));
 sky130_fd_sc_hd__clkbuf_1 _15820_ (.A(_14241_),
    .X(_02111_));
 sky130_fd_sc_hd__mux2_1 _15821_ (.A0(\rvcpu.dp.rf.reg_file_arr[3][26] ),
    .A1(_13198_),
    .S(_14236_),
    .X(_14242_));
 sky130_fd_sc_hd__clkbuf_1 _15822_ (.A(_14242_),
    .X(_02110_));
 sky130_fd_sc_hd__mux2_1 _15823_ (.A0(\rvcpu.dp.rf.reg_file_arr[3][25] ),
    .A1(_13201_),
    .S(_14236_),
    .X(_14243_));
 sky130_fd_sc_hd__clkbuf_1 _15824_ (.A(_14243_),
    .X(_02109_));
 sky130_fd_sc_hd__mux2_1 _15825_ (.A0(\rvcpu.dp.rf.reg_file_arr[3][24] ),
    .A1(_13204_),
    .S(_14236_),
    .X(_14244_));
 sky130_fd_sc_hd__clkbuf_1 _15826_ (.A(_14244_),
    .X(_02108_));
 sky130_fd_sc_hd__mux2_1 _15827_ (.A0(\rvcpu.dp.rf.reg_file_arr[3][23] ),
    .A1(_13207_),
    .S(_14236_),
    .X(_14245_));
 sky130_fd_sc_hd__clkbuf_1 _15828_ (.A(_14245_),
    .X(_02107_));
 sky130_fd_sc_hd__mux2_1 _15829_ (.A0(\rvcpu.dp.rf.reg_file_arr[3][22] ),
    .A1(_13210_),
    .S(_14236_),
    .X(_14246_));
 sky130_fd_sc_hd__clkbuf_1 _15830_ (.A(_14246_),
    .X(_02106_));
 sky130_fd_sc_hd__clkbuf_4 _15831_ (.A(_14235_),
    .X(_14247_));
 sky130_fd_sc_hd__mux2_1 _15832_ (.A0(\rvcpu.dp.rf.reg_file_arr[3][21] ),
    .A1(_13213_),
    .S(_14247_),
    .X(_14248_));
 sky130_fd_sc_hd__clkbuf_1 _15833_ (.A(_14248_),
    .X(_02105_));
 sky130_fd_sc_hd__mux2_1 _15834_ (.A0(\rvcpu.dp.rf.reg_file_arr[3][20] ),
    .A1(_13217_),
    .S(_14247_),
    .X(_14249_));
 sky130_fd_sc_hd__clkbuf_1 _15835_ (.A(_14249_),
    .X(_02104_));
 sky130_fd_sc_hd__mux2_1 _15836_ (.A0(\rvcpu.dp.rf.reg_file_arr[3][19] ),
    .A1(_13220_),
    .S(_14247_),
    .X(_14250_));
 sky130_fd_sc_hd__clkbuf_1 _15837_ (.A(_14250_),
    .X(_02103_));
 sky130_fd_sc_hd__mux2_1 _15838_ (.A0(\rvcpu.dp.rf.reg_file_arr[3][18] ),
    .A1(_13223_),
    .S(_14247_),
    .X(_14251_));
 sky130_fd_sc_hd__clkbuf_1 _15839_ (.A(_14251_),
    .X(_02102_));
 sky130_fd_sc_hd__mux2_1 _15840_ (.A0(\rvcpu.dp.rf.reg_file_arr[3][17] ),
    .A1(_13226_),
    .S(_14247_),
    .X(_14252_));
 sky130_fd_sc_hd__clkbuf_1 _15841_ (.A(_14252_),
    .X(_02101_));
 sky130_fd_sc_hd__mux2_1 _15842_ (.A0(\rvcpu.dp.rf.reg_file_arr[3][16] ),
    .A1(_13229_),
    .S(_14247_),
    .X(_14253_));
 sky130_fd_sc_hd__clkbuf_1 _15843_ (.A(_14253_),
    .X(_02100_));
 sky130_fd_sc_hd__mux2_1 _15844_ (.A0(\rvcpu.dp.rf.reg_file_arr[3][15] ),
    .A1(_13232_),
    .S(_14247_),
    .X(_14254_));
 sky130_fd_sc_hd__clkbuf_1 _15845_ (.A(_14254_),
    .X(_02099_));
 sky130_fd_sc_hd__mux2_1 _15846_ (.A0(\rvcpu.dp.rf.reg_file_arr[3][14] ),
    .A1(_13235_),
    .S(_14247_),
    .X(_14255_));
 sky130_fd_sc_hd__clkbuf_1 _15847_ (.A(_14255_),
    .X(_02098_));
 sky130_fd_sc_hd__mux2_1 _15848_ (.A0(\rvcpu.dp.rf.reg_file_arr[3][13] ),
    .A1(_13238_),
    .S(_14247_),
    .X(_14256_));
 sky130_fd_sc_hd__clkbuf_1 _15849_ (.A(_14256_),
    .X(_02097_));
 sky130_fd_sc_hd__mux2_1 _15850_ (.A0(\rvcpu.dp.rf.reg_file_arr[3][12] ),
    .A1(_13241_),
    .S(_14247_),
    .X(_14257_));
 sky130_fd_sc_hd__clkbuf_1 _15851_ (.A(_14257_),
    .X(_02096_));
 sky130_fd_sc_hd__buf_4 _15852_ (.A(_14235_),
    .X(_14258_));
 sky130_fd_sc_hd__mux2_1 _15853_ (.A0(\rvcpu.dp.rf.reg_file_arr[3][11] ),
    .A1(_13244_),
    .S(_14258_),
    .X(_14259_));
 sky130_fd_sc_hd__clkbuf_1 _15854_ (.A(_14259_),
    .X(_02095_));
 sky130_fd_sc_hd__mux2_1 _15855_ (.A0(\rvcpu.dp.rf.reg_file_arr[3][10] ),
    .A1(_13248_),
    .S(_14258_),
    .X(_14260_));
 sky130_fd_sc_hd__clkbuf_1 _15856_ (.A(_14260_),
    .X(_02094_));
 sky130_fd_sc_hd__mux2_1 _15857_ (.A0(\rvcpu.dp.rf.reg_file_arr[3][9] ),
    .A1(_13251_),
    .S(_14258_),
    .X(_14261_));
 sky130_fd_sc_hd__clkbuf_1 _15858_ (.A(_14261_),
    .X(_02093_));
 sky130_fd_sc_hd__mux2_1 _15859_ (.A0(\rvcpu.dp.rf.reg_file_arr[3][8] ),
    .A1(_13254_),
    .S(_14258_),
    .X(_14262_));
 sky130_fd_sc_hd__clkbuf_1 _15860_ (.A(_14262_),
    .X(_02092_));
 sky130_fd_sc_hd__mux2_1 _15861_ (.A0(\rvcpu.dp.rf.reg_file_arr[3][7] ),
    .A1(_13257_),
    .S(_14258_),
    .X(_14263_));
 sky130_fd_sc_hd__clkbuf_1 _15862_ (.A(_14263_),
    .X(_02091_));
 sky130_fd_sc_hd__mux2_1 _15863_ (.A0(\rvcpu.dp.rf.reg_file_arr[3][6] ),
    .A1(_13260_),
    .S(_14258_),
    .X(_14264_));
 sky130_fd_sc_hd__clkbuf_1 _15864_ (.A(_14264_),
    .X(_02090_));
 sky130_fd_sc_hd__mux2_1 _15865_ (.A0(\rvcpu.dp.rf.reg_file_arr[3][5] ),
    .A1(_13263_),
    .S(_14258_),
    .X(_14265_));
 sky130_fd_sc_hd__clkbuf_1 _15866_ (.A(_14265_),
    .X(_02089_));
 sky130_fd_sc_hd__mux2_1 _15867_ (.A0(\rvcpu.dp.rf.reg_file_arr[3][4] ),
    .A1(_13266_),
    .S(_14258_),
    .X(_14266_));
 sky130_fd_sc_hd__clkbuf_1 _15868_ (.A(_14266_),
    .X(_02088_));
 sky130_fd_sc_hd__mux2_1 _15869_ (.A0(\rvcpu.dp.rf.reg_file_arr[3][3] ),
    .A1(_13269_),
    .S(_14258_),
    .X(_14267_));
 sky130_fd_sc_hd__clkbuf_1 _15870_ (.A(_14267_),
    .X(_02087_));
 sky130_fd_sc_hd__mux2_1 _15871_ (.A0(\rvcpu.dp.rf.reg_file_arr[3][2] ),
    .A1(_13272_),
    .S(_14258_),
    .X(_14268_));
 sky130_fd_sc_hd__clkbuf_1 _15872_ (.A(_14268_),
    .X(_02086_));
 sky130_fd_sc_hd__mux2_1 _15873_ (.A0(\rvcpu.dp.rf.reg_file_arr[3][1] ),
    .A1(_13275_),
    .S(_14235_),
    .X(_14269_));
 sky130_fd_sc_hd__clkbuf_1 _15874_ (.A(_14269_),
    .X(_02085_));
 sky130_fd_sc_hd__mux2_1 _15875_ (.A0(\rvcpu.dp.rf.reg_file_arr[3][0] ),
    .A1(_13278_),
    .S(_14235_),
    .X(_14270_));
 sky130_fd_sc_hd__clkbuf_1 _15876_ (.A(_14270_),
    .X(_02084_));
 sky130_fd_sc_hd__or3b_4 _15877_ (.A(\rvcpu.dp.plmw.RdW[3] ),
    .B(_13176_),
    .C_N(_13174_),
    .X(_14271_));
 sky130_fd_sc_hd__or3b_1 _15878_ (.A(\rvcpu.dp.plmw.RdW[0] ),
    .B(\rvcpu.dp.plmw.RdW[1] ),
    .C_N(\rvcpu.dp.plmw.RegWriteW ),
    .X(_14272_));
 sky130_fd_sc_hd__buf_4 _15879_ (.A(_14272_),
    .X(_14273_));
 sky130_fd_sc_hd__nor2_2 _15880_ (.A(_14271_),
    .B(_14273_),
    .Y(_14274_));
 sky130_fd_sc_hd__clkbuf_4 _15881_ (.A(_14274_),
    .X(_14275_));
 sky130_fd_sc_hd__mux2_1 _15882_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][31] ),
    .A1(_13173_),
    .S(_14275_),
    .X(_14276_));
 sky130_fd_sc_hd__clkbuf_1 _15883_ (.A(_14276_),
    .X(_02083_));
 sky130_fd_sc_hd__mux2_1 _15884_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][30] ),
    .A1(_13184_),
    .S(_14275_),
    .X(_14277_));
 sky130_fd_sc_hd__clkbuf_1 _15885_ (.A(_14277_),
    .X(_02082_));
 sky130_fd_sc_hd__mux2_1 _15886_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][29] ),
    .A1(_13187_),
    .S(_14275_),
    .X(_14278_));
 sky130_fd_sc_hd__clkbuf_1 _15887_ (.A(_14278_),
    .X(_02081_));
 sky130_fd_sc_hd__mux2_1 _15888_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][28] ),
    .A1(_13190_),
    .S(_14275_),
    .X(_14279_));
 sky130_fd_sc_hd__clkbuf_1 _15889_ (.A(_14279_),
    .X(_02080_));
 sky130_fd_sc_hd__mux2_1 _15890_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][27] ),
    .A1(_13195_),
    .S(_14275_),
    .X(_14280_));
 sky130_fd_sc_hd__clkbuf_1 _15891_ (.A(_14280_),
    .X(_02079_));
 sky130_fd_sc_hd__mux2_1 _15892_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][26] ),
    .A1(_13198_),
    .S(_14275_),
    .X(_14281_));
 sky130_fd_sc_hd__clkbuf_1 _15893_ (.A(_14281_),
    .X(_02078_));
 sky130_fd_sc_hd__mux2_1 _15894_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][25] ),
    .A1(_13201_),
    .S(_14275_),
    .X(_14282_));
 sky130_fd_sc_hd__clkbuf_1 _15895_ (.A(_14282_),
    .X(_02077_));
 sky130_fd_sc_hd__mux2_1 _15896_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][24] ),
    .A1(_13204_),
    .S(_14275_),
    .X(_14283_));
 sky130_fd_sc_hd__clkbuf_1 _15897_ (.A(_14283_),
    .X(_02076_));
 sky130_fd_sc_hd__mux2_1 _15898_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][23] ),
    .A1(_13207_),
    .S(_14275_),
    .X(_14284_));
 sky130_fd_sc_hd__clkbuf_1 _15899_ (.A(_14284_),
    .X(_02075_));
 sky130_fd_sc_hd__mux2_1 _15900_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][22] ),
    .A1(_13210_),
    .S(_14275_),
    .X(_14285_));
 sky130_fd_sc_hd__clkbuf_1 _15901_ (.A(_14285_),
    .X(_02074_));
 sky130_fd_sc_hd__buf_4 _15902_ (.A(_14274_),
    .X(_14286_));
 sky130_fd_sc_hd__mux2_1 _15903_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][21] ),
    .A1(_13213_),
    .S(_14286_),
    .X(_14287_));
 sky130_fd_sc_hd__clkbuf_1 _15904_ (.A(_14287_),
    .X(_02073_));
 sky130_fd_sc_hd__mux2_1 _15905_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][20] ),
    .A1(_13217_),
    .S(_14286_),
    .X(_14288_));
 sky130_fd_sc_hd__clkbuf_1 _15906_ (.A(_14288_),
    .X(_02072_));
 sky130_fd_sc_hd__mux2_1 _15907_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][19] ),
    .A1(_13220_),
    .S(_14286_),
    .X(_14289_));
 sky130_fd_sc_hd__clkbuf_1 _15908_ (.A(_14289_),
    .X(_02071_));
 sky130_fd_sc_hd__mux2_1 _15909_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][18] ),
    .A1(_13223_),
    .S(_14286_),
    .X(_14290_));
 sky130_fd_sc_hd__clkbuf_1 _15910_ (.A(_14290_),
    .X(_02070_));
 sky130_fd_sc_hd__mux2_1 _15911_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][17] ),
    .A1(_13226_),
    .S(_14286_),
    .X(_14291_));
 sky130_fd_sc_hd__clkbuf_1 _15912_ (.A(_14291_),
    .X(_02069_));
 sky130_fd_sc_hd__mux2_1 _15913_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][16] ),
    .A1(_13229_),
    .S(_14286_),
    .X(_14292_));
 sky130_fd_sc_hd__clkbuf_1 _15914_ (.A(_14292_),
    .X(_02068_));
 sky130_fd_sc_hd__mux2_1 _15915_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][15] ),
    .A1(_13232_),
    .S(_14286_),
    .X(_14293_));
 sky130_fd_sc_hd__clkbuf_1 _15916_ (.A(_14293_),
    .X(_02067_));
 sky130_fd_sc_hd__mux2_1 _15917_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][14] ),
    .A1(_13235_),
    .S(_14286_),
    .X(_14294_));
 sky130_fd_sc_hd__clkbuf_1 _15918_ (.A(_14294_),
    .X(_02066_));
 sky130_fd_sc_hd__mux2_1 _15919_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][13] ),
    .A1(_13238_),
    .S(_14286_),
    .X(_14295_));
 sky130_fd_sc_hd__clkbuf_1 _15920_ (.A(_14295_),
    .X(_02065_));
 sky130_fd_sc_hd__mux2_1 _15921_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][12] ),
    .A1(_13241_),
    .S(_14286_),
    .X(_14296_));
 sky130_fd_sc_hd__clkbuf_1 _15922_ (.A(_14296_),
    .X(_02064_));
 sky130_fd_sc_hd__buf_4 _15923_ (.A(_14274_),
    .X(_14297_));
 sky130_fd_sc_hd__mux2_1 _15924_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][11] ),
    .A1(_13244_),
    .S(_14297_),
    .X(_14298_));
 sky130_fd_sc_hd__clkbuf_1 _15925_ (.A(_14298_),
    .X(_02063_));
 sky130_fd_sc_hd__mux2_1 _15926_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][10] ),
    .A1(_13248_),
    .S(_14297_),
    .X(_14299_));
 sky130_fd_sc_hd__clkbuf_1 _15927_ (.A(_14299_),
    .X(_02062_));
 sky130_fd_sc_hd__mux2_1 _15928_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][9] ),
    .A1(_13251_),
    .S(_14297_),
    .X(_14300_));
 sky130_fd_sc_hd__clkbuf_1 _15929_ (.A(_14300_),
    .X(_02061_));
 sky130_fd_sc_hd__mux2_1 _15930_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][8] ),
    .A1(_13254_),
    .S(_14297_),
    .X(_14301_));
 sky130_fd_sc_hd__clkbuf_1 _15931_ (.A(_14301_),
    .X(_02060_));
 sky130_fd_sc_hd__mux2_1 _15932_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][7] ),
    .A1(_13257_),
    .S(_14297_),
    .X(_14302_));
 sky130_fd_sc_hd__clkbuf_1 _15933_ (.A(_14302_),
    .X(_02059_));
 sky130_fd_sc_hd__mux2_1 _15934_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][6] ),
    .A1(_13260_),
    .S(_14297_),
    .X(_14303_));
 sky130_fd_sc_hd__clkbuf_1 _15935_ (.A(_14303_),
    .X(_02058_));
 sky130_fd_sc_hd__mux2_1 _15936_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][5] ),
    .A1(_13263_),
    .S(_14297_),
    .X(_14304_));
 sky130_fd_sc_hd__clkbuf_1 _15937_ (.A(_14304_),
    .X(_02057_));
 sky130_fd_sc_hd__mux2_1 _15938_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][4] ),
    .A1(_13266_),
    .S(_14297_),
    .X(_14305_));
 sky130_fd_sc_hd__clkbuf_1 _15939_ (.A(_14305_),
    .X(_02056_));
 sky130_fd_sc_hd__mux2_1 _15940_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][3] ),
    .A1(_13269_),
    .S(_14297_),
    .X(_14306_));
 sky130_fd_sc_hd__clkbuf_1 _15941_ (.A(_14306_),
    .X(_02055_));
 sky130_fd_sc_hd__mux2_1 _15942_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][2] ),
    .A1(_13272_),
    .S(_14297_),
    .X(_14307_));
 sky130_fd_sc_hd__clkbuf_1 _15943_ (.A(_14307_),
    .X(_02054_));
 sky130_fd_sc_hd__mux2_1 _15944_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][1] ),
    .A1(_13275_),
    .S(_14274_),
    .X(_14308_));
 sky130_fd_sc_hd__clkbuf_1 _15945_ (.A(_14308_),
    .X(_02053_));
 sky130_fd_sc_hd__mux2_1 _15946_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][0] ),
    .A1(_13278_),
    .S(_14274_),
    .X(_14309_));
 sky130_fd_sc_hd__clkbuf_1 _15947_ (.A(_14309_),
    .X(_02052_));
 sky130_fd_sc_hd__nor2_2 _15948_ (.A(_13179_),
    .B(_14271_),
    .Y(_14310_));
 sky130_fd_sc_hd__clkbuf_4 _15949_ (.A(_14310_),
    .X(_14311_));
 sky130_fd_sc_hd__mux2_1 _15950_ (.A0(\rvcpu.dp.rf.reg_file_arr[5][31] ),
    .A1(_13173_),
    .S(_14311_),
    .X(_14312_));
 sky130_fd_sc_hd__clkbuf_1 _15951_ (.A(_14312_),
    .X(_02051_));
 sky130_fd_sc_hd__mux2_1 _15952_ (.A0(\rvcpu.dp.rf.reg_file_arr[5][30] ),
    .A1(_13184_),
    .S(_14311_),
    .X(_14313_));
 sky130_fd_sc_hd__clkbuf_1 _15953_ (.A(_14313_),
    .X(_02050_));
 sky130_fd_sc_hd__mux2_1 _15954_ (.A0(\rvcpu.dp.rf.reg_file_arr[5][29] ),
    .A1(_13187_),
    .S(_14311_),
    .X(_14314_));
 sky130_fd_sc_hd__clkbuf_1 _15955_ (.A(_14314_),
    .X(_02049_));
 sky130_fd_sc_hd__mux2_1 _15956_ (.A0(\rvcpu.dp.rf.reg_file_arr[5][28] ),
    .A1(_13190_),
    .S(_14311_),
    .X(_14315_));
 sky130_fd_sc_hd__clkbuf_1 _15957_ (.A(_14315_),
    .X(_02048_));
 sky130_fd_sc_hd__mux2_1 _15958_ (.A0(\rvcpu.dp.rf.reg_file_arr[5][27] ),
    .A1(_13195_),
    .S(_14311_),
    .X(_14316_));
 sky130_fd_sc_hd__clkbuf_1 _15959_ (.A(_14316_),
    .X(_02047_));
 sky130_fd_sc_hd__mux2_1 _15960_ (.A0(\rvcpu.dp.rf.reg_file_arr[5][26] ),
    .A1(_13198_),
    .S(_14311_),
    .X(_14317_));
 sky130_fd_sc_hd__clkbuf_1 _15961_ (.A(_14317_),
    .X(_02046_));
 sky130_fd_sc_hd__mux2_1 _15962_ (.A0(\rvcpu.dp.rf.reg_file_arr[5][25] ),
    .A1(_13201_),
    .S(_14311_),
    .X(_14318_));
 sky130_fd_sc_hd__clkbuf_1 _15963_ (.A(_14318_),
    .X(_02045_));
 sky130_fd_sc_hd__mux2_1 _15964_ (.A0(\rvcpu.dp.rf.reg_file_arr[5][24] ),
    .A1(_13204_),
    .S(_14311_),
    .X(_14319_));
 sky130_fd_sc_hd__clkbuf_1 _15965_ (.A(_14319_),
    .X(_02044_));
 sky130_fd_sc_hd__mux2_1 _15966_ (.A0(\rvcpu.dp.rf.reg_file_arr[5][23] ),
    .A1(_13207_),
    .S(_14311_),
    .X(_14320_));
 sky130_fd_sc_hd__clkbuf_1 _15967_ (.A(_14320_),
    .X(_02043_));
 sky130_fd_sc_hd__mux2_1 _15968_ (.A0(\rvcpu.dp.rf.reg_file_arr[5][22] ),
    .A1(_13210_),
    .S(_14311_),
    .X(_14321_));
 sky130_fd_sc_hd__clkbuf_1 _15969_ (.A(_14321_),
    .X(_02042_));
 sky130_fd_sc_hd__buf_4 _15970_ (.A(_14310_),
    .X(_14322_));
 sky130_fd_sc_hd__mux2_1 _15971_ (.A0(\rvcpu.dp.rf.reg_file_arr[5][21] ),
    .A1(_13213_),
    .S(_14322_),
    .X(_14323_));
 sky130_fd_sc_hd__clkbuf_1 _15972_ (.A(_14323_),
    .X(_02041_));
 sky130_fd_sc_hd__mux2_1 _15973_ (.A0(\rvcpu.dp.rf.reg_file_arr[5][20] ),
    .A1(_13217_),
    .S(_14322_),
    .X(_14324_));
 sky130_fd_sc_hd__clkbuf_1 _15974_ (.A(_14324_),
    .X(_02040_));
 sky130_fd_sc_hd__mux2_1 _15975_ (.A0(\rvcpu.dp.rf.reg_file_arr[5][19] ),
    .A1(_13220_),
    .S(_14322_),
    .X(_14325_));
 sky130_fd_sc_hd__clkbuf_1 _15976_ (.A(_14325_),
    .X(_02039_));
 sky130_fd_sc_hd__mux2_1 _15977_ (.A0(\rvcpu.dp.rf.reg_file_arr[5][18] ),
    .A1(_13223_),
    .S(_14322_),
    .X(_14326_));
 sky130_fd_sc_hd__clkbuf_1 _15978_ (.A(_14326_),
    .X(_02038_));
 sky130_fd_sc_hd__mux2_1 _15979_ (.A0(\rvcpu.dp.rf.reg_file_arr[5][17] ),
    .A1(_13226_),
    .S(_14322_),
    .X(_14327_));
 sky130_fd_sc_hd__clkbuf_1 _15980_ (.A(_14327_),
    .X(_02037_));
 sky130_fd_sc_hd__mux2_1 _15981_ (.A0(\rvcpu.dp.rf.reg_file_arr[5][16] ),
    .A1(_13229_),
    .S(_14322_),
    .X(_14328_));
 sky130_fd_sc_hd__clkbuf_1 _15982_ (.A(_14328_),
    .X(_02036_));
 sky130_fd_sc_hd__mux2_1 _15983_ (.A0(\rvcpu.dp.rf.reg_file_arr[5][15] ),
    .A1(_13232_),
    .S(_14322_),
    .X(_14329_));
 sky130_fd_sc_hd__clkbuf_1 _15984_ (.A(_14329_),
    .X(_02035_));
 sky130_fd_sc_hd__mux2_1 _15985_ (.A0(\rvcpu.dp.rf.reg_file_arr[5][14] ),
    .A1(_13235_),
    .S(_14322_),
    .X(_14330_));
 sky130_fd_sc_hd__clkbuf_1 _15986_ (.A(_14330_),
    .X(_02034_));
 sky130_fd_sc_hd__mux2_1 _15987_ (.A0(\rvcpu.dp.rf.reg_file_arr[5][13] ),
    .A1(_13238_),
    .S(_14322_),
    .X(_14331_));
 sky130_fd_sc_hd__clkbuf_1 _15988_ (.A(_14331_),
    .X(_02033_));
 sky130_fd_sc_hd__mux2_1 _15989_ (.A0(\rvcpu.dp.rf.reg_file_arr[5][12] ),
    .A1(_13241_),
    .S(_14322_),
    .X(_14332_));
 sky130_fd_sc_hd__clkbuf_1 _15990_ (.A(_14332_),
    .X(_02032_));
 sky130_fd_sc_hd__clkbuf_4 _15991_ (.A(_14310_),
    .X(_14333_));
 sky130_fd_sc_hd__mux2_1 _15992_ (.A0(\rvcpu.dp.rf.reg_file_arr[5][11] ),
    .A1(_13244_),
    .S(_14333_),
    .X(_14334_));
 sky130_fd_sc_hd__clkbuf_1 _15993_ (.A(_14334_),
    .X(_02031_));
 sky130_fd_sc_hd__mux2_1 _15994_ (.A0(\rvcpu.dp.rf.reg_file_arr[5][10] ),
    .A1(_13248_),
    .S(_14333_),
    .X(_14335_));
 sky130_fd_sc_hd__clkbuf_1 _15995_ (.A(_14335_),
    .X(_02030_));
 sky130_fd_sc_hd__mux2_1 _15996_ (.A0(\rvcpu.dp.rf.reg_file_arr[5][9] ),
    .A1(_13251_),
    .S(_14333_),
    .X(_14336_));
 sky130_fd_sc_hd__clkbuf_1 _15997_ (.A(_14336_),
    .X(_02029_));
 sky130_fd_sc_hd__mux2_1 _15998_ (.A0(\rvcpu.dp.rf.reg_file_arr[5][8] ),
    .A1(_13254_),
    .S(_14333_),
    .X(_14337_));
 sky130_fd_sc_hd__clkbuf_1 _15999_ (.A(_14337_),
    .X(_02028_));
 sky130_fd_sc_hd__mux2_1 _16000_ (.A0(\rvcpu.dp.rf.reg_file_arr[5][7] ),
    .A1(_13257_),
    .S(_14333_),
    .X(_14338_));
 sky130_fd_sc_hd__clkbuf_1 _16001_ (.A(_14338_),
    .X(_02027_));
 sky130_fd_sc_hd__mux2_1 _16002_ (.A0(\rvcpu.dp.rf.reg_file_arr[5][6] ),
    .A1(_13260_),
    .S(_14333_),
    .X(_14339_));
 sky130_fd_sc_hd__clkbuf_1 _16003_ (.A(_14339_),
    .X(_02026_));
 sky130_fd_sc_hd__mux2_1 _16004_ (.A0(\rvcpu.dp.rf.reg_file_arr[5][5] ),
    .A1(_13263_),
    .S(_14333_),
    .X(_14340_));
 sky130_fd_sc_hd__clkbuf_1 _16005_ (.A(_14340_),
    .X(_02025_));
 sky130_fd_sc_hd__mux2_1 _16006_ (.A0(\rvcpu.dp.rf.reg_file_arr[5][4] ),
    .A1(_13266_),
    .S(_14333_),
    .X(_14341_));
 sky130_fd_sc_hd__clkbuf_1 _16007_ (.A(_14341_),
    .X(_02024_));
 sky130_fd_sc_hd__mux2_1 _16008_ (.A0(\rvcpu.dp.rf.reg_file_arr[5][3] ),
    .A1(_13269_),
    .S(_14333_),
    .X(_14342_));
 sky130_fd_sc_hd__clkbuf_1 _16009_ (.A(_14342_),
    .X(_02023_));
 sky130_fd_sc_hd__mux2_1 _16010_ (.A0(\rvcpu.dp.rf.reg_file_arr[5][2] ),
    .A1(_13272_),
    .S(_14333_),
    .X(_14343_));
 sky130_fd_sc_hd__clkbuf_1 _16011_ (.A(_14343_),
    .X(_02022_));
 sky130_fd_sc_hd__mux2_1 _16012_ (.A0(\rvcpu.dp.rf.reg_file_arr[5][1] ),
    .A1(_13275_),
    .S(_14310_),
    .X(_14344_));
 sky130_fd_sc_hd__clkbuf_1 _16013_ (.A(_14344_),
    .X(_02021_));
 sky130_fd_sc_hd__mux2_1 _16014_ (.A0(\rvcpu.dp.rf.reg_file_arr[5][0] ),
    .A1(_13278_),
    .S(_14310_),
    .X(_14345_));
 sky130_fd_sc_hd__clkbuf_1 _16015_ (.A(_14345_),
    .X(_02020_));
 sky130_fd_sc_hd__inv_2 _16016_ (.A(\rvcpu.dp.plmw.RdW[0] ),
    .Y(_14346_));
 sky130_fd_sc_hd__nand3_4 _16017_ (.A(\rvcpu.dp.plmw.RegWriteW ),
    .B(_14346_),
    .C(\rvcpu.dp.plmw.RdW[1] ),
    .Y(_14347_));
 sky130_fd_sc_hd__nor2_2 _16018_ (.A(_14271_),
    .B(_14347_),
    .Y(_14348_));
 sky130_fd_sc_hd__buf_4 _16019_ (.A(_14348_),
    .X(_14349_));
 sky130_fd_sc_hd__mux2_1 _16020_ (.A0(\rvcpu.dp.rf.reg_file_arr[6][31] ),
    .A1(_13173_),
    .S(_14349_),
    .X(_14350_));
 sky130_fd_sc_hd__clkbuf_1 _16021_ (.A(_14350_),
    .X(_02011_));
 sky130_fd_sc_hd__mux2_1 _16022_ (.A0(\rvcpu.dp.rf.reg_file_arr[6][30] ),
    .A1(_13184_),
    .S(_14349_),
    .X(_14351_));
 sky130_fd_sc_hd__clkbuf_1 _16023_ (.A(_14351_),
    .X(_02010_));
 sky130_fd_sc_hd__mux2_1 _16024_ (.A0(\rvcpu.dp.rf.reg_file_arr[6][29] ),
    .A1(_13187_),
    .S(_14349_),
    .X(_14352_));
 sky130_fd_sc_hd__clkbuf_1 _16025_ (.A(_14352_),
    .X(_02009_));
 sky130_fd_sc_hd__mux2_1 _16026_ (.A0(\rvcpu.dp.rf.reg_file_arr[6][28] ),
    .A1(_13190_),
    .S(_14349_),
    .X(_14353_));
 sky130_fd_sc_hd__clkbuf_1 _16027_ (.A(_14353_),
    .X(_02008_));
 sky130_fd_sc_hd__mux2_1 _16028_ (.A0(\rvcpu.dp.rf.reg_file_arr[6][27] ),
    .A1(_13195_),
    .S(_14349_),
    .X(_14354_));
 sky130_fd_sc_hd__clkbuf_1 _16029_ (.A(_14354_),
    .X(_02007_));
 sky130_fd_sc_hd__mux2_1 _16030_ (.A0(\rvcpu.dp.rf.reg_file_arr[6][26] ),
    .A1(_13198_),
    .S(_14349_),
    .X(_14355_));
 sky130_fd_sc_hd__clkbuf_1 _16031_ (.A(_14355_),
    .X(_02006_));
 sky130_fd_sc_hd__mux2_1 _16032_ (.A0(\rvcpu.dp.rf.reg_file_arr[6][25] ),
    .A1(_13201_),
    .S(_14349_),
    .X(_14356_));
 sky130_fd_sc_hd__clkbuf_1 _16033_ (.A(_14356_),
    .X(_02005_));
 sky130_fd_sc_hd__mux2_1 _16034_ (.A0(\rvcpu.dp.rf.reg_file_arr[6][24] ),
    .A1(_13204_),
    .S(_14349_),
    .X(_14357_));
 sky130_fd_sc_hd__clkbuf_1 _16035_ (.A(_14357_),
    .X(_02004_));
 sky130_fd_sc_hd__mux2_1 _16036_ (.A0(\rvcpu.dp.rf.reg_file_arr[6][23] ),
    .A1(_13207_),
    .S(_14349_),
    .X(_14358_));
 sky130_fd_sc_hd__clkbuf_1 _16037_ (.A(_14358_),
    .X(_02003_));
 sky130_fd_sc_hd__mux2_1 _16038_ (.A0(\rvcpu.dp.rf.reg_file_arr[6][22] ),
    .A1(_13210_),
    .S(_14349_),
    .X(_14359_));
 sky130_fd_sc_hd__clkbuf_1 _16039_ (.A(_14359_),
    .X(_02002_));
 sky130_fd_sc_hd__clkbuf_4 _16040_ (.A(_14348_),
    .X(_14360_));
 sky130_fd_sc_hd__mux2_1 _16041_ (.A0(\rvcpu.dp.rf.reg_file_arr[6][21] ),
    .A1(_13213_),
    .S(_14360_),
    .X(_14361_));
 sky130_fd_sc_hd__clkbuf_1 _16042_ (.A(_14361_),
    .X(_02001_));
 sky130_fd_sc_hd__mux2_1 _16043_ (.A0(\rvcpu.dp.rf.reg_file_arr[6][20] ),
    .A1(_13217_),
    .S(_14360_),
    .X(_14362_));
 sky130_fd_sc_hd__clkbuf_1 _16044_ (.A(_14362_),
    .X(_02000_));
 sky130_fd_sc_hd__mux2_1 _16045_ (.A0(\rvcpu.dp.rf.reg_file_arr[6][19] ),
    .A1(_13220_),
    .S(_14360_),
    .X(_14363_));
 sky130_fd_sc_hd__clkbuf_1 _16046_ (.A(_14363_),
    .X(_01999_));
 sky130_fd_sc_hd__mux2_1 _16047_ (.A0(\rvcpu.dp.rf.reg_file_arr[6][18] ),
    .A1(_13223_),
    .S(_14360_),
    .X(_14364_));
 sky130_fd_sc_hd__clkbuf_1 _16048_ (.A(_14364_),
    .X(_01998_));
 sky130_fd_sc_hd__mux2_1 _16049_ (.A0(\rvcpu.dp.rf.reg_file_arr[6][17] ),
    .A1(_13226_),
    .S(_14360_),
    .X(_14365_));
 sky130_fd_sc_hd__clkbuf_1 _16050_ (.A(_14365_),
    .X(_01997_));
 sky130_fd_sc_hd__mux2_1 _16051_ (.A0(\rvcpu.dp.rf.reg_file_arr[6][16] ),
    .A1(_13229_),
    .S(_14360_),
    .X(_14366_));
 sky130_fd_sc_hd__clkbuf_1 _16052_ (.A(_14366_),
    .X(_01996_));
 sky130_fd_sc_hd__mux2_1 _16053_ (.A0(\rvcpu.dp.rf.reg_file_arr[6][15] ),
    .A1(_13232_),
    .S(_14360_),
    .X(_14367_));
 sky130_fd_sc_hd__clkbuf_1 _16054_ (.A(_14367_),
    .X(_01995_));
 sky130_fd_sc_hd__mux2_1 _16055_ (.A0(\rvcpu.dp.rf.reg_file_arr[6][14] ),
    .A1(_13235_),
    .S(_14360_),
    .X(_14368_));
 sky130_fd_sc_hd__clkbuf_1 _16056_ (.A(_14368_),
    .X(_01994_));
 sky130_fd_sc_hd__mux2_1 _16057_ (.A0(\rvcpu.dp.rf.reg_file_arr[6][13] ),
    .A1(_13238_),
    .S(_14360_),
    .X(_14369_));
 sky130_fd_sc_hd__clkbuf_1 _16058_ (.A(_14369_),
    .X(_01993_));
 sky130_fd_sc_hd__mux2_1 _16059_ (.A0(\rvcpu.dp.rf.reg_file_arr[6][12] ),
    .A1(_13241_),
    .S(_14360_),
    .X(_14370_));
 sky130_fd_sc_hd__clkbuf_1 _16060_ (.A(_14370_),
    .X(_01992_));
 sky130_fd_sc_hd__clkbuf_4 _16061_ (.A(_14348_),
    .X(_14371_));
 sky130_fd_sc_hd__mux2_1 _16062_ (.A0(\rvcpu.dp.rf.reg_file_arr[6][11] ),
    .A1(_13244_),
    .S(_14371_),
    .X(_14372_));
 sky130_fd_sc_hd__clkbuf_1 _16063_ (.A(_14372_),
    .X(_01991_));
 sky130_fd_sc_hd__mux2_1 _16064_ (.A0(\rvcpu.dp.rf.reg_file_arr[6][10] ),
    .A1(_13248_),
    .S(_14371_),
    .X(_14373_));
 sky130_fd_sc_hd__clkbuf_1 _16065_ (.A(_14373_),
    .X(_01990_));
 sky130_fd_sc_hd__mux2_1 _16066_ (.A0(\rvcpu.dp.rf.reg_file_arr[6][9] ),
    .A1(_13251_),
    .S(_14371_),
    .X(_14374_));
 sky130_fd_sc_hd__clkbuf_1 _16067_ (.A(_14374_),
    .X(_01989_));
 sky130_fd_sc_hd__mux2_1 _16068_ (.A0(\rvcpu.dp.rf.reg_file_arr[6][8] ),
    .A1(_13254_),
    .S(_14371_),
    .X(_14375_));
 sky130_fd_sc_hd__clkbuf_1 _16069_ (.A(_14375_),
    .X(_01988_));
 sky130_fd_sc_hd__mux2_1 _16070_ (.A0(\rvcpu.dp.rf.reg_file_arr[6][7] ),
    .A1(_13257_),
    .S(_14371_),
    .X(_14376_));
 sky130_fd_sc_hd__clkbuf_1 _16071_ (.A(_14376_),
    .X(_01987_));
 sky130_fd_sc_hd__mux2_1 _16072_ (.A0(\rvcpu.dp.rf.reg_file_arr[6][6] ),
    .A1(_13260_),
    .S(_14371_),
    .X(_14377_));
 sky130_fd_sc_hd__clkbuf_1 _16073_ (.A(_14377_),
    .X(_01986_));
 sky130_fd_sc_hd__mux2_1 _16074_ (.A0(\rvcpu.dp.rf.reg_file_arr[6][5] ),
    .A1(_13263_),
    .S(_14371_),
    .X(_14378_));
 sky130_fd_sc_hd__clkbuf_1 _16075_ (.A(_14378_),
    .X(_01985_));
 sky130_fd_sc_hd__mux2_1 _16076_ (.A0(\rvcpu.dp.rf.reg_file_arr[6][4] ),
    .A1(_13266_),
    .S(_14371_),
    .X(_14379_));
 sky130_fd_sc_hd__clkbuf_1 _16077_ (.A(_14379_),
    .X(_01984_));
 sky130_fd_sc_hd__mux2_1 _16078_ (.A0(\rvcpu.dp.rf.reg_file_arr[6][3] ),
    .A1(_13269_),
    .S(_14371_),
    .X(_14380_));
 sky130_fd_sc_hd__clkbuf_1 _16079_ (.A(_14380_),
    .X(_01983_));
 sky130_fd_sc_hd__mux2_1 _16080_ (.A0(\rvcpu.dp.rf.reg_file_arr[6][2] ),
    .A1(_13272_),
    .S(_14371_),
    .X(_14381_));
 sky130_fd_sc_hd__clkbuf_1 _16081_ (.A(_14381_),
    .X(_01982_));
 sky130_fd_sc_hd__mux2_1 _16082_ (.A0(\rvcpu.dp.rf.reg_file_arr[6][1] ),
    .A1(_13275_),
    .S(_14348_),
    .X(_14382_));
 sky130_fd_sc_hd__clkbuf_1 _16083_ (.A(_14382_),
    .X(_01981_));
 sky130_fd_sc_hd__mux2_1 _16084_ (.A0(\rvcpu.dp.rf.reg_file_arr[6][0] ),
    .A1(_13278_),
    .S(_14348_),
    .X(_14383_));
 sky130_fd_sc_hd__clkbuf_1 _16085_ (.A(_14383_),
    .X(_01980_));
 sky130_fd_sc_hd__nor2_2 _16086_ (.A(_14090_),
    .B(_14271_),
    .Y(_14384_));
 sky130_fd_sc_hd__buf_4 _16087_ (.A(_14384_),
    .X(_14385_));
 sky130_fd_sc_hd__mux2_1 _16088_ (.A0(\rvcpu.dp.rf.reg_file_arr[7][31] ),
    .A1(_13173_),
    .S(_14385_),
    .X(_14386_));
 sky130_fd_sc_hd__clkbuf_1 _16089_ (.A(_14386_),
    .X(_01979_));
 sky130_fd_sc_hd__mux2_1 _16090_ (.A0(\rvcpu.dp.rf.reg_file_arr[7][30] ),
    .A1(_13184_),
    .S(_14385_),
    .X(_14387_));
 sky130_fd_sc_hd__clkbuf_1 _16091_ (.A(_14387_),
    .X(_01978_));
 sky130_fd_sc_hd__mux2_1 _16092_ (.A0(\rvcpu.dp.rf.reg_file_arr[7][29] ),
    .A1(_13187_),
    .S(_14385_),
    .X(_14388_));
 sky130_fd_sc_hd__clkbuf_1 _16093_ (.A(_14388_),
    .X(_01977_));
 sky130_fd_sc_hd__mux2_1 _16094_ (.A0(\rvcpu.dp.rf.reg_file_arr[7][28] ),
    .A1(_13190_),
    .S(_14385_),
    .X(_14389_));
 sky130_fd_sc_hd__clkbuf_1 _16095_ (.A(_14389_),
    .X(_01976_));
 sky130_fd_sc_hd__mux2_1 _16096_ (.A0(\rvcpu.dp.rf.reg_file_arr[7][27] ),
    .A1(_13195_),
    .S(_14385_),
    .X(_14390_));
 sky130_fd_sc_hd__clkbuf_1 _16097_ (.A(_14390_),
    .X(_01975_));
 sky130_fd_sc_hd__mux2_1 _16098_ (.A0(\rvcpu.dp.rf.reg_file_arr[7][26] ),
    .A1(_13198_),
    .S(_14385_),
    .X(_14391_));
 sky130_fd_sc_hd__clkbuf_1 _16099_ (.A(_14391_),
    .X(_01974_));
 sky130_fd_sc_hd__mux2_1 _16100_ (.A0(\rvcpu.dp.rf.reg_file_arr[7][25] ),
    .A1(_13201_),
    .S(_14385_),
    .X(_14392_));
 sky130_fd_sc_hd__clkbuf_1 _16101_ (.A(_14392_),
    .X(_01973_));
 sky130_fd_sc_hd__mux2_1 _16102_ (.A0(\rvcpu.dp.rf.reg_file_arr[7][24] ),
    .A1(_13204_),
    .S(_14385_),
    .X(_14393_));
 sky130_fd_sc_hd__clkbuf_1 _16103_ (.A(_14393_),
    .X(_01972_));
 sky130_fd_sc_hd__mux2_1 _16104_ (.A0(\rvcpu.dp.rf.reg_file_arr[7][23] ),
    .A1(_13207_),
    .S(_14385_),
    .X(_14394_));
 sky130_fd_sc_hd__clkbuf_1 _16105_ (.A(_14394_),
    .X(_01971_));
 sky130_fd_sc_hd__mux2_1 _16106_ (.A0(\rvcpu.dp.rf.reg_file_arr[7][22] ),
    .A1(_13210_),
    .S(_14385_),
    .X(_14395_));
 sky130_fd_sc_hd__clkbuf_1 _16107_ (.A(_14395_),
    .X(_01970_));
 sky130_fd_sc_hd__buf_4 _16108_ (.A(_14384_),
    .X(_14396_));
 sky130_fd_sc_hd__mux2_1 _16109_ (.A0(\rvcpu.dp.rf.reg_file_arr[7][21] ),
    .A1(_13213_),
    .S(_14396_),
    .X(_14397_));
 sky130_fd_sc_hd__clkbuf_1 _16110_ (.A(_14397_),
    .X(_01969_));
 sky130_fd_sc_hd__mux2_1 _16111_ (.A0(\rvcpu.dp.rf.reg_file_arr[7][20] ),
    .A1(_13217_),
    .S(_14396_),
    .X(_14398_));
 sky130_fd_sc_hd__clkbuf_1 _16112_ (.A(_14398_),
    .X(_01968_));
 sky130_fd_sc_hd__mux2_1 _16113_ (.A0(\rvcpu.dp.rf.reg_file_arr[7][19] ),
    .A1(_13220_),
    .S(_14396_),
    .X(_14399_));
 sky130_fd_sc_hd__clkbuf_1 _16114_ (.A(_14399_),
    .X(_01967_));
 sky130_fd_sc_hd__mux2_1 _16115_ (.A0(\rvcpu.dp.rf.reg_file_arr[7][18] ),
    .A1(_13223_),
    .S(_14396_),
    .X(_14400_));
 sky130_fd_sc_hd__clkbuf_1 _16116_ (.A(_14400_),
    .X(_01966_));
 sky130_fd_sc_hd__mux2_1 _16117_ (.A0(\rvcpu.dp.rf.reg_file_arr[7][17] ),
    .A1(_13226_),
    .S(_14396_),
    .X(_14401_));
 sky130_fd_sc_hd__clkbuf_1 _16118_ (.A(_14401_),
    .X(_01965_));
 sky130_fd_sc_hd__mux2_1 _16119_ (.A0(\rvcpu.dp.rf.reg_file_arr[7][16] ),
    .A1(_13229_),
    .S(_14396_),
    .X(_14402_));
 sky130_fd_sc_hd__clkbuf_1 _16120_ (.A(_14402_),
    .X(_01964_));
 sky130_fd_sc_hd__mux2_1 _16121_ (.A0(\rvcpu.dp.rf.reg_file_arr[7][15] ),
    .A1(_13232_),
    .S(_14396_),
    .X(_14403_));
 sky130_fd_sc_hd__clkbuf_1 _16122_ (.A(_14403_),
    .X(_01963_));
 sky130_fd_sc_hd__mux2_1 _16123_ (.A0(\rvcpu.dp.rf.reg_file_arr[7][14] ),
    .A1(_13235_),
    .S(_14396_),
    .X(_14404_));
 sky130_fd_sc_hd__clkbuf_1 _16124_ (.A(_14404_),
    .X(_01962_));
 sky130_fd_sc_hd__mux2_1 _16125_ (.A0(\rvcpu.dp.rf.reg_file_arr[7][13] ),
    .A1(_13238_),
    .S(_14396_),
    .X(_14405_));
 sky130_fd_sc_hd__clkbuf_1 _16126_ (.A(_14405_),
    .X(_01961_));
 sky130_fd_sc_hd__mux2_1 _16127_ (.A0(\rvcpu.dp.rf.reg_file_arr[7][12] ),
    .A1(_13241_),
    .S(_14396_),
    .X(_14406_));
 sky130_fd_sc_hd__clkbuf_1 _16128_ (.A(_14406_),
    .X(_01960_));
 sky130_fd_sc_hd__clkbuf_4 _16129_ (.A(_14384_),
    .X(_14407_));
 sky130_fd_sc_hd__mux2_1 _16130_ (.A0(\rvcpu.dp.rf.reg_file_arr[7][11] ),
    .A1(_13244_),
    .S(_14407_),
    .X(_14408_));
 sky130_fd_sc_hd__clkbuf_1 _16131_ (.A(_14408_),
    .X(_01959_));
 sky130_fd_sc_hd__mux2_1 _16132_ (.A0(\rvcpu.dp.rf.reg_file_arr[7][10] ),
    .A1(_13248_),
    .S(_14407_),
    .X(_14409_));
 sky130_fd_sc_hd__clkbuf_1 _16133_ (.A(_14409_),
    .X(_01958_));
 sky130_fd_sc_hd__mux2_1 _16134_ (.A0(\rvcpu.dp.rf.reg_file_arr[7][9] ),
    .A1(_13251_),
    .S(_14407_),
    .X(_14410_));
 sky130_fd_sc_hd__clkbuf_1 _16135_ (.A(_14410_),
    .X(_01957_));
 sky130_fd_sc_hd__mux2_1 _16136_ (.A0(\rvcpu.dp.rf.reg_file_arr[7][8] ),
    .A1(_13254_),
    .S(_14407_),
    .X(_14411_));
 sky130_fd_sc_hd__clkbuf_1 _16137_ (.A(_14411_),
    .X(_01956_));
 sky130_fd_sc_hd__mux2_1 _16138_ (.A0(\rvcpu.dp.rf.reg_file_arr[7][7] ),
    .A1(_13257_),
    .S(_14407_),
    .X(_14412_));
 sky130_fd_sc_hd__clkbuf_1 _16139_ (.A(_14412_),
    .X(_01955_));
 sky130_fd_sc_hd__mux2_1 _16140_ (.A0(\rvcpu.dp.rf.reg_file_arr[7][6] ),
    .A1(_13260_),
    .S(_14407_),
    .X(_14413_));
 sky130_fd_sc_hd__clkbuf_1 _16141_ (.A(_14413_),
    .X(_01954_));
 sky130_fd_sc_hd__mux2_1 _16142_ (.A0(\rvcpu.dp.rf.reg_file_arr[7][5] ),
    .A1(_13263_),
    .S(_14407_),
    .X(_14414_));
 sky130_fd_sc_hd__clkbuf_1 _16143_ (.A(_14414_),
    .X(_01953_));
 sky130_fd_sc_hd__mux2_1 _16144_ (.A0(\rvcpu.dp.rf.reg_file_arr[7][4] ),
    .A1(_13266_),
    .S(_14407_),
    .X(_14415_));
 sky130_fd_sc_hd__clkbuf_1 _16145_ (.A(_14415_),
    .X(_01952_));
 sky130_fd_sc_hd__mux2_1 _16146_ (.A0(\rvcpu.dp.rf.reg_file_arr[7][3] ),
    .A1(_13269_),
    .S(_14407_),
    .X(_14416_));
 sky130_fd_sc_hd__clkbuf_1 _16147_ (.A(_14416_),
    .X(_01951_));
 sky130_fd_sc_hd__mux2_1 _16148_ (.A0(\rvcpu.dp.rf.reg_file_arr[7][2] ),
    .A1(_13272_),
    .S(_14407_),
    .X(_14417_));
 sky130_fd_sc_hd__clkbuf_1 _16149_ (.A(_14417_),
    .X(_01950_));
 sky130_fd_sc_hd__mux2_1 _16150_ (.A0(\rvcpu.dp.rf.reg_file_arr[7][1] ),
    .A1(_13275_),
    .S(_14384_),
    .X(_14418_));
 sky130_fd_sc_hd__clkbuf_1 _16151_ (.A(_14418_),
    .X(_01949_));
 sky130_fd_sc_hd__mux2_1 _16152_ (.A0(\rvcpu.dp.rf.reg_file_arr[7][0] ),
    .A1(_13278_),
    .S(_14384_),
    .X(_14419_));
 sky130_fd_sc_hd__clkbuf_1 _16153_ (.A(_14419_),
    .X(_01948_));
 sky130_fd_sc_hd__clkbuf_4 _16154_ (.A(_13172_),
    .X(_14420_));
 sky130_fd_sc_hd__nor2_2 _16155_ (.A(_13177_),
    .B(_14273_),
    .Y(_14421_));
 sky130_fd_sc_hd__buf_4 _16156_ (.A(_14421_),
    .X(_14422_));
 sky130_fd_sc_hd__mux2_1 _16157_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][31] ),
    .A1(_14420_),
    .S(_14422_),
    .X(_14423_));
 sky130_fd_sc_hd__clkbuf_1 _16158_ (.A(_14423_),
    .X(_01947_));
 sky130_fd_sc_hd__clkbuf_4 _16159_ (.A(_13183_),
    .X(_14424_));
 sky130_fd_sc_hd__mux2_1 _16160_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][30] ),
    .A1(_14424_),
    .S(_14422_),
    .X(_14425_));
 sky130_fd_sc_hd__clkbuf_1 _16161_ (.A(_14425_),
    .X(_01946_));
 sky130_fd_sc_hd__clkbuf_4 _16162_ (.A(_13186_),
    .X(_14426_));
 sky130_fd_sc_hd__mux2_1 _16163_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][29] ),
    .A1(_14426_),
    .S(_14422_),
    .X(_14427_));
 sky130_fd_sc_hd__clkbuf_1 _16164_ (.A(_14427_),
    .X(_01945_));
 sky130_fd_sc_hd__clkbuf_4 _16165_ (.A(_13189_),
    .X(_14428_));
 sky130_fd_sc_hd__mux2_1 _16166_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][28] ),
    .A1(_14428_),
    .S(_14422_),
    .X(_14429_));
 sky130_fd_sc_hd__clkbuf_1 _16167_ (.A(_14429_),
    .X(_01944_));
 sky130_fd_sc_hd__clkbuf_4 _16168_ (.A(_13194_),
    .X(_14430_));
 sky130_fd_sc_hd__mux2_1 _16169_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][27] ),
    .A1(_14430_),
    .S(_14422_),
    .X(_14431_));
 sky130_fd_sc_hd__clkbuf_1 _16170_ (.A(_14431_),
    .X(_01943_));
 sky130_fd_sc_hd__buf_4 _16171_ (.A(_13197_),
    .X(_14432_));
 sky130_fd_sc_hd__mux2_1 _16172_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][26] ),
    .A1(_14432_),
    .S(_14422_),
    .X(_14433_));
 sky130_fd_sc_hd__clkbuf_1 _16173_ (.A(_14433_),
    .X(_01942_));
 sky130_fd_sc_hd__buf_4 _16174_ (.A(_13200_),
    .X(_14434_));
 sky130_fd_sc_hd__mux2_1 _16175_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][25] ),
    .A1(_14434_),
    .S(_14422_),
    .X(_14435_));
 sky130_fd_sc_hd__clkbuf_1 _16176_ (.A(_14435_),
    .X(_01941_));
 sky130_fd_sc_hd__clkbuf_4 _16177_ (.A(_13203_),
    .X(_14436_));
 sky130_fd_sc_hd__mux2_1 _16178_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][24] ),
    .A1(_14436_),
    .S(_14422_),
    .X(_14437_));
 sky130_fd_sc_hd__clkbuf_1 _16179_ (.A(_14437_),
    .X(_01940_));
 sky130_fd_sc_hd__buf_4 _16180_ (.A(_13206_),
    .X(_14438_));
 sky130_fd_sc_hd__mux2_1 _16181_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][23] ),
    .A1(_14438_),
    .S(_14422_),
    .X(_14439_));
 sky130_fd_sc_hd__clkbuf_1 _16182_ (.A(_14439_),
    .X(_01939_));
 sky130_fd_sc_hd__clkbuf_4 _16183_ (.A(_13209_),
    .X(_14440_));
 sky130_fd_sc_hd__mux2_1 _16184_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][22] ),
    .A1(_14440_),
    .S(_14422_),
    .X(_14441_));
 sky130_fd_sc_hd__clkbuf_1 _16185_ (.A(_14441_),
    .X(_01938_));
 sky130_fd_sc_hd__buf_4 _16186_ (.A(_13212_),
    .X(_14442_));
 sky130_fd_sc_hd__clkbuf_4 _16187_ (.A(_14421_),
    .X(_14443_));
 sky130_fd_sc_hd__mux2_1 _16188_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][21] ),
    .A1(_14442_),
    .S(_14443_),
    .X(_14444_));
 sky130_fd_sc_hd__clkbuf_1 _16189_ (.A(_14444_),
    .X(_01937_));
 sky130_fd_sc_hd__buf_4 _16190_ (.A(_13216_),
    .X(_14445_));
 sky130_fd_sc_hd__mux2_1 _16191_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][20] ),
    .A1(_14445_),
    .S(_14443_),
    .X(_14446_));
 sky130_fd_sc_hd__clkbuf_1 _16192_ (.A(_14446_),
    .X(_01936_));
 sky130_fd_sc_hd__buf_4 _16193_ (.A(_13219_),
    .X(_14447_));
 sky130_fd_sc_hd__mux2_1 _16194_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][19] ),
    .A1(_14447_),
    .S(_14443_),
    .X(_14448_));
 sky130_fd_sc_hd__clkbuf_1 _16195_ (.A(_14448_),
    .X(_01935_));
 sky130_fd_sc_hd__buf_4 _16196_ (.A(_13222_),
    .X(_14449_));
 sky130_fd_sc_hd__mux2_1 _16197_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][18] ),
    .A1(_14449_),
    .S(_14443_),
    .X(_14450_));
 sky130_fd_sc_hd__clkbuf_1 _16198_ (.A(_14450_),
    .X(_01934_));
 sky130_fd_sc_hd__buf_4 _16199_ (.A(_13225_),
    .X(_14451_));
 sky130_fd_sc_hd__mux2_1 _16200_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][17] ),
    .A1(_14451_),
    .S(_14443_),
    .X(_14452_));
 sky130_fd_sc_hd__clkbuf_1 _16201_ (.A(_14452_),
    .X(_01933_));
 sky130_fd_sc_hd__buf_4 _16202_ (.A(_13228_),
    .X(_14453_));
 sky130_fd_sc_hd__mux2_1 _16203_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][16] ),
    .A1(_14453_),
    .S(_14443_),
    .X(_14454_));
 sky130_fd_sc_hd__clkbuf_1 _16204_ (.A(_14454_),
    .X(_01932_));
 sky130_fd_sc_hd__buf_4 _16205_ (.A(_13231_),
    .X(_14455_));
 sky130_fd_sc_hd__mux2_1 _16206_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][15] ),
    .A1(_14455_),
    .S(_14443_),
    .X(_14456_));
 sky130_fd_sc_hd__clkbuf_1 _16207_ (.A(_14456_),
    .X(_01931_));
 sky130_fd_sc_hd__buf_4 _16208_ (.A(_13234_),
    .X(_14457_));
 sky130_fd_sc_hd__mux2_1 _16209_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][14] ),
    .A1(_14457_),
    .S(_14443_),
    .X(_14458_));
 sky130_fd_sc_hd__clkbuf_1 _16210_ (.A(_14458_),
    .X(_01930_));
 sky130_fd_sc_hd__buf_4 _16211_ (.A(_13237_),
    .X(_14459_));
 sky130_fd_sc_hd__mux2_1 _16212_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][13] ),
    .A1(_14459_),
    .S(_14443_),
    .X(_14460_));
 sky130_fd_sc_hd__clkbuf_1 _16213_ (.A(_14460_),
    .X(_01929_));
 sky130_fd_sc_hd__buf_4 _16214_ (.A(_13240_),
    .X(_14461_));
 sky130_fd_sc_hd__mux2_1 _16215_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][12] ),
    .A1(_14461_),
    .S(_14443_),
    .X(_14462_));
 sky130_fd_sc_hd__clkbuf_1 _16216_ (.A(_14462_),
    .X(_01928_));
 sky130_fd_sc_hd__buf_4 _16217_ (.A(_13243_),
    .X(_14463_));
 sky130_fd_sc_hd__buf_4 _16218_ (.A(_14421_),
    .X(_14464_));
 sky130_fd_sc_hd__mux2_1 _16219_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][11] ),
    .A1(_14463_),
    .S(_14464_),
    .X(_14465_));
 sky130_fd_sc_hd__clkbuf_1 _16220_ (.A(_14465_),
    .X(_01927_));
 sky130_fd_sc_hd__buf_4 _16221_ (.A(_13247_),
    .X(_14466_));
 sky130_fd_sc_hd__mux2_1 _16222_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][10] ),
    .A1(_14466_),
    .S(_14464_),
    .X(_14467_));
 sky130_fd_sc_hd__clkbuf_1 _16223_ (.A(_14467_),
    .X(_01926_));
 sky130_fd_sc_hd__buf_4 _16224_ (.A(_13250_),
    .X(_14468_));
 sky130_fd_sc_hd__mux2_1 _16225_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][9] ),
    .A1(_14468_),
    .S(_14464_),
    .X(_14469_));
 sky130_fd_sc_hd__clkbuf_1 _16226_ (.A(_14469_),
    .X(_01925_));
 sky130_fd_sc_hd__buf_4 _16227_ (.A(_13253_),
    .X(_14470_));
 sky130_fd_sc_hd__mux2_1 _16228_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][8] ),
    .A1(_14470_),
    .S(_14464_),
    .X(_14471_));
 sky130_fd_sc_hd__clkbuf_1 _16229_ (.A(_14471_),
    .X(_01924_));
 sky130_fd_sc_hd__buf_4 _16230_ (.A(_13256_),
    .X(_14472_));
 sky130_fd_sc_hd__mux2_1 _16231_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][7] ),
    .A1(_14472_),
    .S(_14464_),
    .X(_14473_));
 sky130_fd_sc_hd__clkbuf_1 _16232_ (.A(_14473_),
    .X(_01923_));
 sky130_fd_sc_hd__buf_4 _16233_ (.A(_13259_),
    .X(_14474_));
 sky130_fd_sc_hd__mux2_1 _16234_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][6] ),
    .A1(_14474_),
    .S(_14464_),
    .X(_14475_));
 sky130_fd_sc_hd__clkbuf_1 _16235_ (.A(_14475_),
    .X(_01922_));
 sky130_fd_sc_hd__buf_4 _16236_ (.A(_13262_),
    .X(_14476_));
 sky130_fd_sc_hd__mux2_1 _16237_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][5] ),
    .A1(_14476_),
    .S(_14464_),
    .X(_14477_));
 sky130_fd_sc_hd__clkbuf_1 _16238_ (.A(_14477_),
    .X(_01921_));
 sky130_fd_sc_hd__buf_4 _16239_ (.A(_13265_),
    .X(_14478_));
 sky130_fd_sc_hd__mux2_1 _16240_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][4] ),
    .A1(_14478_),
    .S(_14464_),
    .X(_14479_));
 sky130_fd_sc_hd__clkbuf_1 _16241_ (.A(_14479_),
    .X(_01920_));
 sky130_fd_sc_hd__buf_4 _16242_ (.A(_13268_),
    .X(_14480_));
 sky130_fd_sc_hd__mux2_1 _16243_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][3] ),
    .A1(_14480_),
    .S(_14464_),
    .X(_14481_));
 sky130_fd_sc_hd__clkbuf_1 _16244_ (.A(_14481_),
    .X(_01919_));
 sky130_fd_sc_hd__buf_4 _16245_ (.A(_13271_),
    .X(_14482_));
 sky130_fd_sc_hd__mux2_1 _16246_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][2] ),
    .A1(_14482_),
    .S(_14464_),
    .X(_14483_));
 sky130_fd_sc_hd__clkbuf_1 _16247_ (.A(_14483_),
    .X(_01918_));
 sky130_fd_sc_hd__clkbuf_4 _16248_ (.A(_13274_),
    .X(_14484_));
 sky130_fd_sc_hd__mux2_1 _16249_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][1] ),
    .A1(_14484_),
    .S(_14421_),
    .X(_14485_));
 sky130_fd_sc_hd__clkbuf_1 _16250_ (.A(_14485_),
    .X(_01917_));
 sky130_fd_sc_hd__buf_4 _16251_ (.A(_13277_),
    .X(_14486_));
 sky130_fd_sc_hd__mux2_1 _16252_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][0] ),
    .A1(_14486_),
    .S(_14421_),
    .X(_14487_));
 sky130_fd_sc_hd__clkbuf_1 _16253_ (.A(_14487_),
    .X(_01916_));
 sky130_fd_sc_hd__nor2_2 _16254_ (.A(_14234_),
    .B(_14273_),
    .Y(_14488_));
 sky130_fd_sc_hd__clkbuf_4 _16255_ (.A(_14488_),
    .X(_14489_));
 sky130_fd_sc_hd__mux2_1 _16256_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][31] ),
    .A1(_14420_),
    .S(_14489_),
    .X(_14490_));
 sky130_fd_sc_hd__clkbuf_1 _16257_ (.A(_14490_),
    .X(_01907_));
 sky130_fd_sc_hd__mux2_1 _16258_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][30] ),
    .A1(_14424_),
    .S(_14489_),
    .X(_14491_));
 sky130_fd_sc_hd__clkbuf_1 _16259_ (.A(_14491_),
    .X(_01906_));
 sky130_fd_sc_hd__mux2_1 _16260_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][29] ),
    .A1(_14426_),
    .S(_14489_),
    .X(_14492_));
 sky130_fd_sc_hd__clkbuf_1 _16261_ (.A(_14492_),
    .X(_01905_));
 sky130_fd_sc_hd__mux2_1 _16262_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][28] ),
    .A1(_14428_),
    .S(_14489_),
    .X(_14493_));
 sky130_fd_sc_hd__clkbuf_1 _16263_ (.A(_14493_),
    .X(_01904_));
 sky130_fd_sc_hd__mux2_1 _16264_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][27] ),
    .A1(_14430_),
    .S(_14489_),
    .X(_14494_));
 sky130_fd_sc_hd__clkbuf_1 _16265_ (.A(_14494_),
    .X(_01903_));
 sky130_fd_sc_hd__mux2_1 _16266_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][26] ),
    .A1(_14432_),
    .S(_14489_),
    .X(_14495_));
 sky130_fd_sc_hd__clkbuf_1 _16267_ (.A(_14495_),
    .X(_01902_));
 sky130_fd_sc_hd__mux2_1 _16268_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][25] ),
    .A1(_14434_),
    .S(_14489_),
    .X(_14496_));
 sky130_fd_sc_hd__clkbuf_1 _16269_ (.A(_14496_),
    .X(_01901_));
 sky130_fd_sc_hd__mux2_1 _16270_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][24] ),
    .A1(_14436_),
    .S(_14489_),
    .X(_14497_));
 sky130_fd_sc_hd__clkbuf_1 _16271_ (.A(_14497_),
    .X(_01900_));
 sky130_fd_sc_hd__mux2_1 _16272_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][23] ),
    .A1(_14438_),
    .S(_14489_),
    .X(_14498_));
 sky130_fd_sc_hd__clkbuf_1 _16273_ (.A(_14498_),
    .X(_01899_));
 sky130_fd_sc_hd__mux2_1 _16274_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][22] ),
    .A1(_14440_),
    .S(_14489_),
    .X(_14499_));
 sky130_fd_sc_hd__clkbuf_1 _16275_ (.A(_14499_),
    .X(_01898_));
 sky130_fd_sc_hd__buf_4 _16276_ (.A(_14488_),
    .X(_14500_));
 sky130_fd_sc_hd__mux2_1 _16277_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][21] ),
    .A1(_14442_),
    .S(_14500_),
    .X(_14501_));
 sky130_fd_sc_hd__clkbuf_1 _16278_ (.A(_14501_),
    .X(_01897_));
 sky130_fd_sc_hd__mux2_1 _16279_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][20] ),
    .A1(_14445_),
    .S(_14500_),
    .X(_14502_));
 sky130_fd_sc_hd__clkbuf_1 _16280_ (.A(_14502_),
    .X(_01896_));
 sky130_fd_sc_hd__mux2_1 _16281_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][19] ),
    .A1(_14447_),
    .S(_14500_),
    .X(_14503_));
 sky130_fd_sc_hd__clkbuf_1 _16282_ (.A(_14503_),
    .X(_01895_));
 sky130_fd_sc_hd__mux2_1 _16283_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][18] ),
    .A1(_14449_),
    .S(_14500_),
    .X(_14504_));
 sky130_fd_sc_hd__clkbuf_1 _16284_ (.A(_14504_),
    .X(_01894_));
 sky130_fd_sc_hd__mux2_1 _16285_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][17] ),
    .A1(_14451_),
    .S(_14500_),
    .X(_14505_));
 sky130_fd_sc_hd__clkbuf_1 _16286_ (.A(_14505_),
    .X(_01893_));
 sky130_fd_sc_hd__mux2_1 _16287_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][16] ),
    .A1(_14453_),
    .S(_14500_),
    .X(_14506_));
 sky130_fd_sc_hd__clkbuf_1 _16288_ (.A(_14506_),
    .X(_01892_));
 sky130_fd_sc_hd__mux2_1 _16289_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][15] ),
    .A1(_14455_),
    .S(_14500_),
    .X(_14507_));
 sky130_fd_sc_hd__clkbuf_1 _16290_ (.A(_14507_),
    .X(_01891_));
 sky130_fd_sc_hd__mux2_1 _16291_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][14] ),
    .A1(_14457_),
    .S(_14500_),
    .X(_14508_));
 sky130_fd_sc_hd__clkbuf_1 _16292_ (.A(_14508_),
    .X(_01890_));
 sky130_fd_sc_hd__mux2_1 _16293_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][13] ),
    .A1(_14459_),
    .S(_14500_),
    .X(_14509_));
 sky130_fd_sc_hd__clkbuf_1 _16294_ (.A(_14509_),
    .X(_01889_));
 sky130_fd_sc_hd__mux2_1 _16295_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][12] ),
    .A1(_14461_),
    .S(_14500_),
    .X(_14510_));
 sky130_fd_sc_hd__clkbuf_1 _16296_ (.A(_14510_),
    .X(_01888_));
 sky130_fd_sc_hd__clkbuf_4 _16297_ (.A(_14488_),
    .X(_14511_));
 sky130_fd_sc_hd__mux2_1 _16298_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][11] ),
    .A1(_14463_),
    .S(_14511_),
    .X(_14512_));
 sky130_fd_sc_hd__clkbuf_1 _16299_ (.A(_14512_),
    .X(_01887_));
 sky130_fd_sc_hd__mux2_1 _16300_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][10] ),
    .A1(_14466_),
    .S(_14511_),
    .X(_14513_));
 sky130_fd_sc_hd__clkbuf_1 _16301_ (.A(_14513_),
    .X(_01886_));
 sky130_fd_sc_hd__mux2_1 _16302_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][9] ),
    .A1(_14468_),
    .S(_14511_),
    .X(_14514_));
 sky130_fd_sc_hd__clkbuf_1 _16303_ (.A(_14514_),
    .X(_01885_));
 sky130_fd_sc_hd__mux2_1 _16304_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][8] ),
    .A1(_14470_),
    .S(_14511_),
    .X(_14515_));
 sky130_fd_sc_hd__clkbuf_1 _16305_ (.A(_14515_),
    .X(_01884_));
 sky130_fd_sc_hd__mux2_1 _16306_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][7] ),
    .A1(_14472_),
    .S(_14511_),
    .X(_14516_));
 sky130_fd_sc_hd__clkbuf_1 _16307_ (.A(_14516_),
    .X(_01883_));
 sky130_fd_sc_hd__mux2_1 _16308_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][6] ),
    .A1(_14474_),
    .S(_14511_),
    .X(_14517_));
 sky130_fd_sc_hd__clkbuf_1 _16309_ (.A(_14517_),
    .X(_01882_));
 sky130_fd_sc_hd__mux2_1 _16310_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][5] ),
    .A1(_14476_),
    .S(_14511_),
    .X(_14518_));
 sky130_fd_sc_hd__clkbuf_1 _16311_ (.A(_14518_),
    .X(_01881_));
 sky130_fd_sc_hd__mux2_1 _16312_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][4] ),
    .A1(_14478_),
    .S(_14511_),
    .X(_14519_));
 sky130_fd_sc_hd__clkbuf_1 _16313_ (.A(_14519_),
    .X(_01880_));
 sky130_fd_sc_hd__mux2_1 _16314_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][3] ),
    .A1(_14480_),
    .S(_14511_),
    .X(_14520_));
 sky130_fd_sc_hd__clkbuf_1 _16315_ (.A(_14520_),
    .X(_01879_));
 sky130_fd_sc_hd__mux2_1 _16316_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][2] ),
    .A1(_14482_),
    .S(_14511_),
    .X(_14521_));
 sky130_fd_sc_hd__clkbuf_1 _16317_ (.A(_14521_),
    .X(_01878_));
 sky130_fd_sc_hd__mux2_1 _16318_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][1] ),
    .A1(_14484_),
    .S(_14488_),
    .X(_14522_));
 sky130_fd_sc_hd__clkbuf_1 _16319_ (.A(_14522_),
    .X(_01877_));
 sky130_fd_sc_hd__mux2_1 _16320_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][0] ),
    .A1(_14486_),
    .S(_14488_),
    .X(_14523_));
 sky130_fd_sc_hd__clkbuf_1 _16321_ (.A(_14523_),
    .X(_01876_));
 sky130_fd_sc_hd__nor2_2 _16322_ (.A(_13177_),
    .B(_14347_),
    .Y(_14524_));
 sky130_fd_sc_hd__buf_4 _16323_ (.A(_14524_),
    .X(_14525_));
 sky130_fd_sc_hd__mux2_1 _16324_ (.A0(\rvcpu.dp.rf.reg_file_arr[10][31] ),
    .A1(_14420_),
    .S(_14525_),
    .X(_14526_));
 sky130_fd_sc_hd__clkbuf_1 _16325_ (.A(_14526_),
    .X(_01875_));
 sky130_fd_sc_hd__mux2_1 _16326_ (.A0(\rvcpu.dp.rf.reg_file_arr[10][30] ),
    .A1(_14424_),
    .S(_14525_),
    .X(_14527_));
 sky130_fd_sc_hd__clkbuf_1 _16327_ (.A(_14527_),
    .X(_01874_));
 sky130_fd_sc_hd__mux2_1 _16328_ (.A0(\rvcpu.dp.rf.reg_file_arr[10][29] ),
    .A1(_14426_),
    .S(_14525_),
    .X(_14528_));
 sky130_fd_sc_hd__clkbuf_1 _16329_ (.A(_14528_),
    .X(_01873_));
 sky130_fd_sc_hd__mux2_1 _16330_ (.A0(\rvcpu.dp.rf.reg_file_arr[10][28] ),
    .A1(_14428_),
    .S(_14525_),
    .X(_14529_));
 sky130_fd_sc_hd__clkbuf_1 _16331_ (.A(_14529_),
    .X(_01872_));
 sky130_fd_sc_hd__mux2_1 _16332_ (.A0(\rvcpu.dp.rf.reg_file_arr[10][27] ),
    .A1(_14430_),
    .S(_14525_),
    .X(_14530_));
 sky130_fd_sc_hd__clkbuf_1 _16333_ (.A(_14530_),
    .X(_01871_));
 sky130_fd_sc_hd__mux2_1 _16334_ (.A0(\rvcpu.dp.rf.reg_file_arr[10][26] ),
    .A1(_14432_),
    .S(_14525_),
    .X(_14531_));
 sky130_fd_sc_hd__clkbuf_1 _16335_ (.A(_14531_),
    .X(_01870_));
 sky130_fd_sc_hd__mux2_1 _16336_ (.A0(\rvcpu.dp.rf.reg_file_arr[10][25] ),
    .A1(_14434_),
    .S(_14525_),
    .X(_14532_));
 sky130_fd_sc_hd__clkbuf_1 _16337_ (.A(_14532_),
    .X(_01869_));
 sky130_fd_sc_hd__mux2_1 _16338_ (.A0(\rvcpu.dp.rf.reg_file_arr[10][24] ),
    .A1(_14436_),
    .S(_14525_),
    .X(_14533_));
 sky130_fd_sc_hd__clkbuf_1 _16339_ (.A(_14533_),
    .X(_01868_));
 sky130_fd_sc_hd__mux2_1 _16340_ (.A0(\rvcpu.dp.rf.reg_file_arr[10][23] ),
    .A1(_14438_),
    .S(_14525_),
    .X(_14534_));
 sky130_fd_sc_hd__clkbuf_1 _16341_ (.A(_14534_),
    .X(_01867_));
 sky130_fd_sc_hd__mux2_1 _16342_ (.A0(\rvcpu.dp.rf.reg_file_arr[10][22] ),
    .A1(_14440_),
    .S(_14525_),
    .X(_14535_));
 sky130_fd_sc_hd__clkbuf_1 _16343_ (.A(_14535_),
    .X(_01866_));
 sky130_fd_sc_hd__clkbuf_4 _16344_ (.A(_14524_),
    .X(_14536_));
 sky130_fd_sc_hd__mux2_1 _16345_ (.A0(\rvcpu.dp.rf.reg_file_arr[10][21] ),
    .A1(_14442_),
    .S(_14536_),
    .X(_14537_));
 sky130_fd_sc_hd__clkbuf_1 _16346_ (.A(_14537_),
    .X(_01865_));
 sky130_fd_sc_hd__mux2_1 _16347_ (.A0(\rvcpu.dp.rf.reg_file_arr[10][20] ),
    .A1(_14445_),
    .S(_14536_),
    .X(_14538_));
 sky130_fd_sc_hd__clkbuf_1 _16348_ (.A(_14538_),
    .X(_01864_));
 sky130_fd_sc_hd__mux2_1 _16349_ (.A0(\rvcpu.dp.rf.reg_file_arr[10][19] ),
    .A1(_14447_),
    .S(_14536_),
    .X(_14539_));
 sky130_fd_sc_hd__clkbuf_1 _16350_ (.A(_14539_),
    .X(_01863_));
 sky130_fd_sc_hd__mux2_1 _16351_ (.A0(\rvcpu.dp.rf.reg_file_arr[10][18] ),
    .A1(_14449_),
    .S(_14536_),
    .X(_14540_));
 sky130_fd_sc_hd__clkbuf_1 _16352_ (.A(_14540_),
    .X(_01862_));
 sky130_fd_sc_hd__mux2_1 _16353_ (.A0(\rvcpu.dp.rf.reg_file_arr[10][17] ),
    .A1(_14451_),
    .S(_14536_),
    .X(_14541_));
 sky130_fd_sc_hd__clkbuf_1 _16354_ (.A(_14541_),
    .X(_01861_));
 sky130_fd_sc_hd__mux2_1 _16355_ (.A0(\rvcpu.dp.rf.reg_file_arr[10][16] ),
    .A1(_14453_),
    .S(_14536_),
    .X(_14542_));
 sky130_fd_sc_hd__clkbuf_1 _16356_ (.A(_14542_),
    .X(_01860_));
 sky130_fd_sc_hd__mux2_1 _16357_ (.A0(\rvcpu.dp.rf.reg_file_arr[10][15] ),
    .A1(_14455_),
    .S(_14536_),
    .X(_14543_));
 sky130_fd_sc_hd__clkbuf_1 _16358_ (.A(_14543_),
    .X(_01859_));
 sky130_fd_sc_hd__mux2_1 _16359_ (.A0(\rvcpu.dp.rf.reg_file_arr[10][14] ),
    .A1(_14457_),
    .S(_14536_),
    .X(_14544_));
 sky130_fd_sc_hd__clkbuf_1 _16360_ (.A(_14544_),
    .X(_01858_));
 sky130_fd_sc_hd__mux2_1 _16361_ (.A0(\rvcpu.dp.rf.reg_file_arr[10][13] ),
    .A1(_14459_),
    .S(_14536_),
    .X(_14545_));
 sky130_fd_sc_hd__clkbuf_1 _16362_ (.A(_14545_),
    .X(_01857_));
 sky130_fd_sc_hd__mux2_1 _16363_ (.A0(\rvcpu.dp.rf.reg_file_arr[10][12] ),
    .A1(_14461_),
    .S(_14536_),
    .X(_14546_));
 sky130_fd_sc_hd__clkbuf_1 _16364_ (.A(_14546_),
    .X(_01856_));
 sky130_fd_sc_hd__clkbuf_4 _16365_ (.A(_14524_),
    .X(_14547_));
 sky130_fd_sc_hd__mux2_1 _16366_ (.A0(\rvcpu.dp.rf.reg_file_arr[10][11] ),
    .A1(_14463_),
    .S(_14547_),
    .X(_14548_));
 sky130_fd_sc_hd__clkbuf_1 _16367_ (.A(_14548_),
    .X(_01855_));
 sky130_fd_sc_hd__mux2_1 _16368_ (.A0(\rvcpu.dp.rf.reg_file_arr[10][10] ),
    .A1(_14466_),
    .S(_14547_),
    .X(_14549_));
 sky130_fd_sc_hd__clkbuf_1 _16369_ (.A(_14549_),
    .X(_01854_));
 sky130_fd_sc_hd__mux2_1 _16370_ (.A0(\rvcpu.dp.rf.reg_file_arr[10][9] ),
    .A1(_14468_),
    .S(_14547_),
    .X(_14550_));
 sky130_fd_sc_hd__clkbuf_1 _16371_ (.A(_14550_),
    .X(_01853_));
 sky130_fd_sc_hd__mux2_1 _16372_ (.A0(\rvcpu.dp.rf.reg_file_arr[10][8] ),
    .A1(_14470_),
    .S(_14547_),
    .X(_14551_));
 sky130_fd_sc_hd__clkbuf_1 _16373_ (.A(_14551_),
    .X(_01852_));
 sky130_fd_sc_hd__mux2_1 _16374_ (.A0(\rvcpu.dp.rf.reg_file_arr[10][7] ),
    .A1(_14472_),
    .S(_14547_),
    .X(_14552_));
 sky130_fd_sc_hd__clkbuf_1 _16375_ (.A(_14552_),
    .X(_01851_));
 sky130_fd_sc_hd__mux2_1 _16376_ (.A0(\rvcpu.dp.rf.reg_file_arr[10][6] ),
    .A1(_14474_),
    .S(_14547_),
    .X(_14553_));
 sky130_fd_sc_hd__clkbuf_1 _16377_ (.A(_14553_),
    .X(_01850_));
 sky130_fd_sc_hd__mux2_1 _16378_ (.A0(\rvcpu.dp.rf.reg_file_arr[10][5] ),
    .A1(_14476_),
    .S(_14547_),
    .X(_14554_));
 sky130_fd_sc_hd__clkbuf_1 _16379_ (.A(_14554_),
    .X(_01849_));
 sky130_fd_sc_hd__mux2_1 _16380_ (.A0(\rvcpu.dp.rf.reg_file_arr[10][4] ),
    .A1(_14478_),
    .S(_14547_),
    .X(_14555_));
 sky130_fd_sc_hd__clkbuf_1 _16381_ (.A(_14555_),
    .X(_01848_));
 sky130_fd_sc_hd__mux2_1 _16382_ (.A0(\rvcpu.dp.rf.reg_file_arr[10][3] ),
    .A1(_14480_),
    .S(_14547_),
    .X(_14556_));
 sky130_fd_sc_hd__clkbuf_1 _16383_ (.A(_14556_),
    .X(_01847_));
 sky130_fd_sc_hd__mux2_1 _16384_ (.A0(\rvcpu.dp.rf.reg_file_arr[10][2] ),
    .A1(_14482_),
    .S(_14547_),
    .X(_14557_));
 sky130_fd_sc_hd__clkbuf_1 _16385_ (.A(_14557_),
    .X(_01846_));
 sky130_fd_sc_hd__mux2_1 _16386_ (.A0(\rvcpu.dp.rf.reg_file_arr[10][1] ),
    .A1(_14484_),
    .S(_14524_),
    .X(_14558_));
 sky130_fd_sc_hd__clkbuf_1 _16387_ (.A(_14558_),
    .X(_01845_));
 sky130_fd_sc_hd__mux2_1 _16388_ (.A0(\rvcpu.dp.rf.reg_file_arr[10][0] ),
    .A1(_14486_),
    .S(_14524_),
    .X(_14559_));
 sky130_fd_sc_hd__clkbuf_1 _16389_ (.A(_14559_),
    .X(_01844_));
 sky130_fd_sc_hd__nor2_2 _16390_ (.A(_13177_),
    .B(_14090_),
    .Y(_14560_));
 sky130_fd_sc_hd__buf_4 _16391_ (.A(_14560_),
    .X(_14561_));
 sky130_fd_sc_hd__mux2_1 _16392_ (.A0(\rvcpu.dp.rf.reg_file_arr[11][31] ),
    .A1(_14420_),
    .S(_14561_),
    .X(_14562_));
 sky130_fd_sc_hd__clkbuf_1 _16393_ (.A(_14562_),
    .X(_01843_));
 sky130_fd_sc_hd__mux2_1 _16394_ (.A0(\rvcpu.dp.rf.reg_file_arr[11][30] ),
    .A1(_14424_),
    .S(_14561_),
    .X(_14563_));
 sky130_fd_sc_hd__clkbuf_1 _16395_ (.A(_14563_),
    .X(_01842_));
 sky130_fd_sc_hd__mux2_1 _16396_ (.A0(\rvcpu.dp.rf.reg_file_arr[11][29] ),
    .A1(_14426_),
    .S(_14561_),
    .X(_14564_));
 sky130_fd_sc_hd__clkbuf_1 _16397_ (.A(_14564_),
    .X(_01841_));
 sky130_fd_sc_hd__mux2_1 _16398_ (.A0(\rvcpu.dp.rf.reg_file_arr[11][28] ),
    .A1(_14428_),
    .S(_14561_),
    .X(_14565_));
 sky130_fd_sc_hd__clkbuf_1 _16399_ (.A(_14565_),
    .X(_01840_));
 sky130_fd_sc_hd__mux2_1 _16400_ (.A0(\rvcpu.dp.rf.reg_file_arr[11][27] ),
    .A1(_14430_),
    .S(_14561_),
    .X(_14566_));
 sky130_fd_sc_hd__clkbuf_1 _16401_ (.A(_14566_),
    .X(_01839_));
 sky130_fd_sc_hd__mux2_1 _16402_ (.A0(\rvcpu.dp.rf.reg_file_arr[11][26] ),
    .A1(_14432_),
    .S(_14561_),
    .X(_14567_));
 sky130_fd_sc_hd__clkbuf_1 _16403_ (.A(_14567_),
    .X(_01838_));
 sky130_fd_sc_hd__mux2_1 _16404_ (.A0(\rvcpu.dp.rf.reg_file_arr[11][25] ),
    .A1(_14434_),
    .S(_14561_),
    .X(_14568_));
 sky130_fd_sc_hd__clkbuf_1 _16405_ (.A(_14568_),
    .X(_01837_));
 sky130_fd_sc_hd__mux2_1 _16406_ (.A0(\rvcpu.dp.rf.reg_file_arr[11][24] ),
    .A1(_14436_),
    .S(_14561_),
    .X(_14569_));
 sky130_fd_sc_hd__clkbuf_1 _16407_ (.A(_14569_),
    .X(_01836_));
 sky130_fd_sc_hd__mux2_1 _16408_ (.A0(\rvcpu.dp.rf.reg_file_arr[11][23] ),
    .A1(_14438_),
    .S(_14561_),
    .X(_14570_));
 sky130_fd_sc_hd__clkbuf_1 _16409_ (.A(_14570_),
    .X(_01835_));
 sky130_fd_sc_hd__mux2_1 _16410_ (.A0(\rvcpu.dp.rf.reg_file_arr[11][22] ),
    .A1(_14440_),
    .S(_14561_),
    .X(_14571_));
 sky130_fd_sc_hd__clkbuf_1 _16411_ (.A(_14571_),
    .X(_01834_));
 sky130_fd_sc_hd__clkbuf_4 _16412_ (.A(_14560_),
    .X(_14572_));
 sky130_fd_sc_hd__mux2_1 _16413_ (.A0(\rvcpu.dp.rf.reg_file_arr[11][21] ),
    .A1(_14442_),
    .S(_14572_),
    .X(_14573_));
 sky130_fd_sc_hd__clkbuf_1 _16414_ (.A(_14573_),
    .X(_01833_));
 sky130_fd_sc_hd__mux2_1 _16415_ (.A0(\rvcpu.dp.rf.reg_file_arr[11][20] ),
    .A1(_14445_),
    .S(_14572_),
    .X(_14574_));
 sky130_fd_sc_hd__clkbuf_1 _16416_ (.A(_14574_),
    .X(_01832_));
 sky130_fd_sc_hd__mux2_1 _16417_ (.A0(\rvcpu.dp.rf.reg_file_arr[11][19] ),
    .A1(_14447_),
    .S(_14572_),
    .X(_14575_));
 sky130_fd_sc_hd__clkbuf_1 _16418_ (.A(_14575_),
    .X(_01831_));
 sky130_fd_sc_hd__mux2_1 _16419_ (.A0(\rvcpu.dp.rf.reg_file_arr[11][18] ),
    .A1(_14449_),
    .S(_14572_),
    .X(_14576_));
 sky130_fd_sc_hd__clkbuf_1 _16420_ (.A(_14576_),
    .X(_01830_));
 sky130_fd_sc_hd__mux2_1 _16421_ (.A0(\rvcpu.dp.rf.reg_file_arr[11][17] ),
    .A1(_14451_),
    .S(_14572_),
    .X(_14577_));
 sky130_fd_sc_hd__clkbuf_1 _16422_ (.A(_14577_),
    .X(_01829_));
 sky130_fd_sc_hd__mux2_1 _16423_ (.A0(\rvcpu.dp.rf.reg_file_arr[11][16] ),
    .A1(_14453_),
    .S(_14572_),
    .X(_14578_));
 sky130_fd_sc_hd__clkbuf_1 _16424_ (.A(_14578_),
    .X(_01828_));
 sky130_fd_sc_hd__mux2_1 _16425_ (.A0(\rvcpu.dp.rf.reg_file_arr[11][15] ),
    .A1(_14455_),
    .S(_14572_),
    .X(_14579_));
 sky130_fd_sc_hd__clkbuf_1 _16426_ (.A(_14579_),
    .X(_01827_));
 sky130_fd_sc_hd__mux2_1 _16427_ (.A0(\rvcpu.dp.rf.reg_file_arr[11][14] ),
    .A1(_14457_),
    .S(_14572_),
    .X(_14580_));
 sky130_fd_sc_hd__clkbuf_1 _16428_ (.A(_14580_),
    .X(_01826_));
 sky130_fd_sc_hd__mux2_1 _16429_ (.A0(\rvcpu.dp.rf.reg_file_arr[11][13] ),
    .A1(_14459_),
    .S(_14572_),
    .X(_14581_));
 sky130_fd_sc_hd__clkbuf_1 _16430_ (.A(_14581_),
    .X(_01825_));
 sky130_fd_sc_hd__mux2_1 _16431_ (.A0(\rvcpu.dp.rf.reg_file_arr[11][12] ),
    .A1(_14461_),
    .S(_14572_),
    .X(_14582_));
 sky130_fd_sc_hd__clkbuf_1 _16432_ (.A(_14582_),
    .X(_01824_));
 sky130_fd_sc_hd__clkbuf_4 _16433_ (.A(_14560_),
    .X(_04451_));
 sky130_fd_sc_hd__mux2_1 _16434_ (.A0(\rvcpu.dp.rf.reg_file_arr[11][11] ),
    .A1(_14463_),
    .S(_04451_),
    .X(_04452_));
 sky130_fd_sc_hd__clkbuf_1 _16435_ (.A(_04452_),
    .X(_01823_));
 sky130_fd_sc_hd__mux2_1 _16436_ (.A0(\rvcpu.dp.rf.reg_file_arr[11][10] ),
    .A1(_14466_),
    .S(_04451_),
    .X(_04453_));
 sky130_fd_sc_hd__clkbuf_1 _16437_ (.A(_04453_),
    .X(_01822_));
 sky130_fd_sc_hd__mux2_1 _16438_ (.A0(\rvcpu.dp.rf.reg_file_arr[11][9] ),
    .A1(_14468_),
    .S(_04451_),
    .X(_04454_));
 sky130_fd_sc_hd__clkbuf_1 _16439_ (.A(_04454_),
    .X(_01821_));
 sky130_fd_sc_hd__mux2_1 _16440_ (.A0(\rvcpu.dp.rf.reg_file_arr[11][8] ),
    .A1(_14470_),
    .S(_04451_),
    .X(_04455_));
 sky130_fd_sc_hd__clkbuf_1 _16441_ (.A(_04455_),
    .X(_01820_));
 sky130_fd_sc_hd__mux2_1 _16442_ (.A0(\rvcpu.dp.rf.reg_file_arr[11][7] ),
    .A1(_14472_),
    .S(_04451_),
    .X(_04456_));
 sky130_fd_sc_hd__clkbuf_1 _16443_ (.A(_04456_),
    .X(_01819_));
 sky130_fd_sc_hd__mux2_1 _16444_ (.A0(\rvcpu.dp.rf.reg_file_arr[11][6] ),
    .A1(_14474_),
    .S(_04451_),
    .X(_04457_));
 sky130_fd_sc_hd__clkbuf_1 _16445_ (.A(_04457_),
    .X(_01818_));
 sky130_fd_sc_hd__mux2_1 _16446_ (.A0(\rvcpu.dp.rf.reg_file_arr[11][5] ),
    .A1(_14476_),
    .S(_04451_),
    .X(_04458_));
 sky130_fd_sc_hd__clkbuf_1 _16447_ (.A(_04458_),
    .X(_01817_));
 sky130_fd_sc_hd__mux2_1 _16448_ (.A0(\rvcpu.dp.rf.reg_file_arr[11][4] ),
    .A1(_14478_),
    .S(_04451_),
    .X(_04459_));
 sky130_fd_sc_hd__clkbuf_1 _16449_ (.A(_04459_),
    .X(_01816_));
 sky130_fd_sc_hd__mux2_1 _16450_ (.A0(\rvcpu.dp.rf.reg_file_arr[11][3] ),
    .A1(_14480_),
    .S(_04451_),
    .X(_04460_));
 sky130_fd_sc_hd__clkbuf_1 _16451_ (.A(_04460_),
    .X(_01815_));
 sky130_fd_sc_hd__mux2_1 _16452_ (.A0(\rvcpu.dp.rf.reg_file_arr[11][2] ),
    .A1(_14482_),
    .S(_04451_),
    .X(_04461_));
 sky130_fd_sc_hd__clkbuf_1 _16453_ (.A(_04461_),
    .X(_01814_));
 sky130_fd_sc_hd__mux2_1 _16454_ (.A0(\rvcpu.dp.rf.reg_file_arr[11][1] ),
    .A1(_14484_),
    .S(_14560_),
    .X(_04462_));
 sky130_fd_sc_hd__clkbuf_1 _16455_ (.A(_04462_),
    .X(_01813_));
 sky130_fd_sc_hd__mux2_1 _16456_ (.A0(\rvcpu.dp.rf.reg_file_arr[11][0] ),
    .A1(_14486_),
    .S(_14560_),
    .X(_04463_));
 sky130_fd_sc_hd__clkbuf_1 _16457_ (.A(_04463_),
    .X(_01812_));
 sky130_fd_sc_hd__inv_2 _16458_ (.A(_14273_),
    .Y(_04464_));
 sky130_fd_sc_hd__and3b_2 _16459_ (.A_N(_13176_),
    .B(\rvcpu.dp.plmw.RdW[3] ),
    .C(_13174_),
    .X(_04465_));
 sky130_fd_sc_hd__and2_2 _16460_ (.A(_04464_),
    .B(_04465_),
    .X(_04466_));
 sky130_fd_sc_hd__clkbuf_4 _16461_ (.A(_04466_),
    .X(_04467_));
 sky130_fd_sc_hd__mux2_1 _16462_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][31] ),
    .A1(_14420_),
    .S(_04467_),
    .X(_04468_));
 sky130_fd_sc_hd__clkbuf_1 _16463_ (.A(_04468_),
    .X(_01811_));
 sky130_fd_sc_hd__mux2_1 _16464_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][30] ),
    .A1(_14424_),
    .S(_04467_),
    .X(_04469_));
 sky130_fd_sc_hd__clkbuf_1 _16465_ (.A(_04469_),
    .X(_01810_));
 sky130_fd_sc_hd__mux2_1 _16466_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][29] ),
    .A1(_14426_),
    .S(_04467_),
    .X(_04470_));
 sky130_fd_sc_hd__clkbuf_1 _16467_ (.A(_04470_),
    .X(_01809_));
 sky130_fd_sc_hd__mux2_1 _16468_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][28] ),
    .A1(_14428_),
    .S(_04467_),
    .X(_04471_));
 sky130_fd_sc_hd__clkbuf_1 _16469_ (.A(_04471_),
    .X(_01808_));
 sky130_fd_sc_hd__mux2_1 _16470_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][27] ),
    .A1(_14430_),
    .S(_04467_),
    .X(_04472_));
 sky130_fd_sc_hd__clkbuf_1 _16471_ (.A(_04472_),
    .X(_01807_));
 sky130_fd_sc_hd__mux2_1 _16472_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][26] ),
    .A1(_14432_),
    .S(_04467_),
    .X(_04473_));
 sky130_fd_sc_hd__clkbuf_1 _16473_ (.A(_04473_),
    .X(_01806_));
 sky130_fd_sc_hd__mux2_1 _16474_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][25] ),
    .A1(_14434_),
    .S(_04467_),
    .X(_04474_));
 sky130_fd_sc_hd__clkbuf_1 _16475_ (.A(_04474_),
    .X(_01805_));
 sky130_fd_sc_hd__mux2_1 _16476_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][24] ),
    .A1(_14436_),
    .S(_04467_),
    .X(_04475_));
 sky130_fd_sc_hd__clkbuf_1 _16477_ (.A(_04475_),
    .X(_01804_));
 sky130_fd_sc_hd__mux2_1 _16478_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][23] ),
    .A1(_14438_),
    .S(_04467_),
    .X(_04476_));
 sky130_fd_sc_hd__clkbuf_1 _16479_ (.A(_04476_),
    .X(_01803_));
 sky130_fd_sc_hd__mux2_1 _16480_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][22] ),
    .A1(_14440_),
    .S(_04467_),
    .X(_04477_));
 sky130_fd_sc_hd__clkbuf_1 _16481_ (.A(_04477_),
    .X(_01802_));
 sky130_fd_sc_hd__clkbuf_4 _16482_ (.A(_04466_),
    .X(_04478_));
 sky130_fd_sc_hd__mux2_1 _16483_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][21] ),
    .A1(_14442_),
    .S(_04478_),
    .X(_04479_));
 sky130_fd_sc_hd__clkbuf_1 _16484_ (.A(_04479_),
    .X(_01801_));
 sky130_fd_sc_hd__mux2_1 _16485_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][20] ),
    .A1(_14445_),
    .S(_04478_),
    .X(_04480_));
 sky130_fd_sc_hd__clkbuf_1 _16486_ (.A(_04480_),
    .X(_01800_));
 sky130_fd_sc_hd__mux2_1 _16487_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][19] ),
    .A1(_14447_),
    .S(_04478_),
    .X(_04481_));
 sky130_fd_sc_hd__clkbuf_1 _16488_ (.A(_04481_),
    .X(_01799_));
 sky130_fd_sc_hd__mux2_1 _16489_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][18] ),
    .A1(_14449_),
    .S(_04478_),
    .X(_04482_));
 sky130_fd_sc_hd__clkbuf_1 _16490_ (.A(_04482_),
    .X(_01798_));
 sky130_fd_sc_hd__mux2_1 _16491_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][17] ),
    .A1(_14451_),
    .S(_04478_),
    .X(_04483_));
 sky130_fd_sc_hd__clkbuf_1 _16492_ (.A(_04483_),
    .X(_01797_));
 sky130_fd_sc_hd__mux2_1 _16493_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][16] ),
    .A1(_14453_),
    .S(_04478_),
    .X(_04484_));
 sky130_fd_sc_hd__clkbuf_1 _16494_ (.A(_04484_),
    .X(_01796_));
 sky130_fd_sc_hd__mux2_1 _16495_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][15] ),
    .A1(_14455_),
    .S(_04478_),
    .X(_04485_));
 sky130_fd_sc_hd__clkbuf_1 _16496_ (.A(_04485_),
    .X(_01795_));
 sky130_fd_sc_hd__mux2_1 _16497_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][14] ),
    .A1(_14457_),
    .S(_04478_),
    .X(_04486_));
 sky130_fd_sc_hd__clkbuf_1 _16498_ (.A(_04486_),
    .X(_01794_));
 sky130_fd_sc_hd__mux2_1 _16499_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][13] ),
    .A1(_14459_),
    .S(_04478_),
    .X(_04487_));
 sky130_fd_sc_hd__clkbuf_1 _16500_ (.A(_04487_),
    .X(_01793_));
 sky130_fd_sc_hd__mux2_1 _16501_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][12] ),
    .A1(_14461_),
    .S(_04478_),
    .X(_04488_));
 sky130_fd_sc_hd__clkbuf_1 _16502_ (.A(_04488_),
    .X(_01792_));
 sky130_fd_sc_hd__buf_4 _16503_ (.A(_04466_),
    .X(_04489_));
 sky130_fd_sc_hd__mux2_1 _16504_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][11] ),
    .A1(_14463_),
    .S(_04489_),
    .X(_04490_));
 sky130_fd_sc_hd__clkbuf_1 _16505_ (.A(_04490_),
    .X(_01791_));
 sky130_fd_sc_hd__mux2_1 _16506_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][10] ),
    .A1(_14466_),
    .S(_04489_),
    .X(_04491_));
 sky130_fd_sc_hd__clkbuf_1 _16507_ (.A(_04491_),
    .X(_01790_));
 sky130_fd_sc_hd__mux2_1 _16508_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][9] ),
    .A1(_14468_),
    .S(_04489_),
    .X(_04492_));
 sky130_fd_sc_hd__clkbuf_1 _16509_ (.A(_04492_),
    .X(_01789_));
 sky130_fd_sc_hd__mux2_1 _16510_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][8] ),
    .A1(_14470_),
    .S(_04489_),
    .X(_04493_));
 sky130_fd_sc_hd__clkbuf_1 _16511_ (.A(_04493_),
    .X(_01788_));
 sky130_fd_sc_hd__mux2_1 _16512_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][7] ),
    .A1(_14472_),
    .S(_04489_),
    .X(_04494_));
 sky130_fd_sc_hd__clkbuf_1 _16513_ (.A(_04494_),
    .X(_01787_));
 sky130_fd_sc_hd__mux2_1 _16514_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][6] ),
    .A1(_14474_),
    .S(_04489_),
    .X(_04495_));
 sky130_fd_sc_hd__clkbuf_1 _16515_ (.A(_04495_),
    .X(_01786_));
 sky130_fd_sc_hd__mux2_1 _16516_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][5] ),
    .A1(_14476_),
    .S(_04489_),
    .X(_04496_));
 sky130_fd_sc_hd__clkbuf_1 _16517_ (.A(_04496_),
    .X(_01785_));
 sky130_fd_sc_hd__mux2_1 _16518_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][4] ),
    .A1(_14478_),
    .S(_04489_),
    .X(_04497_));
 sky130_fd_sc_hd__clkbuf_1 _16519_ (.A(_04497_),
    .X(_01784_));
 sky130_fd_sc_hd__mux2_1 _16520_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][3] ),
    .A1(_14480_),
    .S(_04489_),
    .X(_04498_));
 sky130_fd_sc_hd__clkbuf_1 _16521_ (.A(_04498_),
    .X(_01783_));
 sky130_fd_sc_hd__mux2_1 _16522_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][2] ),
    .A1(_14482_),
    .S(_04489_),
    .X(_04499_));
 sky130_fd_sc_hd__clkbuf_1 _16523_ (.A(_04499_),
    .X(_01782_));
 sky130_fd_sc_hd__mux2_1 _16524_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][1] ),
    .A1(_14484_),
    .S(_04466_),
    .X(_04500_));
 sky130_fd_sc_hd__clkbuf_1 _16525_ (.A(_04500_),
    .X(_01781_));
 sky130_fd_sc_hd__mux2_1 _16526_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][0] ),
    .A1(_14486_),
    .S(_04466_),
    .X(_04501_));
 sky130_fd_sc_hd__clkbuf_1 _16527_ (.A(_04501_),
    .X(_01780_));
 sky130_fd_sc_hd__nand2_4 _16528_ (.A(_14128_),
    .B(_04465_),
    .Y(_04502_));
 sky130_fd_sc_hd__clkbuf_4 _16529_ (.A(_04502_),
    .X(_04503_));
 sky130_fd_sc_hd__mux2_1 _16530_ (.A0(_14127_),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][31] ),
    .S(_04503_),
    .X(_04504_));
 sky130_fd_sc_hd__clkbuf_1 _16531_ (.A(_04504_),
    .X(_01779_));
 sky130_fd_sc_hd__mux2_1 _16532_ (.A0(_14133_),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][30] ),
    .S(_04503_),
    .X(_04505_));
 sky130_fd_sc_hd__clkbuf_1 _16533_ (.A(_04505_),
    .X(_01778_));
 sky130_fd_sc_hd__mux2_1 _16534_ (.A0(_14135_),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][29] ),
    .S(_04503_),
    .X(_04506_));
 sky130_fd_sc_hd__clkbuf_1 _16535_ (.A(_04506_),
    .X(_01777_));
 sky130_fd_sc_hd__mux2_1 _16536_ (.A0(_14137_),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][28] ),
    .S(_04503_),
    .X(_04507_));
 sky130_fd_sc_hd__clkbuf_1 _16537_ (.A(_04507_),
    .X(_01776_));
 sky130_fd_sc_hd__mux2_1 _16538_ (.A0(_14139_),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][27] ),
    .S(_04503_),
    .X(_04508_));
 sky130_fd_sc_hd__clkbuf_1 _16539_ (.A(_04508_),
    .X(_01775_));
 sky130_fd_sc_hd__mux2_1 _16540_ (.A0(_14141_),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][26] ),
    .S(_04503_),
    .X(_04509_));
 sky130_fd_sc_hd__clkbuf_1 _16541_ (.A(_04509_),
    .X(_01774_));
 sky130_fd_sc_hd__mux2_1 _16542_ (.A0(_14143_),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][25] ),
    .S(_04503_),
    .X(_04510_));
 sky130_fd_sc_hd__clkbuf_1 _16543_ (.A(_04510_),
    .X(_01773_));
 sky130_fd_sc_hd__mux2_1 _16544_ (.A0(_14145_),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][24] ),
    .S(_04503_),
    .X(_04511_));
 sky130_fd_sc_hd__clkbuf_1 _16545_ (.A(_04511_),
    .X(_01772_));
 sky130_fd_sc_hd__mux2_1 _16546_ (.A0(_14147_),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][23] ),
    .S(_04503_),
    .X(_04512_));
 sky130_fd_sc_hd__clkbuf_1 _16547_ (.A(_04512_),
    .X(_01771_));
 sky130_fd_sc_hd__mux2_1 _16548_ (.A0(_14149_),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][22] ),
    .S(_04503_),
    .X(_04513_));
 sky130_fd_sc_hd__clkbuf_1 _16549_ (.A(_04513_),
    .X(_01770_));
 sky130_fd_sc_hd__clkbuf_4 _16550_ (.A(_04502_),
    .X(_04514_));
 sky130_fd_sc_hd__mux2_1 _16551_ (.A0(_14151_),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][21] ),
    .S(_04514_),
    .X(_04515_));
 sky130_fd_sc_hd__clkbuf_1 _16552_ (.A(_04515_),
    .X(_01769_));
 sky130_fd_sc_hd__mux2_1 _16553_ (.A0(_14154_),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][20] ),
    .S(_04514_),
    .X(_04516_));
 sky130_fd_sc_hd__clkbuf_1 _16554_ (.A(_04516_),
    .X(_01768_));
 sky130_fd_sc_hd__mux2_1 _16555_ (.A0(_14156_),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][19] ),
    .S(_04514_),
    .X(_04517_));
 sky130_fd_sc_hd__clkbuf_1 _16556_ (.A(_04517_),
    .X(_01767_));
 sky130_fd_sc_hd__mux2_1 _16557_ (.A0(_14158_),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][18] ),
    .S(_04514_),
    .X(_04518_));
 sky130_fd_sc_hd__clkbuf_1 _16558_ (.A(_04518_),
    .X(_01766_));
 sky130_fd_sc_hd__mux2_1 _16559_ (.A0(_14160_),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][17] ),
    .S(_04514_),
    .X(_04519_));
 sky130_fd_sc_hd__clkbuf_1 _16560_ (.A(_04519_),
    .X(_01765_));
 sky130_fd_sc_hd__mux2_1 _16561_ (.A0(_14162_),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][16] ),
    .S(_04514_),
    .X(_04520_));
 sky130_fd_sc_hd__clkbuf_1 _16562_ (.A(_04520_),
    .X(_01764_));
 sky130_fd_sc_hd__mux2_1 _16563_ (.A0(_14164_),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][15] ),
    .S(_04514_),
    .X(_04521_));
 sky130_fd_sc_hd__clkbuf_1 _16564_ (.A(_04521_),
    .X(_01763_));
 sky130_fd_sc_hd__mux2_1 _16565_ (.A0(_14166_),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][14] ),
    .S(_04514_),
    .X(_04522_));
 sky130_fd_sc_hd__clkbuf_1 _16566_ (.A(_04522_),
    .X(_01762_));
 sky130_fd_sc_hd__mux2_1 _16567_ (.A0(_14168_),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][13] ),
    .S(_04514_),
    .X(_04523_));
 sky130_fd_sc_hd__clkbuf_1 _16568_ (.A(_04523_),
    .X(_01761_));
 sky130_fd_sc_hd__mux2_1 _16569_ (.A0(_14170_),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][12] ),
    .S(_04514_),
    .X(_04524_));
 sky130_fd_sc_hd__clkbuf_1 _16570_ (.A(_04524_),
    .X(_01760_));
 sky130_fd_sc_hd__clkbuf_4 _16571_ (.A(_04502_),
    .X(_04525_));
 sky130_fd_sc_hd__mux2_1 _16572_ (.A0(_14172_),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][11] ),
    .S(_04525_),
    .X(_04526_));
 sky130_fd_sc_hd__clkbuf_1 _16573_ (.A(_04526_),
    .X(_01759_));
 sky130_fd_sc_hd__mux2_1 _16574_ (.A0(_14175_),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][10] ),
    .S(_04525_),
    .X(_04527_));
 sky130_fd_sc_hd__clkbuf_1 _16575_ (.A(_04527_),
    .X(_01758_));
 sky130_fd_sc_hd__mux2_1 _16576_ (.A0(_14177_),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][9] ),
    .S(_04525_),
    .X(_04528_));
 sky130_fd_sc_hd__clkbuf_1 _16577_ (.A(_04528_),
    .X(_01757_));
 sky130_fd_sc_hd__mux2_1 _16578_ (.A0(_14179_),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][8] ),
    .S(_04525_),
    .X(_04529_));
 sky130_fd_sc_hd__clkbuf_1 _16579_ (.A(_04529_),
    .X(_01756_));
 sky130_fd_sc_hd__mux2_1 _16580_ (.A0(_14181_),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][7] ),
    .S(_04525_),
    .X(_04530_));
 sky130_fd_sc_hd__clkbuf_1 _16581_ (.A(_04530_),
    .X(_01755_));
 sky130_fd_sc_hd__mux2_1 _16582_ (.A0(_14183_),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][6] ),
    .S(_04525_),
    .X(_04531_));
 sky130_fd_sc_hd__clkbuf_1 _16583_ (.A(_04531_),
    .X(_01754_));
 sky130_fd_sc_hd__mux2_1 _16584_ (.A0(_14185_),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][5] ),
    .S(_04525_),
    .X(_04532_));
 sky130_fd_sc_hd__clkbuf_1 _16585_ (.A(_04532_),
    .X(_01753_));
 sky130_fd_sc_hd__mux2_1 _16586_ (.A0(_14187_),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][4] ),
    .S(_04525_),
    .X(_04533_));
 sky130_fd_sc_hd__clkbuf_1 _16587_ (.A(_04533_),
    .X(_01752_));
 sky130_fd_sc_hd__mux2_1 _16588_ (.A0(_14189_),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][3] ),
    .S(_04525_),
    .X(_04534_));
 sky130_fd_sc_hd__clkbuf_1 _16589_ (.A(_04534_),
    .X(_01751_));
 sky130_fd_sc_hd__mux2_1 _16590_ (.A0(_14191_),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][2] ),
    .S(_04525_),
    .X(_04535_));
 sky130_fd_sc_hd__clkbuf_1 _16591_ (.A(_04535_),
    .X(_01750_));
 sky130_fd_sc_hd__mux2_1 _16592_ (.A0(_14193_),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][1] ),
    .S(_04502_),
    .X(_04536_));
 sky130_fd_sc_hd__clkbuf_1 _16593_ (.A(_04536_),
    .X(_01749_));
 sky130_fd_sc_hd__mux2_1 _16594_ (.A0(_14195_),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][0] ),
    .S(_04502_),
    .X(_04537_));
 sky130_fd_sc_hd__clkbuf_1 _16595_ (.A(_04537_),
    .X(_01748_));
 sky130_fd_sc_hd__and3_4 _16596_ (.A(\rvcpu.dp.plmw.RegWriteW ),
    .B(_14346_),
    .C(\rvcpu.dp.plmw.RdW[1] ),
    .X(_04538_));
 sky130_fd_sc_hd__nand2_2 _16597_ (.A(_04538_),
    .B(_04465_),
    .Y(_04539_));
 sky130_fd_sc_hd__buf_4 _16598_ (.A(_04539_),
    .X(_04540_));
 sky130_fd_sc_hd__mux2_1 _16599_ (.A0(_14127_),
    .A1(\rvcpu.dp.rf.reg_file_arr[14][31] ),
    .S(_04540_),
    .X(_04541_));
 sky130_fd_sc_hd__clkbuf_1 _16600_ (.A(_04541_),
    .X(_01739_));
 sky130_fd_sc_hd__mux2_1 _16601_ (.A0(_14133_),
    .A1(\rvcpu.dp.rf.reg_file_arr[14][30] ),
    .S(_04540_),
    .X(_04542_));
 sky130_fd_sc_hd__clkbuf_1 _16602_ (.A(_04542_),
    .X(_01738_));
 sky130_fd_sc_hd__mux2_1 _16603_ (.A0(_14135_),
    .A1(\rvcpu.dp.rf.reg_file_arr[14][29] ),
    .S(_04540_),
    .X(_04543_));
 sky130_fd_sc_hd__clkbuf_1 _16604_ (.A(_04543_),
    .X(_01737_));
 sky130_fd_sc_hd__mux2_1 _16605_ (.A0(_14137_),
    .A1(\rvcpu.dp.rf.reg_file_arr[14][28] ),
    .S(_04540_),
    .X(_04544_));
 sky130_fd_sc_hd__clkbuf_1 _16606_ (.A(_04544_),
    .X(_01736_));
 sky130_fd_sc_hd__mux2_1 _16607_ (.A0(_14139_),
    .A1(\rvcpu.dp.rf.reg_file_arr[14][27] ),
    .S(_04540_),
    .X(_04545_));
 sky130_fd_sc_hd__clkbuf_1 _16608_ (.A(_04545_),
    .X(_01735_));
 sky130_fd_sc_hd__mux2_1 _16609_ (.A0(_14141_),
    .A1(\rvcpu.dp.rf.reg_file_arr[14][26] ),
    .S(_04540_),
    .X(_04546_));
 sky130_fd_sc_hd__clkbuf_1 _16610_ (.A(_04546_),
    .X(_01734_));
 sky130_fd_sc_hd__mux2_1 _16611_ (.A0(_14143_),
    .A1(\rvcpu.dp.rf.reg_file_arr[14][25] ),
    .S(_04540_),
    .X(_04547_));
 sky130_fd_sc_hd__clkbuf_1 _16612_ (.A(_04547_),
    .X(_01733_));
 sky130_fd_sc_hd__mux2_1 _16613_ (.A0(_14145_),
    .A1(\rvcpu.dp.rf.reg_file_arr[14][24] ),
    .S(_04540_),
    .X(_04548_));
 sky130_fd_sc_hd__clkbuf_1 _16614_ (.A(_04548_),
    .X(_01732_));
 sky130_fd_sc_hd__mux2_1 _16615_ (.A0(_14147_),
    .A1(\rvcpu.dp.rf.reg_file_arr[14][23] ),
    .S(_04540_),
    .X(_04549_));
 sky130_fd_sc_hd__clkbuf_1 _16616_ (.A(_04549_),
    .X(_01731_));
 sky130_fd_sc_hd__mux2_1 _16617_ (.A0(_14149_),
    .A1(\rvcpu.dp.rf.reg_file_arr[14][22] ),
    .S(_04540_),
    .X(_04550_));
 sky130_fd_sc_hd__clkbuf_1 _16618_ (.A(_04550_),
    .X(_01730_));
 sky130_fd_sc_hd__buf_4 _16619_ (.A(_04539_),
    .X(_04551_));
 sky130_fd_sc_hd__mux2_1 _16620_ (.A0(_14151_),
    .A1(\rvcpu.dp.rf.reg_file_arr[14][21] ),
    .S(_04551_),
    .X(_04552_));
 sky130_fd_sc_hd__clkbuf_1 _16621_ (.A(_04552_),
    .X(_01729_));
 sky130_fd_sc_hd__mux2_1 _16622_ (.A0(_14154_),
    .A1(\rvcpu.dp.rf.reg_file_arr[14][20] ),
    .S(_04551_),
    .X(_04553_));
 sky130_fd_sc_hd__clkbuf_1 _16623_ (.A(_04553_),
    .X(_01728_));
 sky130_fd_sc_hd__mux2_1 _16624_ (.A0(_14156_),
    .A1(\rvcpu.dp.rf.reg_file_arr[14][19] ),
    .S(_04551_),
    .X(_04554_));
 sky130_fd_sc_hd__clkbuf_1 _16625_ (.A(_04554_),
    .X(_01727_));
 sky130_fd_sc_hd__mux2_1 _16626_ (.A0(_14158_),
    .A1(\rvcpu.dp.rf.reg_file_arr[14][18] ),
    .S(_04551_),
    .X(_04555_));
 sky130_fd_sc_hd__clkbuf_1 _16627_ (.A(_04555_),
    .X(_01726_));
 sky130_fd_sc_hd__mux2_1 _16628_ (.A0(_14160_),
    .A1(\rvcpu.dp.rf.reg_file_arr[14][17] ),
    .S(_04551_),
    .X(_04556_));
 sky130_fd_sc_hd__clkbuf_1 _16629_ (.A(_04556_),
    .X(_01725_));
 sky130_fd_sc_hd__mux2_1 _16630_ (.A0(_14162_),
    .A1(\rvcpu.dp.rf.reg_file_arr[14][16] ),
    .S(_04551_),
    .X(_04557_));
 sky130_fd_sc_hd__clkbuf_1 _16631_ (.A(_04557_),
    .X(_01724_));
 sky130_fd_sc_hd__mux2_1 _16632_ (.A0(_14164_),
    .A1(\rvcpu.dp.rf.reg_file_arr[14][15] ),
    .S(_04551_),
    .X(_04558_));
 sky130_fd_sc_hd__clkbuf_1 _16633_ (.A(_04558_),
    .X(_01723_));
 sky130_fd_sc_hd__mux2_1 _16634_ (.A0(_14166_),
    .A1(\rvcpu.dp.rf.reg_file_arr[14][14] ),
    .S(_04551_),
    .X(_04559_));
 sky130_fd_sc_hd__clkbuf_1 _16635_ (.A(_04559_),
    .X(_01722_));
 sky130_fd_sc_hd__mux2_1 _16636_ (.A0(_14168_),
    .A1(\rvcpu.dp.rf.reg_file_arr[14][13] ),
    .S(_04551_),
    .X(_04560_));
 sky130_fd_sc_hd__clkbuf_1 _16637_ (.A(_04560_),
    .X(_01721_));
 sky130_fd_sc_hd__mux2_1 _16638_ (.A0(_14170_),
    .A1(\rvcpu.dp.rf.reg_file_arr[14][12] ),
    .S(_04551_),
    .X(_04561_));
 sky130_fd_sc_hd__clkbuf_1 _16639_ (.A(_04561_),
    .X(_01720_));
 sky130_fd_sc_hd__clkbuf_4 _16640_ (.A(_04539_),
    .X(_04562_));
 sky130_fd_sc_hd__mux2_1 _16641_ (.A0(_14172_),
    .A1(\rvcpu.dp.rf.reg_file_arr[14][11] ),
    .S(_04562_),
    .X(_04563_));
 sky130_fd_sc_hd__clkbuf_1 _16642_ (.A(_04563_),
    .X(_01719_));
 sky130_fd_sc_hd__mux2_1 _16643_ (.A0(_14175_),
    .A1(\rvcpu.dp.rf.reg_file_arr[14][10] ),
    .S(_04562_),
    .X(_04564_));
 sky130_fd_sc_hd__clkbuf_1 _16644_ (.A(_04564_),
    .X(_01718_));
 sky130_fd_sc_hd__mux2_1 _16645_ (.A0(_14177_),
    .A1(\rvcpu.dp.rf.reg_file_arr[14][9] ),
    .S(_04562_),
    .X(_04565_));
 sky130_fd_sc_hd__clkbuf_1 _16646_ (.A(_04565_),
    .X(_01717_));
 sky130_fd_sc_hd__mux2_1 _16647_ (.A0(_14179_),
    .A1(\rvcpu.dp.rf.reg_file_arr[14][8] ),
    .S(_04562_),
    .X(_04566_));
 sky130_fd_sc_hd__clkbuf_1 _16648_ (.A(_04566_),
    .X(_01716_));
 sky130_fd_sc_hd__mux2_1 _16649_ (.A0(_14181_),
    .A1(\rvcpu.dp.rf.reg_file_arr[14][7] ),
    .S(_04562_),
    .X(_04567_));
 sky130_fd_sc_hd__clkbuf_1 _16650_ (.A(_04567_),
    .X(_01715_));
 sky130_fd_sc_hd__mux2_1 _16651_ (.A0(_14183_),
    .A1(\rvcpu.dp.rf.reg_file_arr[14][6] ),
    .S(_04562_),
    .X(_04568_));
 sky130_fd_sc_hd__clkbuf_1 _16652_ (.A(_04568_),
    .X(_01714_));
 sky130_fd_sc_hd__mux2_1 _16653_ (.A0(_14185_),
    .A1(\rvcpu.dp.rf.reg_file_arr[14][5] ),
    .S(_04562_),
    .X(_04569_));
 sky130_fd_sc_hd__clkbuf_1 _16654_ (.A(_04569_),
    .X(_01713_));
 sky130_fd_sc_hd__mux2_1 _16655_ (.A0(_14187_),
    .A1(\rvcpu.dp.rf.reg_file_arr[14][4] ),
    .S(_04562_),
    .X(_04570_));
 sky130_fd_sc_hd__clkbuf_1 _16656_ (.A(_04570_),
    .X(_01712_));
 sky130_fd_sc_hd__mux2_1 _16657_ (.A0(_14189_),
    .A1(\rvcpu.dp.rf.reg_file_arr[14][3] ),
    .S(_04562_),
    .X(_04571_));
 sky130_fd_sc_hd__clkbuf_1 _16658_ (.A(_04571_),
    .X(_01711_));
 sky130_fd_sc_hd__mux2_1 _16659_ (.A0(_14191_),
    .A1(\rvcpu.dp.rf.reg_file_arr[14][2] ),
    .S(_04562_),
    .X(_04572_));
 sky130_fd_sc_hd__clkbuf_1 _16660_ (.A(_04572_),
    .X(_01710_));
 sky130_fd_sc_hd__mux2_1 _16661_ (.A0(_14193_),
    .A1(\rvcpu.dp.rf.reg_file_arr[14][1] ),
    .S(_04539_),
    .X(_04573_));
 sky130_fd_sc_hd__clkbuf_1 _16662_ (.A(_04573_),
    .X(_01709_));
 sky130_fd_sc_hd__mux2_1 _16663_ (.A0(_14195_),
    .A1(\rvcpu.dp.rf.reg_file_arr[14][0] ),
    .S(_04539_),
    .X(_04574_));
 sky130_fd_sc_hd__clkbuf_1 _16664_ (.A(_04574_),
    .X(_01708_));
 sky130_fd_sc_hd__nand2_2 _16665_ (.A(_14197_),
    .B(_04465_),
    .Y(_04575_));
 sky130_fd_sc_hd__clkbuf_4 _16666_ (.A(_04575_),
    .X(_04576_));
 sky130_fd_sc_hd__mux2_1 _16667_ (.A0(_14127_),
    .A1(\rvcpu.dp.rf.reg_file_arr[15][31] ),
    .S(_04576_),
    .X(_04577_));
 sky130_fd_sc_hd__clkbuf_1 _16668_ (.A(_04577_),
    .X(_01707_));
 sky130_fd_sc_hd__mux2_1 _16669_ (.A0(_14133_),
    .A1(\rvcpu.dp.rf.reg_file_arr[15][30] ),
    .S(_04576_),
    .X(_04578_));
 sky130_fd_sc_hd__clkbuf_1 _16670_ (.A(_04578_),
    .X(_01706_));
 sky130_fd_sc_hd__mux2_1 _16671_ (.A0(_14135_),
    .A1(\rvcpu.dp.rf.reg_file_arr[15][29] ),
    .S(_04576_),
    .X(_04579_));
 sky130_fd_sc_hd__clkbuf_1 _16672_ (.A(_04579_),
    .X(_01705_));
 sky130_fd_sc_hd__mux2_1 _16673_ (.A0(_14137_),
    .A1(\rvcpu.dp.rf.reg_file_arr[15][28] ),
    .S(_04576_),
    .X(_04580_));
 sky130_fd_sc_hd__clkbuf_1 _16674_ (.A(_04580_),
    .X(_01704_));
 sky130_fd_sc_hd__mux2_1 _16675_ (.A0(_14139_),
    .A1(\rvcpu.dp.rf.reg_file_arr[15][27] ),
    .S(_04576_),
    .X(_04581_));
 sky130_fd_sc_hd__clkbuf_1 _16676_ (.A(_04581_),
    .X(_01703_));
 sky130_fd_sc_hd__mux2_1 _16677_ (.A0(_14141_),
    .A1(\rvcpu.dp.rf.reg_file_arr[15][26] ),
    .S(_04576_),
    .X(_04582_));
 sky130_fd_sc_hd__clkbuf_1 _16678_ (.A(_04582_),
    .X(_01702_));
 sky130_fd_sc_hd__mux2_1 _16679_ (.A0(_14143_),
    .A1(\rvcpu.dp.rf.reg_file_arr[15][25] ),
    .S(_04576_),
    .X(_04583_));
 sky130_fd_sc_hd__clkbuf_1 _16680_ (.A(_04583_),
    .X(_01701_));
 sky130_fd_sc_hd__mux2_1 _16681_ (.A0(_14145_),
    .A1(\rvcpu.dp.rf.reg_file_arr[15][24] ),
    .S(_04576_),
    .X(_04584_));
 sky130_fd_sc_hd__clkbuf_1 _16682_ (.A(_04584_),
    .X(_01700_));
 sky130_fd_sc_hd__mux2_1 _16683_ (.A0(_14147_),
    .A1(\rvcpu.dp.rf.reg_file_arr[15][23] ),
    .S(_04576_),
    .X(_04585_));
 sky130_fd_sc_hd__clkbuf_1 _16684_ (.A(_04585_),
    .X(_01699_));
 sky130_fd_sc_hd__mux2_1 _16685_ (.A0(_14149_),
    .A1(\rvcpu.dp.rf.reg_file_arr[15][22] ),
    .S(_04576_),
    .X(_04586_));
 sky130_fd_sc_hd__clkbuf_1 _16686_ (.A(_04586_),
    .X(_01698_));
 sky130_fd_sc_hd__buf_4 _16687_ (.A(_04575_),
    .X(_04587_));
 sky130_fd_sc_hd__mux2_1 _16688_ (.A0(_14151_),
    .A1(\rvcpu.dp.rf.reg_file_arr[15][21] ),
    .S(_04587_),
    .X(_04588_));
 sky130_fd_sc_hd__clkbuf_1 _16689_ (.A(_04588_),
    .X(_01697_));
 sky130_fd_sc_hd__mux2_1 _16690_ (.A0(_14154_),
    .A1(\rvcpu.dp.rf.reg_file_arr[15][20] ),
    .S(_04587_),
    .X(_04589_));
 sky130_fd_sc_hd__clkbuf_1 _16691_ (.A(_04589_),
    .X(_01696_));
 sky130_fd_sc_hd__mux2_1 _16692_ (.A0(_14156_),
    .A1(\rvcpu.dp.rf.reg_file_arr[15][19] ),
    .S(_04587_),
    .X(_04590_));
 sky130_fd_sc_hd__clkbuf_1 _16693_ (.A(_04590_),
    .X(_01695_));
 sky130_fd_sc_hd__mux2_1 _16694_ (.A0(_14158_),
    .A1(\rvcpu.dp.rf.reg_file_arr[15][18] ),
    .S(_04587_),
    .X(_04591_));
 sky130_fd_sc_hd__clkbuf_1 _16695_ (.A(_04591_),
    .X(_01694_));
 sky130_fd_sc_hd__mux2_1 _16696_ (.A0(_14160_),
    .A1(\rvcpu.dp.rf.reg_file_arr[15][17] ),
    .S(_04587_),
    .X(_04592_));
 sky130_fd_sc_hd__clkbuf_1 _16697_ (.A(_04592_),
    .X(_01693_));
 sky130_fd_sc_hd__mux2_1 _16698_ (.A0(_14162_),
    .A1(\rvcpu.dp.rf.reg_file_arr[15][16] ),
    .S(_04587_),
    .X(_04593_));
 sky130_fd_sc_hd__clkbuf_1 _16699_ (.A(_04593_),
    .X(_01692_));
 sky130_fd_sc_hd__mux2_1 _16700_ (.A0(_14164_),
    .A1(\rvcpu.dp.rf.reg_file_arr[15][15] ),
    .S(_04587_),
    .X(_04594_));
 sky130_fd_sc_hd__clkbuf_1 _16701_ (.A(_04594_),
    .X(_01691_));
 sky130_fd_sc_hd__mux2_1 _16702_ (.A0(_14166_),
    .A1(\rvcpu.dp.rf.reg_file_arr[15][14] ),
    .S(_04587_),
    .X(_04595_));
 sky130_fd_sc_hd__clkbuf_1 _16703_ (.A(_04595_),
    .X(_01690_));
 sky130_fd_sc_hd__mux2_1 _16704_ (.A0(_14168_),
    .A1(\rvcpu.dp.rf.reg_file_arr[15][13] ),
    .S(_04587_),
    .X(_04596_));
 sky130_fd_sc_hd__clkbuf_1 _16705_ (.A(_04596_),
    .X(_01689_));
 sky130_fd_sc_hd__mux2_1 _16706_ (.A0(_14170_),
    .A1(\rvcpu.dp.rf.reg_file_arr[15][12] ),
    .S(_04587_),
    .X(_04597_));
 sky130_fd_sc_hd__clkbuf_1 _16707_ (.A(_04597_),
    .X(_01688_));
 sky130_fd_sc_hd__clkbuf_4 _16708_ (.A(_04575_),
    .X(_04598_));
 sky130_fd_sc_hd__mux2_1 _16709_ (.A0(_14172_),
    .A1(\rvcpu.dp.rf.reg_file_arr[15][11] ),
    .S(_04598_),
    .X(_04599_));
 sky130_fd_sc_hd__clkbuf_1 _16710_ (.A(_04599_),
    .X(_01687_));
 sky130_fd_sc_hd__mux2_1 _16711_ (.A0(_14175_),
    .A1(\rvcpu.dp.rf.reg_file_arr[15][10] ),
    .S(_04598_),
    .X(_04600_));
 sky130_fd_sc_hd__clkbuf_1 _16712_ (.A(_04600_),
    .X(_01686_));
 sky130_fd_sc_hd__mux2_1 _16713_ (.A0(_14177_),
    .A1(\rvcpu.dp.rf.reg_file_arr[15][9] ),
    .S(_04598_),
    .X(_04601_));
 sky130_fd_sc_hd__clkbuf_1 _16714_ (.A(_04601_),
    .X(_01685_));
 sky130_fd_sc_hd__mux2_1 _16715_ (.A0(_14179_),
    .A1(\rvcpu.dp.rf.reg_file_arr[15][8] ),
    .S(_04598_),
    .X(_04602_));
 sky130_fd_sc_hd__clkbuf_1 _16716_ (.A(_04602_),
    .X(_01684_));
 sky130_fd_sc_hd__mux2_1 _16717_ (.A0(_14181_),
    .A1(\rvcpu.dp.rf.reg_file_arr[15][7] ),
    .S(_04598_),
    .X(_04603_));
 sky130_fd_sc_hd__clkbuf_1 _16718_ (.A(_04603_),
    .X(_01683_));
 sky130_fd_sc_hd__mux2_1 _16719_ (.A0(_14183_),
    .A1(\rvcpu.dp.rf.reg_file_arr[15][6] ),
    .S(_04598_),
    .X(_04604_));
 sky130_fd_sc_hd__clkbuf_1 _16720_ (.A(_04604_),
    .X(_01682_));
 sky130_fd_sc_hd__mux2_1 _16721_ (.A0(_14185_),
    .A1(\rvcpu.dp.rf.reg_file_arr[15][5] ),
    .S(_04598_),
    .X(_04605_));
 sky130_fd_sc_hd__clkbuf_1 _16722_ (.A(_04605_),
    .X(_01681_));
 sky130_fd_sc_hd__mux2_1 _16723_ (.A0(_14187_),
    .A1(\rvcpu.dp.rf.reg_file_arr[15][4] ),
    .S(_04598_),
    .X(_04606_));
 sky130_fd_sc_hd__clkbuf_1 _16724_ (.A(_04606_),
    .X(_01680_));
 sky130_fd_sc_hd__mux2_1 _16725_ (.A0(_14189_),
    .A1(\rvcpu.dp.rf.reg_file_arr[15][3] ),
    .S(_04598_),
    .X(_04607_));
 sky130_fd_sc_hd__clkbuf_1 _16726_ (.A(_04607_),
    .X(_01679_));
 sky130_fd_sc_hd__mux2_1 _16727_ (.A0(_14191_),
    .A1(\rvcpu.dp.rf.reg_file_arr[15][2] ),
    .S(_04598_),
    .X(_04608_));
 sky130_fd_sc_hd__clkbuf_1 _16728_ (.A(_04608_),
    .X(_01678_));
 sky130_fd_sc_hd__mux2_1 _16729_ (.A0(_14193_),
    .A1(\rvcpu.dp.rf.reg_file_arr[15][1] ),
    .S(_04575_),
    .X(_04609_));
 sky130_fd_sc_hd__clkbuf_1 _16730_ (.A(_04609_),
    .X(_01677_));
 sky130_fd_sc_hd__mux2_1 _16731_ (.A0(_14195_),
    .A1(\rvcpu.dp.rf.reg_file_arr[15][0] ),
    .S(_04575_),
    .X(_04610_));
 sky130_fd_sc_hd__clkbuf_1 _16732_ (.A(_04610_),
    .X(_01676_));
 sky130_fd_sc_hd__nor2_2 _16733_ (.A(_14089_),
    .B(_14273_),
    .Y(_04611_));
 sky130_fd_sc_hd__clkbuf_4 _16734_ (.A(_04611_),
    .X(_04612_));
 sky130_fd_sc_hd__mux2_1 _16735_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][31] ),
    .A1(_14420_),
    .S(_04612_),
    .X(_04613_));
 sky130_fd_sc_hd__clkbuf_1 _16736_ (.A(_04613_),
    .X(_01675_));
 sky130_fd_sc_hd__mux2_1 _16737_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][30] ),
    .A1(_14424_),
    .S(_04612_),
    .X(_04614_));
 sky130_fd_sc_hd__clkbuf_1 _16738_ (.A(_04614_),
    .X(_01674_));
 sky130_fd_sc_hd__mux2_1 _16739_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][29] ),
    .A1(_14426_),
    .S(_04612_),
    .X(_04615_));
 sky130_fd_sc_hd__clkbuf_1 _16740_ (.A(_04615_),
    .X(_01673_));
 sky130_fd_sc_hd__mux2_1 _16741_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][28] ),
    .A1(_14428_),
    .S(_04612_),
    .X(_04616_));
 sky130_fd_sc_hd__clkbuf_1 _16742_ (.A(_04616_),
    .X(_01672_));
 sky130_fd_sc_hd__mux2_1 _16743_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][27] ),
    .A1(_14430_),
    .S(_04612_),
    .X(_04617_));
 sky130_fd_sc_hd__clkbuf_1 _16744_ (.A(_04617_),
    .X(_01671_));
 sky130_fd_sc_hd__mux2_1 _16745_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][26] ),
    .A1(_14432_),
    .S(_04612_),
    .X(_04618_));
 sky130_fd_sc_hd__clkbuf_1 _16746_ (.A(_04618_),
    .X(_01670_));
 sky130_fd_sc_hd__mux2_1 _16747_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][25] ),
    .A1(_14434_),
    .S(_04612_),
    .X(_04619_));
 sky130_fd_sc_hd__clkbuf_1 _16748_ (.A(_04619_),
    .X(_01669_));
 sky130_fd_sc_hd__mux2_1 _16749_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][24] ),
    .A1(_14436_),
    .S(_04612_),
    .X(_04620_));
 sky130_fd_sc_hd__clkbuf_1 _16750_ (.A(_04620_),
    .X(_01668_));
 sky130_fd_sc_hd__mux2_1 _16751_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][23] ),
    .A1(_14438_),
    .S(_04612_),
    .X(_04621_));
 sky130_fd_sc_hd__clkbuf_1 _16752_ (.A(_04621_),
    .X(_01667_));
 sky130_fd_sc_hd__mux2_1 _16753_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][22] ),
    .A1(_14440_),
    .S(_04612_),
    .X(_04622_));
 sky130_fd_sc_hd__clkbuf_1 _16754_ (.A(_04622_),
    .X(_01666_));
 sky130_fd_sc_hd__clkbuf_4 _16755_ (.A(_04611_),
    .X(_04623_));
 sky130_fd_sc_hd__mux2_1 _16756_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][21] ),
    .A1(_14442_),
    .S(_04623_),
    .X(_04624_));
 sky130_fd_sc_hd__clkbuf_1 _16757_ (.A(_04624_),
    .X(_01665_));
 sky130_fd_sc_hd__mux2_1 _16758_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][20] ),
    .A1(_14445_),
    .S(_04623_),
    .X(_04625_));
 sky130_fd_sc_hd__clkbuf_1 _16759_ (.A(_04625_),
    .X(_01664_));
 sky130_fd_sc_hd__mux2_1 _16760_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][19] ),
    .A1(_14447_),
    .S(_04623_),
    .X(_04626_));
 sky130_fd_sc_hd__clkbuf_1 _16761_ (.A(_04626_),
    .X(_01663_));
 sky130_fd_sc_hd__mux2_1 _16762_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][18] ),
    .A1(_14449_),
    .S(_04623_),
    .X(_04627_));
 sky130_fd_sc_hd__clkbuf_1 _16763_ (.A(_04627_),
    .X(_01662_));
 sky130_fd_sc_hd__mux2_1 _16764_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][17] ),
    .A1(_14451_),
    .S(_04623_),
    .X(_04628_));
 sky130_fd_sc_hd__clkbuf_1 _16765_ (.A(_04628_),
    .X(_01661_));
 sky130_fd_sc_hd__mux2_1 _16766_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][16] ),
    .A1(_14453_),
    .S(_04623_),
    .X(_04629_));
 sky130_fd_sc_hd__clkbuf_1 _16767_ (.A(_04629_),
    .X(_01660_));
 sky130_fd_sc_hd__mux2_1 _16768_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][15] ),
    .A1(_14455_),
    .S(_04623_),
    .X(_04630_));
 sky130_fd_sc_hd__clkbuf_1 _16769_ (.A(_04630_),
    .X(_01659_));
 sky130_fd_sc_hd__mux2_1 _16770_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][14] ),
    .A1(_14457_),
    .S(_04623_),
    .X(_04631_));
 sky130_fd_sc_hd__clkbuf_1 _16771_ (.A(_04631_),
    .X(_01658_));
 sky130_fd_sc_hd__mux2_1 _16772_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][13] ),
    .A1(_14459_),
    .S(_04623_),
    .X(_04632_));
 sky130_fd_sc_hd__clkbuf_1 _16773_ (.A(_04632_),
    .X(_01657_));
 sky130_fd_sc_hd__mux2_1 _16774_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][12] ),
    .A1(_14461_),
    .S(_04623_),
    .X(_04633_));
 sky130_fd_sc_hd__clkbuf_1 _16775_ (.A(_04633_),
    .X(_01656_));
 sky130_fd_sc_hd__buf_4 _16776_ (.A(_04611_),
    .X(_04634_));
 sky130_fd_sc_hd__mux2_1 _16777_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][11] ),
    .A1(_14463_),
    .S(_04634_),
    .X(_04635_));
 sky130_fd_sc_hd__clkbuf_1 _16778_ (.A(_04635_),
    .X(_01655_));
 sky130_fd_sc_hd__mux2_1 _16779_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][10] ),
    .A1(_14466_),
    .S(_04634_),
    .X(_04636_));
 sky130_fd_sc_hd__clkbuf_1 _16780_ (.A(_04636_),
    .X(_01654_));
 sky130_fd_sc_hd__mux2_1 _16781_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][9] ),
    .A1(_14468_),
    .S(_04634_),
    .X(_04637_));
 sky130_fd_sc_hd__clkbuf_1 _16782_ (.A(_04637_),
    .X(_01653_));
 sky130_fd_sc_hd__mux2_1 _16783_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][8] ),
    .A1(_14470_),
    .S(_04634_),
    .X(_04638_));
 sky130_fd_sc_hd__clkbuf_1 _16784_ (.A(_04638_),
    .X(_01652_));
 sky130_fd_sc_hd__mux2_1 _16785_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][7] ),
    .A1(_14472_),
    .S(_04634_),
    .X(_04639_));
 sky130_fd_sc_hd__clkbuf_1 _16786_ (.A(_04639_),
    .X(_01651_));
 sky130_fd_sc_hd__mux2_1 _16787_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][6] ),
    .A1(_14474_),
    .S(_04634_),
    .X(_04640_));
 sky130_fd_sc_hd__clkbuf_1 _16788_ (.A(_04640_),
    .X(_01650_));
 sky130_fd_sc_hd__mux2_1 _16789_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][5] ),
    .A1(_14476_),
    .S(_04634_),
    .X(_04641_));
 sky130_fd_sc_hd__clkbuf_1 _16790_ (.A(_04641_),
    .X(_01649_));
 sky130_fd_sc_hd__mux2_1 _16791_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][4] ),
    .A1(_14478_),
    .S(_04634_),
    .X(_04642_));
 sky130_fd_sc_hd__clkbuf_1 _16792_ (.A(_04642_),
    .X(_01648_));
 sky130_fd_sc_hd__mux2_1 _16793_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][3] ),
    .A1(_14480_),
    .S(_04634_),
    .X(_04643_));
 sky130_fd_sc_hd__clkbuf_1 _16794_ (.A(_04643_),
    .X(_01647_));
 sky130_fd_sc_hd__mux2_1 _16795_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][2] ),
    .A1(_14482_),
    .S(_04634_),
    .X(_04644_));
 sky130_fd_sc_hd__clkbuf_1 _16796_ (.A(_04644_),
    .X(_01646_));
 sky130_fd_sc_hd__mux2_1 _16797_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][1] ),
    .A1(_14484_),
    .S(_04611_),
    .X(_04645_));
 sky130_fd_sc_hd__clkbuf_1 _16798_ (.A(_04645_),
    .X(_01645_));
 sky130_fd_sc_hd__mux2_1 _16799_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][0] ),
    .A1(_14486_),
    .S(_04611_),
    .X(_04646_));
 sky130_fd_sc_hd__clkbuf_1 _16800_ (.A(_04646_),
    .X(_01644_));
 sky130_fd_sc_hd__nor2_2 _16801_ (.A(_13179_),
    .B(_14089_),
    .Y(_04647_));
 sky130_fd_sc_hd__buf_4 _16802_ (.A(_04647_),
    .X(_04648_));
 sky130_fd_sc_hd__mux2_1 _16803_ (.A0(\rvcpu.dp.rf.reg_file_arr[17][31] ),
    .A1(_14420_),
    .S(_04648_),
    .X(_04649_));
 sky130_fd_sc_hd__clkbuf_1 _16804_ (.A(_04649_),
    .X(_01635_));
 sky130_fd_sc_hd__mux2_1 _16805_ (.A0(\rvcpu.dp.rf.reg_file_arr[17][30] ),
    .A1(_14424_),
    .S(_04648_),
    .X(_04650_));
 sky130_fd_sc_hd__clkbuf_1 _16806_ (.A(_04650_),
    .X(_01634_));
 sky130_fd_sc_hd__mux2_1 _16807_ (.A0(\rvcpu.dp.rf.reg_file_arr[17][29] ),
    .A1(_14426_),
    .S(_04648_),
    .X(_04651_));
 sky130_fd_sc_hd__clkbuf_1 _16808_ (.A(_04651_),
    .X(_01633_));
 sky130_fd_sc_hd__mux2_1 _16809_ (.A0(\rvcpu.dp.rf.reg_file_arr[17][28] ),
    .A1(_14428_),
    .S(_04648_),
    .X(_04652_));
 sky130_fd_sc_hd__clkbuf_1 _16810_ (.A(_04652_),
    .X(_01632_));
 sky130_fd_sc_hd__mux2_1 _16811_ (.A0(\rvcpu.dp.rf.reg_file_arr[17][27] ),
    .A1(_14430_),
    .S(_04648_),
    .X(_04653_));
 sky130_fd_sc_hd__clkbuf_1 _16812_ (.A(_04653_),
    .X(_01631_));
 sky130_fd_sc_hd__mux2_1 _16813_ (.A0(\rvcpu.dp.rf.reg_file_arr[17][26] ),
    .A1(_14432_),
    .S(_04648_),
    .X(_04654_));
 sky130_fd_sc_hd__clkbuf_1 _16814_ (.A(_04654_),
    .X(_01630_));
 sky130_fd_sc_hd__mux2_1 _16815_ (.A0(\rvcpu.dp.rf.reg_file_arr[17][25] ),
    .A1(_14434_),
    .S(_04648_),
    .X(_04655_));
 sky130_fd_sc_hd__clkbuf_1 _16816_ (.A(_04655_),
    .X(_01629_));
 sky130_fd_sc_hd__mux2_1 _16817_ (.A0(\rvcpu.dp.rf.reg_file_arr[17][24] ),
    .A1(_14436_),
    .S(_04648_),
    .X(_04656_));
 sky130_fd_sc_hd__clkbuf_1 _16818_ (.A(_04656_),
    .X(_01628_));
 sky130_fd_sc_hd__mux2_1 _16819_ (.A0(\rvcpu.dp.rf.reg_file_arr[17][23] ),
    .A1(_14438_),
    .S(_04648_),
    .X(_04657_));
 sky130_fd_sc_hd__clkbuf_1 _16820_ (.A(_04657_),
    .X(_01627_));
 sky130_fd_sc_hd__mux2_1 _16821_ (.A0(\rvcpu.dp.rf.reg_file_arr[17][22] ),
    .A1(_14440_),
    .S(_04648_),
    .X(_04658_));
 sky130_fd_sc_hd__clkbuf_1 _16822_ (.A(_04658_),
    .X(_01626_));
 sky130_fd_sc_hd__buf_4 _16823_ (.A(_04647_),
    .X(_04659_));
 sky130_fd_sc_hd__mux2_1 _16824_ (.A0(\rvcpu.dp.rf.reg_file_arr[17][21] ),
    .A1(_14442_),
    .S(_04659_),
    .X(_04660_));
 sky130_fd_sc_hd__clkbuf_1 _16825_ (.A(_04660_),
    .X(_01625_));
 sky130_fd_sc_hd__mux2_1 _16826_ (.A0(\rvcpu.dp.rf.reg_file_arr[17][20] ),
    .A1(_14445_),
    .S(_04659_),
    .X(_04661_));
 sky130_fd_sc_hd__clkbuf_1 _16827_ (.A(_04661_),
    .X(_01624_));
 sky130_fd_sc_hd__mux2_1 _16828_ (.A0(\rvcpu.dp.rf.reg_file_arr[17][19] ),
    .A1(_14447_),
    .S(_04659_),
    .X(_04662_));
 sky130_fd_sc_hd__clkbuf_1 _16829_ (.A(_04662_),
    .X(_01623_));
 sky130_fd_sc_hd__mux2_1 _16830_ (.A0(\rvcpu.dp.rf.reg_file_arr[17][18] ),
    .A1(_14449_),
    .S(_04659_),
    .X(_04663_));
 sky130_fd_sc_hd__clkbuf_1 _16831_ (.A(_04663_),
    .X(_01622_));
 sky130_fd_sc_hd__mux2_1 _16832_ (.A0(\rvcpu.dp.rf.reg_file_arr[17][17] ),
    .A1(_14451_),
    .S(_04659_),
    .X(_04664_));
 sky130_fd_sc_hd__clkbuf_1 _16833_ (.A(_04664_),
    .X(_01621_));
 sky130_fd_sc_hd__mux2_1 _16834_ (.A0(\rvcpu.dp.rf.reg_file_arr[17][16] ),
    .A1(_14453_),
    .S(_04659_),
    .X(_04665_));
 sky130_fd_sc_hd__clkbuf_1 _16835_ (.A(_04665_),
    .X(_01620_));
 sky130_fd_sc_hd__mux2_1 _16836_ (.A0(\rvcpu.dp.rf.reg_file_arr[17][15] ),
    .A1(_14455_),
    .S(_04659_),
    .X(_04666_));
 sky130_fd_sc_hd__clkbuf_1 _16837_ (.A(_04666_),
    .X(_01619_));
 sky130_fd_sc_hd__mux2_1 _16838_ (.A0(\rvcpu.dp.rf.reg_file_arr[17][14] ),
    .A1(_14457_),
    .S(_04659_),
    .X(_04667_));
 sky130_fd_sc_hd__clkbuf_1 _16839_ (.A(_04667_),
    .X(_01618_));
 sky130_fd_sc_hd__mux2_1 _16840_ (.A0(\rvcpu.dp.rf.reg_file_arr[17][13] ),
    .A1(_14459_),
    .S(_04659_),
    .X(_04668_));
 sky130_fd_sc_hd__clkbuf_1 _16841_ (.A(_04668_),
    .X(_01617_));
 sky130_fd_sc_hd__mux2_1 _16842_ (.A0(\rvcpu.dp.rf.reg_file_arr[17][12] ),
    .A1(_14461_),
    .S(_04659_),
    .X(_04669_));
 sky130_fd_sc_hd__clkbuf_1 _16843_ (.A(_04669_),
    .X(_01616_));
 sky130_fd_sc_hd__buf_4 _16844_ (.A(_04647_),
    .X(_04670_));
 sky130_fd_sc_hd__mux2_1 _16845_ (.A0(\rvcpu.dp.rf.reg_file_arr[17][11] ),
    .A1(_14463_),
    .S(_04670_),
    .X(_04671_));
 sky130_fd_sc_hd__clkbuf_1 _16846_ (.A(_04671_),
    .X(_01615_));
 sky130_fd_sc_hd__mux2_1 _16847_ (.A0(\rvcpu.dp.rf.reg_file_arr[17][10] ),
    .A1(_14466_),
    .S(_04670_),
    .X(_04672_));
 sky130_fd_sc_hd__clkbuf_1 _16848_ (.A(_04672_),
    .X(_01614_));
 sky130_fd_sc_hd__mux2_1 _16849_ (.A0(\rvcpu.dp.rf.reg_file_arr[17][9] ),
    .A1(_14468_),
    .S(_04670_),
    .X(_04673_));
 sky130_fd_sc_hd__clkbuf_1 _16850_ (.A(_04673_),
    .X(_01613_));
 sky130_fd_sc_hd__mux2_1 _16851_ (.A0(\rvcpu.dp.rf.reg_file_arr[17][8] ),
    .A1(_14470_),
    .S(_04670_),
    .X(_04674_));
 sky130_fd_sc_hd__clkbuf_1 _16852_ (.A(_04674_),
    .X(_01612_));
 sky130_fd_sc_hd__mux2_1 _16853_ (.A0(\rvcpu.dp.rf.reg_file_arr[17][7] ),
    .A1(_14472_),
    .S(_04670_),
    .X(_04675_));
 sky130_fd_sc_hd__clkbuf_1 _16854_ (.A(_04675_),
    .X(_01611_));
 sky130_fd_sc_hd__mux2_1 _16855_ (.A0(\rvcpu.dp.rf.reg_file_arr[17][6] ),
    .A1(_14474_),
    .S(_04670_),
    .X(_04676_));
 sky130_fd_sc_hd__clkbuf_1 _16856_ (.A(_04676_),
    .X(_01610_));
 sky130_fd_sc_hd__mux2_1 _16857_ (.A0(\rvcpu.dp.rf.reg_file_arr[17][5] ),
    .A1(_14476_),
    .S(_04670_),
    .X(_04677_));
 sky130_fd_sc_hd__clkbuf_1 _16858_ (.A(_04677_),
    .X(_01609_));
 sky130_fd_sc_hd__mux2_1 _16859_ (.A0(\rvcpu.dp.rf.reg_file_arr[17][4] ),
    .A1(_14478_),
    .S(_04670_),
    .X(_04678_));
 sky130_fd_sc_hd__clkbuf_1 _16860_ (.A(_04678_),
    .X(_01608_));
 sky130_fd_sc_hd__mux2_1 _16861_ (.A0(\rvcpu.dp.rf.reg_file_arr[17][3] ),
    .A1(_14480_),
    .S(_04670_),
    .X(_04679_));
 sky130_fd_sc_hd__clkbuf_1 _16862_ (.A(_04679_),
    .X(_01607_));
 sky130_fd_sc_hd__mux2_1 _16863_ (.A0(\rvcpu.dp.rf.reg_file_arr[17][2] ),
    .A1(_14482_),
    .S(_04670_),
    .X(_04680_));
 sky130_fd_sc_hd__clkbuf_1 _16864_ (.A(_04680_),
    .X(_01606_));
 sky130_fd_sc_hd__mux2_1 _16865_ (.A0(\rvcpu.dp.rf.reg_file_arr[17][1] ),
    .A1(_14484_),
    .S(_04647_),
    .X(_04681_));
 sky130_fd_sc_hd__clkbuf_1 _16866_ (.A(_04681_),
    .X(_01605_));
 sky130_fd_sc_hd__mux2_1 _16867_ (.A0(\rvcpu.dp.rf.reg_file_arr[17][0] ),
    .A1(_14486_),
    .S(_04647_),
    .X(_04682_));
 sky130_fd_sc_hd__clkbuf_1 _16868_ (.A(_04682_),
    .X(_01604_));
 sky130_fd_sc_hd__nor2_2 _16869_ (.A(_14089_),
    .B(_14347_),
    .Y(_04683_));
 sky130_fd_sc_hd__clkbuf_4 _16870_ (.A(_04683_),
    .X(_04684_));
 sky130_fd_sc_hd__mux2_1 _16871_ (.A0(\rvcpu.dp.rf.reg_file_arr[18][31] ),
    .A1(_14420_),
    .S(_04684_),
    .X(_04685_));
 sky130_fd_sc_hd__clkbuf_1 _16872_ (.A(_04685_),
    .X(_01603_));
 sky130_fd_sc_hd__mux2_1 _16873_ (.A0(\rvcpu.dp.rf.reg_file_arr[18][30] ),
    .A1(_14424_),
    .S(_04684_),
    .X(_04686_));
 sky130_fd_sc_hd__clkbuf_1 _16874_ (.A(_04686_),
    .X(_01602_));
 sky130_fd_sc_hd__mux2_1 _16875_ (.A0(\rvcpu.dp.rf.reg_file_arr[18][29] ),
    .A1(_14426_),
    .S(_04684_),
    .X(_04687_));
 sky130_fd_sc_hd__clkbuf_1 _16876_ (.A(_04687_),
    .X(_01601_));
 sky130_fd_sc_hd__mux2_1 _16877_ (.A0(\rvcpu.dp.rf.reg_file_arr[18][28] ),
    .A1(_14428_),
    .S(_04684_),
    .X(_04688_));
 sky130_fd_sc_hd__clkbuf_1 _16878_ (.A(_04688_),
    .X(_01600_));
 sky130_fd_sc_hd__mux2_1 _16879_ (.A0(\rvcpu.dp.rf.reg_file_arr[18][27] ),
    .A1(_14430_),
    .S(_04684_),
    .X(_04689_));
 sky130_fd_sc_hd__clkbuf_1 _16880_ (.A(_04689_),
    .X(_01599_));
 sky130_fd_sc_hd__mux2_1 _16881_ (.A0(\rvcpu.dp.rf.reg_file_arr[18][26] ),
    .A1(_14432_),
    .S(_04684_),
    .X(_04690_));
 sky130_fd_sc_hd__clkbuf_1 _16882_ (.A(_04690_),
    .X(_01598_));
 sky130_fd_sc_hd__mux2_1 _16883_ (.A0(\rvcpu.dp.rf.reg_file_arr[18][25] ),
    .A1(_14434_),
    .S(_04684_),
    .X(_04691_));
 sky130_fd_sc_hd__clkbuf_1 _16884_ (.A(_04691_),
    .X(_01597_));
 sky130_fd_sc_hd__mux2_1 _16885_ (.A0(\rvcpu.dp.rf.reg_file_arr[18][24] ),
    .A1(_14436_),
    .S(_04684_),
    .X(_04692_));
 sky130_fd_sc_hd__clkbuf_1 _16886_ (.A(_04692_),
    .X(_01596_));
 sky130_fd_sc_hd__mux2_1 _16887_ (.A0(\rvcpu.dp.rf.reg_file_arr[18][23] ),
    .A1(_14438_),
    .S(_04684_),
    .X(_04693_));
 sky130_fd_sc_hd__clkbuf_1 _16888_ (.A(_04693_),
    .X(_01595_));
 sky130_fd_sc_hd__mux2_1 _16889_ (.A0(\rvcpu.dp.rf.reg_file_arr[18][22] ),
    .A1(_14440_),
    .S(_04684_),
    .X(_04694_));
 sky130_fd_sc_hd__clkbuf_1 _16890_ (.A(_04694_),
    .X(_01594_));
 sky130_fd_sc_hd__buf_4 _16891_ (.A(_04683_),
    .X(_04695_));
 sky130_fd_sc_hd__mux2_1 _16892_ (.A0(\rvcpu.dp.rf.reg_file_arr[18][21] ),
    .A1(_14442_),
    .S(_04695_),
    .X(_04696_));
 sky130_fd_sc_hd__clkbuf_1 _16893_ (.A(_04696_),
    .X(_01593_));
 sky130_fd_sc_hd__mux2_1 _16894_ (.A0(\rvcpu.dp.rf.reg_file_arr[18][20] ),
    .A1(_14445_),
    .S(_04695_),
    .X(_04697_));
 sky130_fd_sc_hd__clkbuf_1 _16895_ (.A(_04697_),
    .X(_01592_));
 sky130_fd_sc_hd__mux2_1 _16896_ (.A0(\rvcpu.dp.rf.reg_file_arr[18][19] ),
    .A1(_14447_),
    .S(_04695_),
    .X(_04698_));
 sky130_fd_sc_hd__clkbuf_1 _16897_ (.A(_04698_),
    .X(_01591_));
 sky130_fd_sc_hd__mux2_1 _16898_ (.A0(\rvcpu.dp.rf.reg_file_arr[18][18] ),
    .A1(_14449_),
    .S(_04695_),
    .X(_04699_));
 sky130_fd_sc_hd__clkbuf_1 _16899_ (.A(_04699_),
    .X(_01590_));
 sky130_fd_sc_hd__mux2_1 _16900_ (.A0(\rvcpu.dp.rf.reg_file_arr[18][17] ),
    .A1(_14451_),
    .S(_04695_),
    .X(_04700_));
 sky130_fd_sc_hd__clkbuf_1 _16901_ (.A(_04700_),
    .X(_01589_));
 sky130_fd_sc_hd__mux2_1 _16902_ (.A0(\rvcpu.dp.rf.reg_file_arr[18][16] ),
    .A1(_14453_),
    .S(_04695_),
    .X(_04701_));
 sky130_fd_sc_hd__clkbuf_1 _16903_ (.A(_04701_),
    .X(_01588_));
 sky130_fd_sc_hd__mux2_1 _16904_ (.A0(\rvcpu.dp.rf.reg_file_arr[18][15] ),
    .A1(_14455_),
    .S(_04695_),
    .X(_04702_));
 sky130_fd_sc_hd__clkbuf_1 _16905_ (.A(_04702_),
    .X(_01587_));
 sky130_fd_sc_hd__mux2_1 _16906_ (.A0(\rvcpu.dp.rf.reg_file_arr[18][14] ),
    .A1(_14457_),
    .S(_04695_),
    .X(_04703_));
 sky130_fd_sc_hd__clkbuf_1 _16907_ (.A(_04703_),
    .X(_01586_));
 sky130_fd_sc_hd__mux2_1 _16908_ (.A0(\rvcpu.dp.rf.reg_file_arr[18][13] ),
    .A1(_14459_),
    .S(_04695_),
    .X(_04704_));
 sky130_fd_sc_hd__clkbuf_1 _16909_ (.A(_04704_),
    .X(_01585_));
 sky130_fd_sc_hd__mux2_1 _16910_ (.A0(\rvcpu.dp.rf.reg_file_arr[18][12] ),
    .A1(_14461_),
    .S(_04695_),
    .X(_04705_));
 sky130_fd_sc_hd__clkbuf_1 _16911_ (.A(_04705_),
    .X(_01584_));
 sky130_fd_sc_hd__buf_4 _16912_ (.A(_04683_),
    .X(_04706_));
 sky130_fd_sc_hd__mux2_1 _16913_ (.A0(\rvcpu.dp.rf.reg_file_arr[18][11] ),
    .A1(_14463_),
    .S(_04706_),
    .X(_04707_));
 sky130_fd_sc_hd__clkbuf_1 _16914_ (.A(_04707_),
    .X(_01583_));
 sky130_fd_sc_hd__mux2_1 _16915_ (.A0(\rvcpu.dp.rf.reg_file_arr[18][10] ),
    .A1(_14466_),
    .S(_04706_),
    .X(_04708_));
 sky130_fd_sc_hd__clkbuf_1 _16916_ (.A(_04708_),
    .X(_01582_));
 sky130_fd_sc_hd__mux2_1 _16917_ (.A0(\rvcpu.dp.rf.reg_file_arr[18][9] ),
    .A1(_14468_),
    .S(_04706_),
    .X(_04709_));
 sky130_fd_sc_hd__clkbuf_1 _16918_ (.A(_04709_),
    .X(_01581_));
 sky130_fd_sc_hd__mux2_1 _16919_ (.A0(\rvcpu.dp.rf.reg_file_arr[18][8] ),
    .A1(_14470_),
    .S(_04706_),
    .X(_04710_));
 sky130_fd_sc_hd__clkbuf_1 _16920_ (.A(_04710_),
    .X(_01580_));
 sky130_fd_sc_hd__mux2_1 _16921_ (.A0(\rvcpu.dp.rf.reg_file_arr[18][7] ),
    .A1(_14472_),
    .S(_04706_),
    .X(_04711_));
 sky130_fd_sc_hd__clkbuf_1 _16922_ (.A(_04711_),
    .X(_01579_));
 sky130_fd_sc_hd__mux2_1 _16923_ (.A0(\rvcpu.dp.rf.reg_file_arr[18][6] ),
    .A1(_14474_),
    .S(_04706_),
    .X(_04712_));
 sky130_fd_sc_hd__clkbuf_1 _16924_ (.A(_04712_),
    .X(_01578_));
 sky130_fd_sc_hd__mux2_1 _16925_ (.A0(\rvcpu.dp.rf.reg_file_arr[18][5] ),
    .A1(_14476_),
    .S(_04706_),
    .X(_04713_));
 sky130_fd_sc_hd__clkbuf_1 _16926_ (.A(_04713_),
    .X(_01577_));
 sky130_fd_sc_hd__mux2_1 _16927_ (.A0(\rvcpu.dp.rf.reg_file_arr[18][4] ),
    .A1(_14478_),
    .S(_04706_),
    .X(_04714_));
 sky130_fd_sc_hd__clkbuf_1 _16928_ (.A(_04714_),
    .X(_01576_));
 sky130_fd_sc_hd__mux2_1 _16929_ (.A0(\rvcpu.dp.rf.reg_file_arr[18][3] ),
    .A1(_14480_),
    .S(_04706_),
    .X(_04715_));
 sky130_fd_sc_hd__clkbuf_1 _16930_ (.A(_04715_),
    .X(_01575_));
 sky130_fd_sc_hd__mux2_1 _16931_ (.A0(\rvcpu.dp.rf.reg_file_arr[18][2] ),
    .A1(_14482_),
    .S(_04706_),
    .X(_04716_));
 sky130_fd_sc_hd__clkbuf_1 _16932_ (.A(_04716_),
    .X(_01574_));
 sky130_fd_sc_hd__mux2_1 _16933_ (.A0(\rvcpu.dp.rf.reg_file_arr[18][1] ),
    .A1(_14484_),
    .S(_04683_),
    .X(_04717_));
 sky130_fd_sc_hd__clkbuf_1 _16934_ (.A(_04717_),
    .X(_01573_));
 sky130_fd_sc_hd__mux2_1 _16935_ (.A0(\rvcpu.dp.rf.reg_file_arr[18][0] ),
    .A1(_14486_),
    .S(_04683_),
    .X(_04718_));
 sky130_fd_sc_hd__clkbuf_1 _16936_ (.A(_04718_),
    .X(_01572_));
 sky130_fd_sc_hd__nor2_2 _16937_ (.A(_13179_),
    .B(_14234_),
    .Y(_04719_));
 sky130_fd_sc_hd__buf_4 _16938_ (.A(_04719_),
    .X(_04720_));
 sky130_fd_sc_hd__mux2_1 _16939_ (.A0(\rvcpu.dp.rf.reg_file_arr[1][31] ),
    .A1(_14420_),
    .S(_04720_),
    .X(_04721_));
 sky130_fd_sc_hd__clkbuf_1 _16940_ (.A(_04721_),
    .X(_01571_));
 sky130_fd_sc_hd__mux2_1 _16941_ (.A0(\rvcpu.dp.rf.reg_file_arr[1][30] ),
    .A1(_14424_),
    .S(_04720_),
    .X(_04722_));
 sky130_fd_sc_hd__clkbuf_1 _16942_ (.A(_04722_),
    .X(_01570_));
 sky130_fd_sc_hd__mux2_1 _16943_ (.A0(\rvcpu.dp.rf.reg_file_arr[1][29] ),
    .A1(_14426_),
    .S(_04720_),
    .X(_04723_));
 sky130_fd_sc_hd__clkbuf_1 _16944_ (.A(_04723_),
    .X(_01569_));
 sky130_fd_sc_hd__mux2_1 _16945_ (.A0(\rvcpu.dp.rf.reg_file_arr[1][28] ),
    .A1(_14428_),
    .S(_04720_),
    .X(_04724_));
 sky130_fd_sc_hd__clkbuf_1 _16946_ (.A(_04724_),
    .X(_01568_));
 sky130_fd_sc_hd__mux2_1 _16947_ (.A0(\rvcpu.dp.rf.reg_file_arr[1][27] ),
    .A1(_14430_),
    .S(_04720_),
    .X(_04725_));
 sky130_fd_sc_hd__clkbuf_1 _16948_ (.A(_04725_),
    .X(_01567_));
 sky130_fd_sc_hd__mux2_1 _16949_ (.A0(\rvcpu.dp.rf.reg_file_arr[1][26] ),
    .A1(_14432_),
    .S(_04720_),
    .X(_04726_));
 sky130_fd_sc_hd__clkbuf_1 _16950_ (.A(_04726_),
    .X(_01566_));
 sky130_fd_sc_hd__mux2_1 _16951_ (.A0(\rvcpu.dp.rf.reg_file_arr[1][25] ),
    .A1(_14434_),
    .S(_04720_),
    .X(_04727_));
 sky130_fd_sc_hd__clkbuf_1 _16952_ (.A(_04727_),
    .X(_01565_));
 sky130_fd_sc_hd__mux2_1 _16953_ (.A0(\rvcpu.dp.rf.reg_file_arr[1][24] ),
    .A1(_14436_),
    .S(_04720_),
    .X(_04728_));
 sky130_fd_sc_hd__clkbuf_1 _16954_ (.A(_04728_),
    .X(_01564_));
 sky130_fd_sc_hd__mux2_1 _16955_ (.A0(\rvcpu.dp.rf.reg_file_arr[1][23] ),
    .A1(_14438_),
    .S(_04720_),
    .X(_04729_));
 sky130_fd_sc_hd__clkbuf_1 _16956_ (.A(_04729_),
    .X(_01563_));
 sky130_fd_sc_hd__mux2_1 _16957_ (.A0(\rvcpu.dp.rf.reg_file_arr[1][22] ),
    .A1(_14440_),
    .S(_04720_),
    .X(_04730_));
 sky130_fd_sc_hd__clkbuf_1 _16958_ (.A(_04730_),
    .X(_01562_));
 sky130_fd_sc_hd__buf_4 _16959_ (.A(_04719_),
    .X(_04731_));
 sky130_fd_sc_hd__mux2_1 _16960_ (.A0(\rvcpu.dp.rf.reg_file_arr[1][21] ),
    .A1(_14442_),
    .S(_04731_),
    .X(_04732_));
 sky130_fd_sc_hd__clkbuf_1 _16961_ (.A(_04732_),
    .X(_01561_));
 sky130_fd_sc_hd__mux2_1 _16962_ (.A0(\rvcpu.dp.rf.reg_file_arr[1][20] ),
    .A1(_14445_),
    .S(_04731_),
    .X(_04733_));
 sky130_fd_sc_hd__clkbuf_1 _16963_ (.A(_04733_),
    .X(_01560_));
 sky130_fd_sc_hd__mux2_1 _16964_ (.A0(\rvcpu.dp.rf.reg_file_arr[1][19] ),
    .A1(_14447_),
    .S(_04731_),
    .X(_04734_));
 sky130_fd_sc_hd__clkbuf_1 _16965_ (.A(_04734_),
    .X(_01559_));
 sky130_fd_sc_hd__mux2_1 _16966_ (.A0(\rvcpu.dp.rf.reg_file_arr[1][18] ),
    .A1(_14449_),
    .S(_04731_),
    .X(_04735_));
 sky130_fd_sc_hd__clkbuf_1 _16967_ (.A(_04735_),
    .X(_01558_));
 sky130_fd_sc_hd__mux2_1 _16968_ (.A0(\rvcpu.dp.rf.reg_file_arr[1][17] ),
    .A1(_14451_),
    .S(_04731_),
    .X(_04736_));
 sky130_fd_sc_hd__clkbuf_1 _16969_ (.A(_04736_),
    .X(_01557_));
 sky130_fd_sc_hd__mux2_1 _16970_ (.A0(\rvcpu.dp.rf.reg_file_arr[1][16] ),
    .A1(_14453_),
    .S(_04731_),
    .X(_04737_));
 sky130_fd_sc_hd__clkbuf_1 _16971_ (.A(_04737_),
    .X(_01556_));
 sky130_fd_sc_hd__mux2_1 _16972_ (.A0(\rvcpu.dp.rf.reg_file_arr[1][15] ),
    .A1(_14455_),
    .S(_04731_),
    .X(_04738_));
 sky130_fd_sc_hd__clkbuf_1 _16973_ (.A(_04738_),
    .X(_01555_));
 sky130_fd_sc_hd__mux2_1 _16974_ (.A0(\rvcpu.dp.rf.reg_file_arr[1][14] ),
    .A1(_14457_),
    .S(_04731_),
    .X(_04739_));
 sky130_fd_sc_hd__clkbuf_1 _16975_ (.A(_04739_),
    .X(_01554_));
 sky130_fd_sc_hd__mux2_1 _16976_ (.A0(\rvcpu.dp.rf.reg_file_arr[1][13] ),
    .A1(_14459_),
    .S(_04731_),
    .X(_04740_));
 sky130_fd_sc_hd__clkbuf_1 _16977_ (.A(_04740_),
    .X(_01553_));
 sky130_fd_sc_hd__mux2_1 _16978_ (.A0(\rvcpu.dp.rf.reg_file_arr[1][12] ),
    .A1(_14461_),
    .S(_04731_),
    .X(_04741_));
 sky130_fd_sc_hd__clkbuf_1 _16979_ (.A(_04741_),
    .X(_01552_));
 sky130_fd_sc_hd__buf_4 _16980_ (.A(_04719_),
    .X(_04742_));
 sky130_fd_sc_hd__mux2_1 _16981_ (.A0(\rvcpu.dp.rf.reg_file_arr[1][11] ),
    .A1(_14463_),
    .S(_04742_),
    .X(_04743_));
 sky130_fd_sc_hd__clkbuf_1 _16982_ (.A(_04743_),
    .X(_01551_));
 sky130_fd_sc_hd__mux2_1 _16983_ (.A0(\rvcpu.dp.rf.reg_file_arr[1][10] ),
    .A1(_14466_),
    .S(_04742_),
    .X(_04744_));
 sky130_fd_sc_hd__clkbuf_1 _16984_ (.A(_04744_),
    .X(_01550_));
 sky130_fd_sc_hd__mux2_1 _16985_ (.A0(\rvcpu.dp.rf.reg_file_arr[1][9] ),
    .A1(_14468_),
    .S(_04742_),
    .X(_04745_));
 sky130_fd_sc_hd__clkbuf_1 _16986_ (.A(_04745_),
    .X(_01549_));
 sky130_fd_sc_hd__mux2_1 _16987_ (.A0(\rvcpu.dp.rf.reg_file_arr[1][8] ),
    .A1(_14470_),
    .S(_04742_),
    .X(_04746_));
 sky130_fd_sc_hd__clkbuf_1 _16988_ (.A(_04746_),
    .X(_01548_));
 sky130_fd_sc_hd__mux2_1 _16989_ (.A0(\rvcpu.dp.rf.reg_file_arr[1][7] ),
    .A1(_14472_),
    .S(_04742_),
    .X(_04747_));
 sky130_fd_sc_hd__clkbuf_1 _16990_ (.A(_04747_),
    .X(_01547_));
 sky130_fd_sc_hd__mux2_1 _16991_ (.A0(\rvcpu.dp.rf.reg_file_arr[1][6] ),
    .A1(_14474_),
    .S(_04742_),
    .X(_04748_));
 sky130_fd_sc_hd__clkbuf_1 _16992_ (.A(_04748_),
    .X(_01546_));
 sky130_fd_sc_hd__mux2_1 _16993_ (.A0(\rvcpu.dp.rf.reg_file_arr[1][5] ),
    .A1(_14476_),
    .S(_04742_),
    .X(_04749_));
 sky130_fd_sc_hd__clkbuf_1 _16994_ (.A(_04749_),
    .X(_01545_));
 sky130_fd_sc_hd__mux2_1 _16995_ (.A0(\rvcpu.dp.rf.reg_file_arr[1][4] ),
    .A1(_14478_),
    .S(_04742_),
    .X(_04750_));
 sky130_fd_sc_hd__clkbuf_1 _16996_ (.A(_04750_),
    .X(_01544_));
 sky130_fd_sc_hd__mux2_1 _16997_ (.A0(\rvcpu.dp.rf.reg_file_arr[1][3] ),
    .A1(_14480_),
    .S(_04742_),
    .X(_04751_));
 sky130_fd_sc_hd__clkbuf_1 _16998_ (.A(_04751_),
    .X(_01543_));
 sky130_fd_sc_hd__mux2_1 _16999_ (.A0(\rvcpu.dp.rf.reg_file_arr[1][2] ),
    .A1(_14482_),
    .S(_04742_),
    .X(_04752_));
 sky130_fd_sc_hd__clkbuf_1 _17000_ (.A(_04752_),
    .X(_01542_));
 sky130_fd_sc_hd__mux2_1 _17001_ (.A0(\rvcpu.dp.rf.reg_file_arr[1][1] ),
    .A1(_14484_),
    .S(_04719_),
    .X(_04753_));
 sky130_fd_sc_hd__clkbuf_1 _17002_ (.A(_04753_),
    .X(_01541_));
 sky130_fd_sc_hd__mux2_1 _17003_ (.A0(\rvcpu.dp.rf.reg_file_arr[1][0] ),
    .A1(_14486_),
    .S(_04719_),
    .X(_04754_));
 sky130_fd_sc_hd__clkbuf_1 _17004_ (.A(_04754_),
    .X(_01540_));
 sky130_fd_sc_hd__and3_2 _17005_ (.A(_13174_),
    .B(_13175_),
    .C(_13176_),
    .X(_04755_));
 sky130_fd_sc_hd__and2_2 _17006_ (.A(_04464_),
    .B(_04755_),
    .X(_04756_));
 sky130_fd_sc_hd__buf_4 _17007_ (.A(_04756_),
    .X(_04757_));
 sky130_fd_sc_hd__mux2_1 _17008_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][31] ),
    .A1(_14420_),
    .S(_04757_),
    .X(_04758_));
 sky130_fd_sc_hd__clkbuf_1 _17009_ (.A(_04758_),
    .X(_01531_));
 sky130_fd_sc_hd__mux2_1 _17010_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][30] ),
    .A1(_14424_),
    .S(_04757_),
    .X(_04759_));
 sky130_fd_sc_hd__clkbuf_1 _17011_ (.A(_04759_),
    .X(_01530_));
 sky130_fd_sc_hd__mux2_1 _17012_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][29] ),
    .A1(_14426_),
    .S(_04757_),
    .X(_04760_));
 sky130_fd_sc_hd__clkbuf_1 _17013_ (.A(_04760_),
    .X(_01529_));
 sky130_fd_sc_hd__mux2_1 _17014_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][28] ),
    .A1(_14428_),
    .S(_04757_),
    .X(_04761_));
 sky130_fd_sc_hd__clkbuf_1 _17015_ (.A(_04761_),
    .X(_01528_));
 sky130_fd_sc_hd__mux2_1 _17016_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][27] ),
    .A1(_14430_),
    .S(_04757_),
    .X(_04762_));
 sky130_fd_sc_hd__clkbuf_1 _17017_ (.A(_04762_),
    .X(_01527_));
 sky130_fd_sc_hd__mux2_1 _17018_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][26] ),
    .A1(_14432_),
    .S(_04757_),
    .X(_04763_));
 sky130_fd_sc_hd__clkbuf_1 _17019_ (.A(_04763_),
    .X(_01526_));
 sky130_fd_sc_hd__mux2_1 _17020_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][25] ),
    .A1(_14434_),
    .S(_04757_),
    .X(_04764_));
 sky130_fd_sc_hd__clkbuf_1 _17021_ (.A(_04764_),
    .X(_01525_));
 sky130_fd_sc_hd__mux2_1 _17022_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][24] ),
    .A1(_14436_),
    .S(_04757_),
    .X(_04765_));
 sky130_fd_sc_hd__clkbuf_1 _17023_ (.A(_04765_),
    .X(_01524_));
 sky130_fd_sc_hd__mux2_1 _17024_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][23] ),
    .A1(_14438_),
    .S(_04757_),
    .X(_04766_));
 sky130_fd_sc_hd__clkbuf_1 _17025_ (.A(_04766_),
    .X(_01523_));
 sky130_fd_sc_hd__mux2_1 _17026_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][22] ),
    .A1(_14440_),
    .S(_04757_),
    .X(_04767_));
 sky130_fd_sc_hd__clkbuf_1 _17027_ (.A(_04767_),
    .X(_01522_));
 sky130_fd_sc_hd__buf_4 _17028_ (.A(_04756_),
    .X(_04768_));
 sky130_fd_sc_hd__mux2_1 _17029_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][21] ),
    .A1(_14442_),
    .S(_04768_),
    .X(_04769_));
 sky130_fd_sc_hd__clkbuf_1 _17030_ (.A(_04769_),
    .X(_01521_));
 sky130_fd_sc_hd__mux2_1 _17031_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][20] ),
    .A1(_14445_),
    .S(_04768_),
    .X(_04770_));
 sky130_fd_sc_hd__clkbuf_1 _17032_ (.A(_04770_),
    .X(_01520_));
 sky130_fd_sc_hd__mux2_1 _17033_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][19] ),
    .A1(_14447_),
    .S(_04768_),
    .X(_04771_));
 sky130_fd_sc_hd__clkbuf_1 _17034_ (.A(_04771_),
    .X(_01519_));
 sky130_fd_sc_hd__mux2_1 _17035_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][18] ),
    .A1(_14449_),
    .S(_04768_),
    .X(_04772_));
 sky130_fd_sc_hd__clkbuf_1 _17036_ (.A(_04772_),
    .X(_01518_));
 sky130_fd_sc_hd__mux2_1 _17037_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][17] ),
    .A1(_14451_),
    .S(_04768_),
    .X(_04773_));
 sky130_fd_sc_hd__clkbuf_1 _17038_ (.A(_04773_),
    .X(_01517_));
 sky130_fd_sc_hd__mux2_1 _17039_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][16] ),
    .A1(_14453_),
    .S(_04768_),
    .X(_04774_));
 sky130_fd_sc_hd__clkbuf_1 _17040_ (.A(_04774_),
    .X(_01516_));
 sky130_fd_sc_hd__mux2_1 _17041_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][15] ),
    .A1(_14455_),
    .S(_04768_),
    .X(_04775_));
 sky130_fd_sc_hd__clkbuf_1 _17042_ (.A(_04775_),
    .X(_01515_));
 sky130_fd_sc_hd__mux2_1 _17043_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][14] ),
    .A1(_14457_),
    .S(_04768_),
    .X(_04776_));
 sky130_fd_sc_hd__clkbuf_1 _17044_ (.A(_04776_),
    .X(_01514_));
 sky130_fd_sc_hd__mux2_1 _17045_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][13] ),
    .A1(_14459_),
    .S(_04768_),
    .X(_04777_));
 sky130_fd_sc_hd__clkbuf_1 _17046_ (.A(_04777_),
    .X(_01513_));
 sky130_fd_sc_hd__mux2_1 _17047_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][12] ),
    .A1(_14461_),
    .S(_04768_),
    .X(_04778_));
 sky130_fd_sc_hd__clkbuf_1 _17048_ (.A(_04778_),
    .X(_01512_));
 sky130_fd_sc_hd__buf_4 _17049_ (.A(_04756_),
    .X(_04779_));
 sky130_fd_sc_hd__mux2_1 _17050_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][11] ),
    .A1(_14463_),
    .S(_04779_),
    .X(_04780_));
 sky130_fd_sc_hd__clkbuf_1 _17051_ (.A(_04780_),
    .X(_01511_));
 sky130_fd_sc_hd__mux2_1 _17052_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][10] ),
    .A1(_14466_),
    .S(_04779_),
    .X(_04781_));
 sky130_fd_sc_hd__clkbuf_1 _17053_ (.A(_04781_),
    .X(_01510_));
 sky130_fd_sc_hd__mux2_1 _17054_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][9] ),
    .A1(_14468_),
    .S(_04779_),
    .X(_04782_));
 sky130_fd_sc_hd__clkbuf_1 _17055_ (.A(_04782_),
    .X(_01509_));
 sky130_fd_sc_hd__mux2_1 _17056_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][8] ),
    .A1(_14470_),
    .S(_04779_),
    .X(_04783_));
 sky130_fd_sc_hd__clkbuf_1 _17057_ (.A(_04783_),
    .X(_01508_));
 sky130_fd_sc_hd__mux2_1 _17058_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][7] ),
    .A1(_14472_),
    .S(_04779_),
    .X(_04784_));
 sky130_fd_sc_hd__clkbuf_1 _17059_ (.A(_04784_),
    .X(_01507_));
 sky130_fd_sc_hd__mux2_1 _17060_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][6] ),
    .A1(_14474_),
    .S(_04779_),
    .X(_04785_));
 sky130_fd_sc_hd__clkbuf_1 _17061_ (.A(_04785_),
    .X(_01506_));
 sky130_fd_sc_hd__mux2_1 _17062_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][5] ),
    .A1(_14476_),
    .S(_04779_),
    .X(_04786_));
 sky130_fd_sc_hd__clkbuf_1 _17063_ (.A(_04786_),
    .X(_01505_));
 sky130_fd_sc_hd__mux2_1 _17064_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][4] ),
    .A1(_14478_),
    .S(_04779_),
    .X(_04787_));
 sky130_fd_sc_hd__clkbuf_1 _17065_ (.A(_04787_),
    .X(_01504_));
 sky130_fd_sc_hd__mux2_1 _17066_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][3] ),
    .A1(_14480_),
    .S(_04779_),
    .X(_04788_));
 sky130_fd_sc_hd__clkbuf_1 _17067_ (.A(_04788_),
    .X(_01503_));
 sky130_fd_sc_hd__mux2_1 _17068_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][2] ),
    .A1(_14482_),
    .S(_04779_),
    .X(_04789_));
 sky130_fd_sc_hd__clkbuf_1 _17069_ (.A(_04789_),
    .X(_01502_));
 sky130_fd_sc_hd__mux2_1 _17070_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][1] ),
    .A1(_14484_),
    .S(_04756_),
    .X(_04790_));
 sky130_fd_sc_hd__clkbuf_1 _17071_ (.A(_04790_),
    .X(_01501_));
 sky130_fd_sc_hd__mux2_1 _17072_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][0] ),
    .A1(_14486_),
    .S(_04756_),
    .X(_04791_));
 sky130_fd_sc_hd__clkbuf_1 _17073_ (.A(_04791_),
    .X(_01500_));
 sky130_fd_sc_hd__nand2_4 _17074_ (.A(_14128_),
    .B(_04755_),
    .Y(_04792_));
 sky130_fd_sc_hd__clkbuf_4 _17075_ (.A(_04792_),
    .X(_04793_));
 sky130_fd_sc_hd__mux2_1 _17076_ (.A0(_14127_),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][31] ),
    .S(_04793_),
    .X(_04794_));
 sky130_fd_sc_hd__clkbuf_1 _17077_ (.A(_04794_),
    .X(_01499_));
 sky130_fd_sc_hd__mux2_1 _17078_ (.A0(_14133_),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][30] ),
    .S(_04793_),
    .X(_04795_));
 sky130_fd_sc_hd__clkbuf_1 _17079_ (.A(_04795_),
    .X(_01498_));
 sky130_fd_sc_hd__mux2_1 _17080_ (.A0(_14135_),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][29] ),
    .S(_04793_),
    .X(_04796_));
 sky130_fd_sc_hd__clkbuf_1 _17081_ (.A(_04796_),
    .X(_01497_));
 sky130_fd_sc_hd__mux2_1 _17082_ (.A0(_14137_),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][28] ),
    .S(_04793_),
    .X(_04797_));
 sky130_fd_sc_hd__clkbuf_1 _17083_ (.A(_04797_),
    .X(_01496_));
 sky130_fd_sc_hd__mux2_1 _17084_ (.A0(_14139_),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][27] ),
    .S(_04793_),
    .X(_04798_));
 sky130_fd_sc_hd__clkbuf_1 _17085_ (.A(_04798_),
    .X(_01495_));
 sky130_fd_sc_hd__mux2_1 _17086_ (.A0(_14141_),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][26] ),
    .S(_04793_),
    .X(_04799_));
 sky130_fd_sc_hd__clkbuf_1 _17087_ (.A(_04799_),
    .X(_01494_));
 sky130_fd_sc_hd__mux2_1 _17088_ (.A0(_14143_),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][25] ),
    .S(_04793_),
    .X(_04800_));
 sky130_fd_sc_hd__clkbuf_1 _17089_ (.A(_04800_),
    .X(_01493_));
 sky130_fd_sc_hd__mux2_1 _17090_ (.A0(_14145_),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][24] ),
    .S(_04793_),
    .X(_04801_));
 sky130_fd_sc_hd__clkbuf_1 _17091_ (.A(_04801_),
    .X(_01492_));
 sky130_fd_sc_hd__mux2_1 _17092_ (.A0(_14147_),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][23] ),
    .S(_04793_),
    .X(_04802_));
 sky130_fd_sc_hd__clkbuf_1 _17093_ (.A(_04802_),
    .X(_01491_));
 sky130_fd_sc_hd__mux2_1 _17094_ (.A0(_14149_),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][22] ),
    .S(_04793_),
    .X(_04803_));
 sky130_fd_sc_hd__clkbuf_1 _17095_ (.A(_04803_),
    .X(_01490_));
 sky130_fd_sc_hd__clkbuf_4 _17096_ (.A(_04792_),
    .X(_04804_));
 sky130_fd_sc_hd__mux2_1 _17097_ (.A0(_14151_),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][21] ),
    .S(_04804_),
    .X(_04805_));
 sky130_fd_sc_hd__clkbuf_1 _17098_ (.A(_04805_),
    .X(_01489_));
 sky130_fd_sc_hd__mux2_1 _17099_ (.A0(_14154_),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][20] ),
    .S(_04804_),
    .X(_04806_));
 sky130_fd_sc_hd__clkbuf_1 _17100_ (.A(_04806_),
    .X(_01488_));
 sky130_fd_sc_hd__mux2_1 _17101_ (.A0(_14156_),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][19] ),
    .S(_04804_),
    .X(_04807_));
 sky130_fd_sc_hd__clkbuf_1 _17102_ (.A(_04807_),
    .X(_01487_));
 sky130_fd_sc_hd__mux2_1 _17103_ (.A0(_14158_),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][18] ),
    .S(_04804_),
    .X(_04808_));
 sky130_fd_sc_hd__clkbuf_1 _17104_ (.A(_04808_),
    .X(_01486_));
 sky130_fd_sc_hd__mux2_1 _17105_ (.A0(_14160_),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][17] ),
    .S(_04804_),
    .X(_04809_));
 sky130_fd_sc_hd__clkbuf_1 _17106_ (.A(_04809_),
    .X(_01485_));
 sky130_fd_sc_hd__mux2_1 _17107_ (.A0(_14162_),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][16] ),
    .S(_04804_),
    .X(_04810_));
 sky130_fd_sc_hd__clkbuf_1 _17108_ (.A(_04810_),
    .X(_01484_));
 sky130_fd_sc_hd__mux2_1 _17109_ (.A0(_14164_),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][15] ),
    .S(_04804_),
    .X(_04811_));
 sky130_fd_sc_hd__clkbuf_1 _17110_ (.A(_04811_),
    .X(_01483_));
 sky130_fd_sc_hd__mux2_1 _17111_ (.A0(_14166_),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][14] ),
    .S(_04804_),
    .X(_04812_));
 sky130_fd_sc_hd__clkbuf_1 _17112_ (.A(_04812_),
    .X(_01482_));
 sky130_fd_sc_hd__mux2_1 _17113_ (.A0(_14168_),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][13] ),
    .S(_04804_),
    .X(_04813_));
 sky130_fd_sc_hd__clkbuf_1 _17114_ (.A(_04813_),
    .X(_01481_));
 sky130_fd_sc_hd__mux2_1 _17115_ (.A0(_14170_),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][12] ),
    .S(_04804_),
    .X(_04814_));
 sky130_fd_sc_hd__clkbuf_1 _17116_ (.A(_04814_),
    .X(_01480_));
 sky130_fd_sc_hd__clkbuf_4 _17117_ (.A(_04792_),
    .X(_04815_));
 sky130_fd_sc_hd__mux2_1 _17118_ (.A0(_14172_),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][11] ),
    .S(_04815_),
    .X(_04816_));
 sky130_fd_sc_hd__clkbuf_1 _17119_ (.A(_04816_),
    .X(_01479_));
 sky130_fd_sc_hd__mux2_1 _17120_ (.A0(_14175_),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][10] ),
    .S(_04815_),
    .X(_04817_));
 sky130_fd_sc_hd__clkbuf_1 _17121_ (.A(_04817_),
    .X(_01478_));
 sky130_fd_sc_hd__mux2_1 _17122_ (.A0(_14177_),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][9] ),
    .S(_04815_),
    .X(_04818_));
 sky130_fd_sc_hd__clkbuf_1 _17123_ (.A(_04818_),
    .X(_01477_));
 sky130_fd_sc_hd__mux2_1 _17124_ (.A0(_14179_),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][8] ),
    .S(_04815_),
    .X(_04819_));
 sky130_fd_sc_hd__clkbuf_1 _17125_ (.A(_04819_),
    .X(_01476_));
 sky130_fd_sc_hd__mux2_1 _17126_ (.A0(_14181_),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][7] ),
    .S(_04815_),
    .X(_04820_));
 sky130_fd_sc_hd__clkbuf_1 _17127_ (.A(_04820_),
    .X(_01475_));
 sky130_fd_sc_hd__mux2_1 _17128_ (.A0(_14183_),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][6] ),
    .S(_04815_),
    .X(_04821_));
 sky130_fd_sc_hd__clkbuf_1 _17129_ (.A(_04821_),
    .X(_01474_));
 sky130_fd_sc_hd__mux2_1 _17130_ (.A0(_14185_),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][5] ),
    .S(_04815_),
    .X(_04822_));
 sky130_fd_sc_hd__clkbuf_1 _17131_ (.A(_04822_),
    .X(_01473_));
 sky130_fd_sc_hd__mux2_1 _17132_ (.A0(_14187_),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][4] ),
    .S(_04815_),
    .X(_04823_));
 sky130_fd_sc_hd__clkbuf_1 _17133_ (.A(_04823_),
    .X(_01472_));
 sky130_fd_sc_hd__mux2_1 _17134_ (.A0(_14189_),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][3] ),
    .S(_04815_),
    .X(_04824_));
 sky130_fd_sc_hd__clkbuf_1 _17135_ (.A(_04824_),
    .X(_01471_));
 sky130_fd_sc_hd__mux2_1 _17136_ (.A0(_14191_),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][2] ),
    .S(_04815_),
    .X(_04825_));
 sky130_fd_sc_hd__clkbuf_1 _17137_ (.A(_04825_),
    .X(_01470_));
 sky130_fd_sc_hd__mux2_1 _17138_ (.A0(_14193_),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][1] ),
    .S(_04792_),
    .X(_04826_));
 sky130_fd_sc_hd__clkbuf_1 _17139_ (.A(_04826_),
    .X(_01469_));
 sky130_fd_sc_hd__mux2_1 _17140_ (.A0(_14195_),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][0] ),
    .S(_04792_),
    .X(_04827_));
 sky130_fd_sc_hd__clkbuf_1 _17141_ (.A(_04827_),
    .X(_01468_));
 sky130_fd_sc_hd__nand2_2 _17142_ (.A(_04538_),
    .B(_04755_),
    .Y(_04828_));
 sky130_fd_sc_hd__buf_4 _17143_ (.A(_04828_),
    .X(_04829_));
 sky130_fd_sc_hd__mux2_1 _17144_ (.A0(_14127_),
    .A1(\rvcpu.dp.rf.reg_file_arr[22][31] ),
    .S(_04829_),
    .X(_04830_));
 sky130_fd_sc_hd__clkbuf_1 _17145_ (.A(_04830_),
    .X(_01467_));
 sky130_fd_sc_hd__mux2_1 _17146_ (.A0(_14133_),
    .A1(\rvcpu.dp.rf.reg_file_arr[22][30] ),
    .S(_04829_),
    .X(_04831_));
 sky130_fd_sc_hd__clkbuf_1 _17147_ (.A(_04831_),
    .X(_01466_));
 sky130_fd_sc_hd__mux2_1 _17148_ (.A0(_14135_),
    .A1(\rvcpu.dp.rf.reg_file_arr[22][29] ),
    .S(_04829_),
    .X(_04832_));
 sky130_fd_sc_hd__clkbuf_1 _17149_ (.A(_04832_),
    .X(_01465_));
 sky130_fd_sc_hd__mux2_1 _17150_ (.A0(_14137_),
    .A1(\rvcpu.dp.rf.reg_file_arr[22][28] ),
    .S(_04829_),
    .X(_04833_));
 sky130_fd_sc_hd__clkbuf_1 _17151_ (.A(_04833_),
    .X(_01464_));
 sky130_fd_sc_hd__mux2_1 _17152_ (.A0(_14139_),
    .A1(\rvcpu.dp.rf.reg_file_arr[22][27] ),
    .S(_04829_),
    .X(_04834_));
 sky130_fd_sc_hd__clkbuf_1 _17153_ (.A(_04834_),
    .X(_01463_));
 sky130_fd_sc_hd__mux2_1 _17154_ (.A0(_14141_),
    .A1(\rvcpu.dp.rf.reg_file_arr[22][26] ),
    .S(_04829_),
    .X(_04835_));
 sky130_fd_sc_hd__clkbuf_1 _17155_ (.A(_04835_),
    .X(_01462_));
 sky130_fd_sc_hd__mux2_1 _17156_ (.A0(_14143_),
    .A1(\rvcpu.dp.rf.reg_file_arr[22][25] ),
    .S(_04829_),
    .X(_04836_));
 sky130_fd_sc_hd__clkbuf_1 _17157_ (.A(_04836_),
    .X(_01461_));
 sky130_fd_sc_hd__mux2_1 _17158_ (.A0(_14145_),
    .A1(\rvcpu.dp.rf.reg_file_arr[22][24] ),
    .S(_04829_),
    .X(_04837_));
 sky130_fd_sc_hd__clkbuf_1 _17159_ (.A(_04837_),
    .X(_01460_));
 sky130_fd_sc_hd__mux2_1 _17160_ (.A0(_14147_),
    .A1(\rvcpu.dp.rf.reg_file_arr[22][23] ),
    .S(_04829_),
    .X(_04838_));
 sky130_fd_sc_hd__clkbuf_1 _17161_ (.A(_04838_),
    .X(_01459_));
 sky130_fd_sc_hd__mux2_1 _17162_ (.A0(_14149_),
    .A1(\rvcpu.dp.rf.reg_file_arr[22][22] ),
    .S(_04829_),
    .X(_04839_));
 sky130_fd_sc_hd__clkbuf_1 _17163_ (.A(_04839_),
    .X(_01458_));
 sky130_fd_sc_hd__buf_4 _17164_ (.A(_04828_),
    .X(_04840_));
 sky130_fd_sc_hd__mux2_1 _17165_ (.A0(_14151_),
    .A1(\rvcpu.dp.rf.reg_file_arr[22][21] ),
    .S(_04840_),
    .X(_04841_));
 sky130_fd_sc_hd__clkbuf_1 _17166_ (.A(_04841_),
    .X(_01457_));
 sky130_fd_sc_hd__mux2_1 _17167_ (.A0(_14154_),
    .A1(\rvcpu.dp.rf.reg_file_arr[22][20] ),
    .S(_04840_),
    .X(_04842_));
 sky130_fd_sc_hd__clkbuf_1 _17168_ (.A(_04842_),
    .X(_01456_));
 sky130_fd_sc_hd__mux2_1 _17169_ (.A0(_14156_),
    .A1(\rvcpu.dp.rf.reg_file_arr[22][19] ),
    .S(_04840_),
    .X(_04843_));
 sky130_fd_sc_hd__clkbuf_1 _17170_ (.A(_04843_),
    .X(_01455_));
 sky130_fd_sc_hd__mux2_1 _17171_ (.A0(_14158_),
    .A1(\rvcpu.dp.rf.reg_file_arr[22][18] ),
    .S(_04840_),
    .X(_04844_));
 sky130_fd_sc_hd__clkbuf_1 _17172_ (.A(_04844_),
    .X(_01454_));
 sky130_fd_sc_hd__mux2_1 _17173_ (.A0(_14160_),
    .A1(\rvcpu.dp.rf.reg_file_arr[22][17] ),
    .S(_04840_),
    .X(_04845_));
 sky130_fd_sc_hd__clkbuf_1 _17174_ (.A(_04845_),
    .X(_01453_));
 sky130_fd_sc_hd__mux2_1 _17175_ (.A0(_14162_),
    .A1(\rvcpu.dp.rf.reg_file_arr[22][16] ),
    .S(_04840_),
    .X(_04846_));
 sky130_fd_sc_hd__clkbuf_1 _17176_ (.A(_04846_),
    .X(_01452_));
 sky130_fd_sc_hd__mux2_1 _17177_ (.A0(_14164_),
    .A1(\rvcpu.dp.rf.reg_file_arr[22][15] ),
    .S(_04840_),
    .X(_04847_));
 sky130_fd_sc_hd__clkbuf_1 _17178_ (.A(_04847_),
    .X(_01451_));
 sky130_fd_sc_hd__mux2_1 _17179_ (.A0(_14166_),
    .A1(\rvcpu.dp.rf.reg_file_arr[22][14] ),
    .S(_04840_),
    .X(_04848_));
 sky130_fd_sc_hd__clkbuf_1 _17180_ (.A(_04848_),
    .X(_01450_));
 sky130_fd_sc_hd__mux2_1 _17181_ (.A0(_14168_),
    .A1(\rvcpu.dp.rf.reg_file_arr[22][13] ),
    .S(_04840_),
    .X(_04849_));
 sky130_fd_sc_hd__clkbuf_1 _17182_ (.A(_04849_),
    .X(_01449_));
 sky130_fd_sc_hd__mux2_1 _17183_ (.A0(_14170_),
    .A1(\rvcpu.dp.rf.reg_file_arr[22][12] ),
    .S(_04840_),
    .X(_04850_));
 sky130_fd_sc_hd__clkbuf_1 _17184_ (.A(_04850_),
    .X(_01448_));
 sky130_fd_sc_hd__clkbuf_4 _17185_ (.A(_04828_),
    .X(_04851_));
 sky130_fd_sc_hd__mux2_1 _17186_ (.A0(_14172_),
    .A1(\rvcpu.dp.rf.reg_file_arr[22][11] ),
    .S(_04851_),
    .X(_04852_));
 sky130_fd_sc_hd__clkbuf_1 _17187_ (.A(_04852_),
    .X(_01447_));
 sky130_fd_sc_hd__mux2_1 _17188_ (.A0(_14175_),
    .A1(\rvcpu.dp.rf.reg_file_arr[22][10] ),
    .S(_04851_),
    .X(_04853_));
 sky130_fd_sc_hd__clkbuf_1 _17189_ (.A(_04853_),
    .X(_01446_));
 sky130_fd_sc_hd__mux2_1 _17190_ (.A0(_14177_),
    .A1(\rvcpu.dp.rf.reg_file_arr[22][9] ),
    .S(_04851_),
    .X(_04854_));
 sky130_fd_sc_hd__clkbuf_1 _17191_ (.A(_04854_),
    .X(_01445_));
 sky130_fd_sc_hd__mux2_1 _17192_ (.A0(_14179_),
    .A1(\rvcpu.dp.rf.reg_file_arr[22][8] ),
    .S(_04851_),
    .X(_04855_));
 sky130_fd_sc_hd__clkbuf_1 _17193_ (.A(_04855_),
    .X(_01444_));
 sky130_fd_sc_hd__mux2_1 _17194_ (.A0(_14181_),
    .A1(\rvcpu.dp.rf.reg_file_arr[22][7] ),
    .S(_04851_),
    .X(_04856_));
 sky130_fd_sc_hd__clkbuf_1 _17195_ (.A(_04856_),
    .X(_01443_));
 sky130_fd_sc_hd__mux2_1 _17196_ (.A0(_14183_),
    .A1(\rvcpu.dp.rf.reg_file_arr[22][6] ),
    .S(_04851_),
    .X(_04857_));
 sky130_fd_sc_hd__clkbuf_1 _17197_ (.A(_04857_),
    .X(_01442_));
 sky130_fd_sc_hd__mux2_1 _17198_ (.A0(_14185_),
    .A1(\rvcpu.dp.rf.reg_file_arr[22][5] ),
    .S(_04851_),
    .X(_04858_));
 sky130_fd_sc_hd__clkbuf_1 _17199_ (.A(_04858_),
    .X(_01441_));
 sky130_fd_sc_hd__mux2_1 _17200_ (.A0(_14187_),
    .A1(\rvcpu.dp.rf.reg_file_arr[22][4] ),
    .S(_04851_),
    .X(_04859_));
 sky130_fd_sc_hd__clkbuf_1 _17201_ (.A(_04859_),
    .X(_01440_));
 sky130_fd_sc_hd__mux2_1 _17202_ (.A0(_14189_),
    .A1(\rvcpu.dp.rf.reg_file_arr[22][3] ),
    .S(_04851_),
    .X(_04860_));
 sky130_fd_sc_hd__clkbuf_1 _17203_ (.A(_04860_),
    .X(_01439_));
 sky130_fd_sc_hd__mux2_1 _17204_ (.A0(_14191_),
    .A1(\rvcpu.dp.rf.reg_file_arr[22][2] ),
    .S(_04851_),
    .X(_04861_));
 sky130_fd_sc_hd__clkbuf_1 _17205_ (.A(_04861_),
    .X(_01438_));
 sky130_fd_sc_hd__mux2_1 _17206_ (.A0(_14193_),
    .A1(\rvcpu.dp.rf.reg_file_arr[22][1] ),
    .S(_04828_),
    .X(_04862_));
 sky130_fd_sc_hd__clkbuf_1 _17207_ (.A(_04862_),
    .X(_01437_));
 sky130_fd_sc_hd__mux2_1 _17208_ (.A0(_14195_),
    .A1(\rvcpu.dp.rf.reg_file_arr[22][0] ),
    .S(_04828_),
    .X(_04863_));
 sky130_fd_sc_hd__clkbuf_1 _17209_ (.A(_04863_),
    .X(_01436_));
 sky130_fd_sc_hd__nand2_2 _17210_ (.A(_14197_),
    .B(_04755_),
    .Y(_04864_));
 sky130_fd_sc_hd__buf_4 _17211_ (.A(_04864_),
    .X(_04865_));
 sky130_fd_sc_hd__mux2_1 _17212_ (.A0(_14127_),
    .A1(\rvcpu.dp.rf.reg_file_arr[23][31] ),
    .S(_04865_),
    .X(_04866_));
 sky130_fd_sc_hd__clkbuf_1 _17213_ (.A(_04866_),
    .X(_01435_));
 sky130_fd_sc_hd__mux2_1 _17214_ (.A0(_14133_),
    .A1(\rvcpu.dp.rf.reg_file_arr[23][30] ),
    .S(_04865_),
    .X(_04867_));
 sky130_fd_sc_hd__clkbuf_1 _17215_ (.A(_04867_),
    .X(_01434_));
 sky130_fd_sc_hd__mux2_1 _17216_ (.A0(_14135_),
    .A1(\rvcpu.dp.rf.reg_file_arr[23][29] ),
    .S(_04865_),
    .X(_04868_));
 sky130_fd_sc_hd__clkbuf_1 _17217_ (.A(_04868_),
    .X(_01433_));
 sky130_fd_sc_hd__mux2_1 _17218_ (.A0(_14137_),
    .A1(\rvcpu.dp.rf.reg_file_arr[23][28] ),
    .S(_04865_),
    .X(_04869_));
 sky130_fd_sc_hd__clkbuf_1 _17219_ (.A(_04869_),
    .X(_01432_));
 sky130_fd_sc_hd__mux2_1 _17220_ (.A0(_14139_),
    .A1(\rvcpu.dp.rf.reg_file_arr[23][27] ),
    .S(_04865_),
    .X(_04870_));
 sky130_fd_sc_hd__clkbuf_1 _17221_ (.A(_04870_),
    .X(_01431_));
 sky130_fd_sc_hd__mux2_1 _17222_ (.A0(_14141_),
    .A1(\rvcpu.dp.rf.reg_file_arr[23][26] ),
    .S(_04865_),
    .X(_04871_));
 sky130_fd_sc_hd__clkbuf_1 _17223_ (.A(_04871_),
    .X(_01430_));
 sky130_fd_sc_hd__mux2_1 _17224_ (.A0(_14143_),
    .A1(\rvcpu.dp.rf.reg_file_arr[23][25] ),
    .S(_04865_),
    .X(_04872_));
 sky130_fd_sc_hd__clkbuf_1 _17225_ (.A(_04872_),
    .X(_01429_));
 sky130_fd_sc_hd__mux2_1 _17226_ (.A0(_14145_),
    .A1(\rvcpu.dp.rf.reg_file_arr[23][24] ),
    .S(_04865_),
    .X(_04873_));
 sky130_fd_sc_hd__clkbuf_1 _17227_ (.A(_04873_),
    .X(_01428_));
 sky130_fd_sc_hd__mux2_1 _17228_ (.A0(_14147_),
    .A1(\rvcpu.dp.rf.reg_file_arr[23][23] ),
    .S(_04865_),
    .X(_04874_));
 sky130_fd_sc_hd__clkbuf_1 _17229_ (.A(_04874_),
    .X(_01427_));
 sky130_fd_sc_hd__mux2_1 _17230_ (.A0(_14149_),
    .A1(\rvcpu.dp.rf.reg_file_arr[23][22] ),
    .S(_04865_),
    .X(_04875_));
 sky130_fd_sc_hd__clkbuf_1 _17231_ (.A(_04875_),
    .X(_01426_));
 sky130_fd_sc_hd__buf_4 _17232_ (.A(_04864_),
    .X(_04876_));
 sky130_fd_sc_hd__mux2_1 _17233_ (.A0(_14151_),
    .A1(\rvcpu.dp.rf.reg_file_arr[23][21] ),
    .S(_04876_),
    .X(_04877_));
 sky130_fd_sc_hd__clkbuf_1 _17234_ (.A(_04877_),
    .X(_01425_));
 sky130_fd_sc_hd__mux2_1 _17235_ (.A0(_14154_),
    .A1(\rvcpu.dp.rf.reg_file_arr[23][20] ),
    .S(_04876_),
    .X(_04878_));
 sky130_fd_sc_hd__clkbuf_1 _17236_ (.A(_04878_),
    .X(_01424_));
 sky130_fd_sc_hd__mux2_1 _17237_ (.A0(_14156_),
    .A1(\rvcpu.dp.rf.reg_file_arr[23][19] ),
    .S(_04876_),
    .X(_04879_));
 sky130_fd_sc_hd__clkbuf_1 _17238_ (.A(_04879_),
    .X(_01423_));
 sky130_fd_sc_hd__mux2_1 _17239_ (.A0(_14158_),
    .A1(\rvcpu.dp.rf.reg_file_arr[23][18] ),
    .S(_04876_),
    .X(_04880_));
 sky130_fd_sc_hd__clkbuf_1 _17240_ (.A(_04880_),
    .X(_01422_));
 sky130_fd_sc_hd__mux2_1 _17241_ (.A0(_14160_),
    .A1(\rvcpu.dp.rf.reg_file_arr[23][17] ),
    .S(_04876_),
    .X(_04881_));
 sky130_fd_sc_hd__clkbuf_1 _17242_ (.A(_04881_),
    .X(_01421_));
 sky130_fd_sc_hd__mux2_1 _17243_ (.A0(_14162_),
    .A1(\rvcpu.dp.rf.reg_file_arr[23][16] ),
    .S(_04876_),
    .X(_04882_));
 sky130_fd_sc_hd__clkbuf_1 _17244_ (.A(_04882_),
    .X(_01420_));
 sky130_fd_sc_hd__mux2_1 _17245_ (.A0(_14164_),
    .A1(\rvcpu.dp.rf.reg_file_arr[23][15] ),
    .S(_04876_),
    .X(_04883_));
 sky130_fd_sc_hd__clkbuf_1 _17246_ (.A(_04883_),
    .X(_01419_));
 sky130_fd_sc_hd__mux2_1 _17247_ (.A0(_14166_),
    .A1(\rvcpu.dp.rf.reg_file_arr[23][14] ),
    .S(_04876_),
    .X(_04884_));
 sky130_fd_sc_hd__clkbuf_1 _17248_ (.A(_04884_),
    .X(_01418_));
 sky130_fd_sc_hd__mux2_1 _17249_ (.A0(_14168_),
    .A1(\rvcpu.dp.rf.reg_file_arr[23][13] ),
    .S(_04876_),
    .X(_04885_));
 sky130_fd_sc_hd__clkbuf_1 _17250_ (.A(_04885_),
    .X(_01417_));
 sky130_fd_sc_hd__mux2_1 _17251_ (.A0(_14170_),
    .A1(\rvcpu.dp.rf.reg_file_arr[23][12] ),
    .S(_04876_),
    .X(_04886_));
 sky130_fd_sc_hd__clkbuf_1 _17252_ (.A(_04886_),
    .X(_01416_));
 sky130_fd_sc_hd__clkbuf_4 _17253_ (.A(_04864_),
    .X(_04887_));
 sky130_fd_sc_hd__mux2_1 _17254_ (.A0(_14172_),
    .A1(\rvcpu.dp.rf.reg_file_arr[23][11] ),
    .S(_04887_),
    .X(_04888_));
 sky130_fd_sc_hd__clkbuf_1 _17255_ (.A(_04888_),
    .X(_01415_));
 sky130_fd_sc_hd__mux2_1 _17256_ (.A0(_14175_),
    .A1(\rvcpu.dp.rf.reg_file_arr[23][10] ),
    .S(_04887_),
    .X(_04889_));
 sky130_fd_sc_hd__clkbuf_1 _17257_ (.A(_04889_),
    .X(_01414_));
 sky130_fd_sc_hd__mux2_1 _17258_ (.A0(_14177_),
    .A1(\rvcpu.dp.rf.reg_file_arr[23][9] ),
    .S(_04887_),
    .X(_04890_));
 sky130_fd_sc_hd__clkbuf_1 _17259_ (.A(_04890_),
    .X(_01413_));
 sky130_fd_sc_hd__mux2_1 _17260_ (.A0(_14179_),
    .A1(\rvcpu.dp.rf.reg_file_arr[23][8] ),
    .S(_04887_),
    .X(_04891_));
 sky130_fd_sc_hd__clkbuf_1 _17261_ (.A(_04891_),
    .X(_01412_));
 sky130_fd_sc_hd__mux2_1 _17262_ (.A0(_14181_),
    .A1(\rvcpu.dp.rf.reg_file_arr[23][7] ),
    .S(_04887_),
    .X(_04892_));
 sky130_fd_sc_hd__clkbuf_1 _17263_ (.A(_04892_),
    .X(_01411_));
 sky130_fd_sc_hd__mux2_1 _17264_ (.A0(_14183_),
    .A1(\rvcpu.dp.rf.reg_file_arr[23][6] ),
    .S(_04887_),
    .X(_04893_));
 sky130_fd_sc_hd__clkbuf_1 _17265_ (.A(_04893_),
    .X(_01410_));
 sky130_fd_sc_hd__mux2_1 _17266_ (.A0(_14185_),
    .A1(\rvcpu.dp.rf.reg_file_arr[23][5] ),
    .S(_04887_),
    .X(_04894_));
 sky130_fd_sc_hd__clkbuf_1 _17267_ (.A(_04894_),
    .X(_01409_));
 sky130_fd_sc_hd__mux2_1 _17268_ (.A0(_14187_),
    .A1(\rvcpu.dp.rf.reg_file_arr[23][4] ),
    .S(_04887_),
    .X(_04895_));
 sky130_fd_sc_hd__clkbuf_1 _17269_ (.A(_04895_),
    .X(_01408_));
 sky130_fd_sc_hd__mux2_1 _17270_ (.A0(_14189_),
    .A1(\rvcpu.dp.rf.reg_file_arr[23][3] ),
    .S(_04887_),
    .X(_04896_));
 sky130_fd_sc_hd__clkbuf_1 _17271_ (.A(_04896_),
    .X(_01407_));
 sky130_fd_sc_hd__mux2_1 _17272_ (.A0(_14191_),
    .A1(\rvcpu.dp.rf.reg_file_arr[23][2] ),
    .S(_04887_),
    .X(_04897_));
 sky130_fd_sc_hd__clkbuf_1 _17273_ (.A(_04897_),
    .X(_01406_));
 sky130_fd_sc_hd__mux2_1 _17274_ (.A0(_14193_),
    .A1(\rvcpu.dp.rf.reg_file_arr[23][1] ),
    .S(_04864_),
    .X(_04898_));
 sky130_fd_sc_hd__clkbuf_1 _17275_ (.A(_04898_),
    .X(_01405_));
 sky130_fd_sc_hd__mux2_1 _17276_ (.A0(_14195_),
    .A1(\rvcpu.dp.rf.reg_file_arr[23][0] ),
    .S(_04864_),
    .X(_04899_));
 sky130_fd_sc_hd__clkbuf_1 _17277_ (.A(_04899_),
    .X(_01404_));
 sky130_fd_sc_hd__and3b_1 _17278_ (.A_N(_13174_),
    .B(\rvcpu.dp.plmw.RdW[3] ),
    .C(_13176_),
    .X(_04900_));
 sky130_fd_sc_hd__and2_2 _17279_ (.A(_04464_),
    .B(_04900_),
    .X(_04901_));
 sky130_fd_sc_hd__clkbuf_4 _17280_ (.A(_04901_),
    .X(_04902_));
 sky130_fd_sc_hd__mux2_1 _17281_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][31] ),
    .A1(_13172_),
    .S(_04902_),
    .X(_04903_));
 sky130_fd_sc_hd__clkbuf_1 _17282_ (.A(_04903_),
    .X(_01403_));
 sky130_fd_sc_hd__mux2_1 _17283_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][30] ),
    .A1(_13183_),
    .S(_04902_),
    .X(_04904_));
 sky130_fd_sc_hd__clkbuf_1 _17284_ (.A(_04904_),
    .X(_01402_));
 sky130_fd_sc_hd__mux2_1 _17285_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][29] ),
    .A1(_13186_),
    .S(_04902_),
    .X(_04905_));
 sky130_fd_sc_hd__clkbuf_1 _17286_ (.A(_04905_),
    .X(_01401_));
 sky130_fd_sc_hd__mux2_1 _17287_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][28] ),
    .A1(_13189_),
    .S(_04902_),
    .X(_04906_));
 sky130_fd_sc_hd__clkbuf_1 _17288_ (.A(_04906_),
    .X(_01400_));
 sky130_fd_sc_hd__mux2_1 _17289_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][27] ),
    .A1(_13194_),
    .S(_04902_),
    .X(_04907_));
 sky130_fd_sc_hd__clkbuf_1 _17290_ (.A(_04907_),
    .X(_01399_));
 sky130_fd_sc_hd__mux2_1 _17291_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][26] ),
    .A1(_13197_),
    .S(_04902_),
    .X(_04908_));
 sky130_fd_sc_hd__clkbuf_1 _17292_ (.A(_04908_),
    .X(_01398_));
 sky130_fd_sc_hd__mux2_1 _17293_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][25] ),
    .A1(_13200_),
    .S(_04902_),
    .X(_04909_));
 sky130_fd_sc_hd__clkbuf_1 _17294_ (.A(_04909_),
    .X(_01397_));
 sky130_fd_sc_hd__mux2_1 _17295_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][24] ),
    .A1(_13203_),
    .S(_04902_),
    .X(_04910_));
 sky130_fd_sc_hd__clkbuf_1 _17296_ (.A(_04910_),
    .X(_01396_));
 sky130_fd_sc_hd__mux2_1 _17297_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][23] ),
    .A1(_13206_),
    .S(_04902_),
    .X(_04911_));
 sky130_fd_sc_hd__clkbuf_1 _17298_ (.A(_04911_),
    .X(_01395_));
 sky130_fd_sc_hd__mux2_1 _17299_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][22] ),
    .A1(_13209_),
    .S(_04902_),
    .X(_04912_));
 sky130_fd_sc_hd__clkbuf_1 _17300_ (.A(_04912_),
    .X(_01394_));
 sky130_fd_sc_hd__buf_4 _17301_ (.A(_04901_),
    .X(_04913_));
 sky130_fd_sc_hd__mux2_1 _17302_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][21] ),
    .A1(_13212_),
    .S(_04913_),
    .X(_04914_));
 sky130_fd_sc_hd__clkbuf_1 _17303_ (.A(_04914_),
    .X(_01393_));
 sky130_fd_sc_hd__mux2_1 _17304_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][20] ),
    .A1(_13216_),
    .S(_04913_),
    .X(_04915_));
 sky130_fd_sc_hd__clkbuf_1 _17305_ (.A(_04915_),
    .X(_01392_));
 sky130_fd_sc_hd__mux2_1 _17306_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][19] ),
    .A1(_13219_),
    .S(_04913_),
    .X(_04916_));
 sky130_fd_sc_hd__clkbuf_1 _17307_ (.A(_04916_),
    .X(_01391_));
 sky130_fd_sc_hd__mux2_1 _17308_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][18] ),
    .A1(_13222_),
    .S(_04913_),
    .X(_04917_));
 sky130_fd_sc_hd__clkbuf_1 _17309_ (.A(_04917_),
    .X(_01390_));
 sky130_fd_sc_hd__mux2_1 _17310_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][17] ),
    .A1(_13225_),
    .S(_04913_),
    .X(_04918_));
 sky130_fd_sc_hd__clkbuf_1 _17311_ (.A(_04918_),
    .X(_01389_));
 sky130_fd_sc_hd__mux2_1 _17312_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][16] ),
    .A1(_13228_),
    .S(_04913_),
    .X(_04919_));
 sky130_fd_sc_hd__clkbuf_1 _17313_ (.A(_04919_),
    .X(_01388_));
 sky130_fd_sc_hd__mux2_1 _17314_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][15] ),
    .A1(_13231_),
    .S(_04913_),
    .X(_04920_));
 sky130_fd_sc_hd__clkbuf_1 _17315_ (.A(_04920_),
    .X(_01387_));
 sky130_fd_sc_hd__mux2_1 _17316_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][14] ),
    .A1(_13234_),
    .S(_04913_),
    .X(_04921_));
 sky130_fd_sc_hd__clkbuf_1 _17317_ (.A(_04921_),
    .X(_01386_));
 sky130_fd_sc_hd__mux2_1 _17318_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][13] ),
    .A1(_13237_),
    .S(_04913_),
    .X(_04922_));
 sky130_fd_sc_hd__clkbuf_1 _17319_ (.A(_04922_),
    .X(_01385_));
 sky130_fd_sc_hd__mux2_1 _17320_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][12] ),
    .A1(_13240_),
    .S(_04913_),
    .X(_04923_));
 sky130_fd_sc_hd__clkbuf_1 _17321_ (.A(_04923_),
    .X(_01384_));
 sky130_fd_sc_hd__clkbuf_4 _17322_ (.A(_04901_),
    .X(_04924_));
 sky130_fd_sc_hd__mux2_1 _17323_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][11] ),
    .A1(_13243_),
    .S(_04924_),
    .X(_04925_));
 sky130_fd_sc_hd__clkbuf_1 _17324_ (.A(_04925_),
    .X(_01383_));
 sky130_fd_sc_hd__mux2_1 _17325_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][10] ),
    .A1(_13247_),
    .S(_04924_),
    .X(_04926_));
 sky130_fd_sc_hd__clkbuf_1 _17326_ (.A(_04926_),
    .X(_01382_));
 sky130_fd_sc_hd__mux2_1 _17327_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][9] ),
    .A1(_13250_),
    .S(_04924_),
    .X(_04927_));
 sky130_fd_sc_hd__clkbuf_1 _17328_ (.A(_04927_),
    .X(_01381_));
 sky130_fd_sc_hd__mux2_1 _17329_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][8] ),
    .A1(_13253_),
    .S(_04924_),
    .X(_04928_));
 sky130_fd_sc_hd__clkbuf_1 _17330_ (.A(_04928_),
    .X(_01380_));
 sky130_fd_sc_hd__mux2_1 _17331_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][7] ),
    .A1(_13256_),
    .S(_04924_),
    .X(_04929_));
 sky130_fd_sc_hd__clkbuf_1 _17332_ (.A(_04929_),
    .X(_01379_));
 sky130_fd_sc_hd__mux2_1 _17333_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][6] ),
    .A1(_13259_),
    .S(_04924_),
    .X(_04930_));
 sky130_fd_sc_hd__clkbuf_1 _17334_ (.A(_04930_),
    .X(_01378_));
 sky130_fd_sc_hd__mux2_1 _17335_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][5] ),
    .A1(_13262_),
    .S(_04924_),
    .X(_04931_));
 sky130_fd_sc_hd__clkbuf_1 _17336_ (.A(_04931_),
    .X(_01377_));
 sky130_fd_sc_hd__mux2_1 _17337_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][4] ),
    .A1(_13265_),
    .S(_04924_),
    .X(_04932_));
 sky130_fd_sc_hd__clkbuf_1 _17338_ (.A(_04932_),
    .X(_01376_));
 sky130_fd_sc_hd__mux2_1 _17339_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][3] ),
    .A1(_13268_),
    .S(_04924_),
    .X(_04933_));
 sky130_fd_sc_hd__clkbuf_1 _17340_ (.A(_04933_),
    .X(_01375_));
 sky130_fd_sc_hd__mux2_1 _17341_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][2] ),
    .A1(_13271_),
    .S(_04924_),
    .X(_04934_));
 sky130_fd_sc_hd__clkbuf_1 _17342_ (.A(_04934_),
    .X(_01374_));
 sky130_fd_sc_hd__mux2_1 _17343_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][1] ),
    .A1(_13274_),
    .S(_04901_),
    .X(_04935_));
 sky130_fd_sc_hd__clkbuf_1 _17344_ (.A(_04935_),
    .X(_01373_));
 sky130_fd_sc_hd__mux2_1 _17345_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][0] ),
    .A1(_13277_),
    .S(_04901_),
    .X(_04936_));
 sky130_fd_sc_hd__clkbuf_1 _17346_ (.A(_04936_),
    .X(_01372_));
 sky130_fd_sc_hd__nand2_2 _17347_ (.A(_14128_),
    .B(_04900_),
    .Y(_04937_));
 sky130_fd_sc_hd__clkbuf_4 _17348_ (.A(_04937_),
    .X(_04938_));
 sky130_fd_sc_hd__mux2_1 _17349_ (.A0(_14127_),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][31] ),
    .S(_04938_),
    .X(_04939_));
 sky130_fd_sc_hd__clkbuf_1 _17350_ (.A(_04939_),
    .X(_01363_));
 sky130_fd_sc_hd__mux2_1 _17351_ (.A0(_14133_),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][30] ),
    .S(_04938_),
    .X(_04940_));
 sky130_fd_sc_hd__clkbuf_1 _17352_ (.A(_04940_),
    .X(_01362_));
 sky130_fd_sc_hd__mux2_1 _17353_ (.A0(_14135_),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][29] ),
    .S(_04938_),
    .X(_04941_));
 sky130_fd_sc_hd__clkbuf_1 _17354_ (.A(_04941_),
    .X(_01361_));
 sky130_fd_sc_hd__mux2_1 _17355_ (.A0(_14137_),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][28] ),
    .S(_04938_),
    .X(_04942_));
 sky130_fd_sc_hd__clkbuf_1 _17356_ (.A(_04942_),
    .X(_01360_));
 sky130_fd_sc_hd__mux2_1 _17357_ (.A0(_14139_),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][27] ),
    .S(_04938_),
    .X(_04943_));
 sky130_fd_sc_hd__clkbuf_1 _17358_ (.A(_04943_),
    .X(_01359_));
 sky130_fd_sc_hd__mux2_1 _17359_ (.A0(_14141_),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][26] ),
    .S(_04938_),
    .X(_04944_));
 sky130_fd_sc_hd__clkbuf_1 _17360_ (.A(_04944_),
    .X(_01358_));
 sky130_fd_sc_hd__mux2_1 _17361_ (.A0(_14143_),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][25] ),
    .S(_04938_),
    .X(_04945_));
 sky130_fd_sc_hd__clkbuf_1 _17362_ (.A(_04945_),
    .X(_01357_));
 sky130_fd_sc_hd__mux2_1 _17363_ (.A0(_14145_),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][24] ),
    .S(_04938_),
    .X(_04946_));
 sky130_fd_sc_hd__clkbuf_1 _17364_ (.A(_04946_),
    .X(_01356_));
 sky130_fd_sc_hd__mux2_1 _17365_ (.A0(_14147_),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][23] ),
    .S(_04938_),
    .X(_04947_));
 sky130_fd_sc_hd__clkbuf_1 _17366_ (.A(_04947_),
    .X(_01355_));
 sky130_fd_sc_hd__mux2_1 _17367_ (.A0(_14149_),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][22] ),
    .S(_04938_),
    .X(_04948_));
 sky130_fd_sc_hd__clkbuf_1 _17368_ (.A(_04948_),
    .X(_01354_));
 sky130_fd_sc_hd__buf_4 _17369_ (.A(_04937_),
    .X(_04949_));
 sky130_fd_sc_hd__mux2_1 _17370_ (.A0(_14151_),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][21] ),
    .S(_04949_),
    .X(_04950_));
 sky130_fd_sc_hd__clkbuf_1 _17371_ (.A(_04950_),
    .X(_01353_));
 sky130_fd_sc_hd__mux2_1 _17372_ (.A0(_14154_),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][20] ),
    .S(_04949_),
    .X(_04951_));
 sky130_fd_sc_hd__clkbuf_1 _17373_ (.A(_04951_),
    .X(_01352_));
 sky130_fd_sc_hd__mux2_1 _17374_ (.A0(_14156_),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][19] ),
    .S(_04949_),
    .X(_04952_));
 sky130_fd_sc_hd__clkbuf_1 _17375_ (.A(_04952_),
    .X(_01351_));
 sky130_fd_sc_hd__mux2_1 _17376_ (.A0(_14158_),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][18] ),
    .S(_04949_),
    .X(_04953_));
 sky130_fd_sc_hd__clkbuf_1 _17377_ (.A(_04953_),
    .X(_01350_));
 sky130_fd_sc_hd__mux2_1 _17378_ (.A0(_14160_),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][17] ),
    .S(_04949_),
    .X(_04954_));
 sky130_fd_sc_hd__clkbuf_1 _17379_ (.A(_04954_),
    .X(_01349_));
 sky130_fd_sc_hd__mux2_1 _17380_ (.A0(_14162_),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][16] ),
    .S(_04949_),
    .X(_04955_));
 sky130_fd_sc_hd__clkbuf_1 _17381_ (.A(_04955_),
    .X(_01348_));
 sky130_fd_sc_hd__mux2_1 _17382_ (.A0(_14164_),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][15] ),
    .S(_04949_),
    .X(_04956_));
 sky130_fd_sc_hd__clkbuf_1 _17383_ (.A(_04956_),
    .X(_01347_));
 sky130_fd_sc_hd__mux2_1 _17384_ (.A0(_14166_),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][14] ),
    .S(_04949_),
    .X(_04957_));
 sky130_fd_sc_hd__clkbuf_1 _17385_ (.A(_04957_),
    .X(_01346_));
 sky130_fd_sc_hd__mux2_1 _17386_ (.A0(_14168_),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][13] ),
    .S(_04949_),
    .X(_04958_));
 sky130_fd_sc_hd__clkbuf_1 _17387_ (.A(_04958_),
    .X(_01345_));
 sky130_fd_sc_hd__mux2_1 _17388_ (.A0(_14170_),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][12] ),
    .S(_04949_),
    .X(_04959_));
 sky130_fd_sc_hd__clkbuf_1 _17389_ (.A(_04959_),
    .X(_01344_));
 sky130_fd_sc_hd__clkbuf_4 _17390_ (.A(_04937_),
    .X(_04960_));
 sky130_fd_sc_hd__mux2_1 _17391_ (.A0(_14172_),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][11] ),
    .S(_04960_),
    .X(_04961_));
 sky130_fd_sc_hd__clkbuf_1 _17392_ (.A(_04961_),
    .X(_01343_));
 sky130_fd_sc_hd__mux2_1 _17393_ (.A0(_14175_),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][10] ),
    .S(_04960_),
    .X(_04962_));
 sky130_fd_sc_hd__clkbuf_1 _17394_ (.A(_04962_),
    .X(_01342_));
 sky130_fd_sc_hd__mux2_1 _17395_ (.A0(_14177_),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][9] ),
    .S(_04960_),
    .X(_04963_));
 sky130_fd_sc_hd__clkbuf_1 _17396_ (.A(_04963_),
    .X(_01341_));
 sky130_fd_sc_hd__mux2_1 _17397_ (.A0(_14179_),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][8] ),
    .S(_04960_),
    .X(_04964_));
 sky130_fd_sc_hd__clkbuf_1 _17398_ (.A(_04964_),
    .X(_01340_));
 sky130_fd_sc_hd__mux2_1 _17399_ (.A0(_14181_),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][7] ),
    .S(_04960_),
    .X(_04965_));
 sky130_fd_sc_hd__clkbuf_1 _17400_ (.A(_04965_),
    .X(_01339_));
 sky130_fd_sc_hd__mux2_1 _17401_ (.A0(_14183_),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][6] ),
    .S(_04960_),
    .X(_04966_));
 sky130_fd_sc_hd__clkbuf_1 _17402_ (.A(_04966_),
    .X(_01338_));
 sky130_fd_sc_hd__mux2_1 _17403_ (.A0(_14185_),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][5] ),
    .S(_04960_),
    .X(_04967_));
 sky130_fd_sc_hd__clkbuf_1 _17404_ (.A(_04967_),
    .X(_01337_));
 sky130_fd_sc_hd__mux2_1 _17405_ (.A0(_14187_),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][4] ),
    .S(_04960_),
    .X(_04968_));
 sky130_fd_sc_hd__clkbuf_1 _17406_ (.A(_04968_),
    .X(_01336_));
 sky130_fd_sc_hd__mux2_1 _17407_ (.A0(_14189_),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][3] ),
    .S(_04960_),
    .X(_04969_));
 sky130_fd_sc_hd__clkbuf_1 _17408_ (.A(_04969_),
    .X(_01335_));
 sky130_fd_sc_hd__mux2_1 _17409_ (.A0(_14191_),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][2] ),
    .S(_04960_),
    .X(_04970_));
 sky130_fd_sc_hd__clkbuf_1 _17410_ (.A(_04970_),
    .X(_01334_));
 sky130_fd_sc_hd__mux2_1 _17411_ (.A0(_14193_),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][1] ),
    .S(_04937_),
    .X(_04971_));
 sky130_fd_sc_hd__clkbuf_1 _17412_ (.A(_04971_),
    .X(_01333_));
 sky130_fd_sc_hd__mux2_1 _17413_ (.A0(_14195_),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][0] ),
    .S(_04937_),
    .X(_04972_));
 sky130_fd_sc_hd__clkbuf_1 _17414_ (.A(_04972_),
    .X(_01332_));
 sky130_fd_sc_hd__nand2_2 _17415_ (.A(_04538_),
    .B(_04900_),
    .Y(_04973_));
 sky130_fd_sc_hd__clkbuf_4 _17416_ (.A(_04973_),
    .X(_04974_));
 sky130_fd_sc_hd__mux2_1 _17417_ (.A0(_14127_),
    .A1(\rvcpu.dp.rf.reg_file_arr[26][31] ),
    .S(_04974_),
    .X(_04975_));
 sky130_fd_sc_hd__clkbuf_1 _17418_ (.A(_04975_),
    .X(_01331_));
 sky130_fd_sc_hd__mux2_1 _17419_ (.A0(_14133_),
    .A1(\rvcpu.dp.rf.reg_file_arr[26][30] ),
    .S(_04974_),
    .X(_04976_));
 sky130_fd_sc_hd__clkbuf_1 _17420_ (.A(_04976_),
    .X(_01330_));
 sky130_fd_sc_hd__mux2_1 _17421_ (.A0(_14135_),
    .A1(\rvcpu.dp.rf.reg_file_arr[26][29] ),
    .S(_04974_),
    .X(_04977_));
 sky130_fd_sc_hd__clkbuf_1 _17422_ (.A(_04977_),
    .X(_01329_));
 sky130_fd_sc_hd__mux2_1 _17423_ (.A0(_14137_),
    .A1(\rvcpu.dp.rf.reg_file_arr[26][28] ),
    .S(_04974_),
    .X(_04978_));
 sky130_fd_sc_hd__clkbuf_1 _17424_ (.A(_04978_),
    .X(_01328_));
 sky130_fd_sc_hd__mux2_1 _17425_ (.A0(_14139_),
    .A1(\rvcpu.dp.rf.reg_file_arr[26][27] ),
    .S(_04974_),
    .X(_04979_));
 sky130_fd_sc_hd__clkbuf_1 _17426_ (.A(_04979_),
    .X(_01327_));
 sky130_fd_sc_hd__mux2_1 _17427_ (.A0(_14141_),
    .A1(\rvcpu.dp.rf.reg_file_arr[26][26] ),
    .S(_04974_),
    .X(_04980_));
 sky130_fd_sc_hd__clkbuf_1 _17428_ (.A(_04980_),
    .X(_01326_));
 sky130_fd_sc_hd__mux2_1 _17429_ (.A0(_14143_),
    .A1(\rvcpu.dp.rf.reg_file_arr[26][25] ),
    .S(_04974_),
    .X(_04981_));
 sky130_fd_sc_hd__clkbuf_1 _17430_ (.A(_04981_),
    .X(_01325_));
 sky130_fd_sc_hd__mux2_1 _17431_ (.A0(_14145_),
    .A1(\rvcpu.dp.rf.reg_file_arr[26][24] ),
    .S(_04974_),
    .X(_04982_));
 sky130_fd_sc_hd__clkbuf_1 _17432_ (.A(_04982_),
    .X(_01324_));
 sky130_fd_sc_hd__mux2_1 _17433_ (.A0(_14147_),
    .A1(\rvcpu.dp.rf.reg_file_arr[26][23] ),
    .S(_04974_),
    .X(_04983_));
 sky130_fd_sc_hd__clkbuf_1 _17434_ (.A(_04983_),
    .X(_01323_));
 sky130_fd_sc_hd__mux2_1 _17435_ (.A0(_14149_),
    .A1(\rvcpu.dp.rf.reg_file_arr[26][22] ),
    .S(_04974_),
    .X(_04984_));
 sky130_fd_sc_hd__clkbuf_1 _17436_ (.A(_04984_),
    .X(_01322_));
 sky130_fd_sc_hd__buf_4 _17437_ (.A(_04973_),
    .X(_04985_));
 sky130_fd_sc_hd__mux2_1 _17438_ (.A0(_14151_),
    .A1(\rvcpu.dp.rf.reg_file_arr[26][21] ),
    .S(_04985_),
    .X(_04986_));
 sky130_fd_sc_hd__clkbuf_1 _17439_ (.A(_04986_),
    .X(_01321_));
 sky130_fd_sc_hd__mux2_1 _17440_ (.A0(_14154_),
    .A1(\rvcpu.dp.rf.reg_file_arr[26][20] ),
    .S(_04985_),
    .X(_04987_));
 sky130_fd_sc_hd__clkbuf_1 _17441_ (.A(_04987_),
    .X(_01320_));
 sky130_fd_sc_hd__mux2_1 _17442_ (.A0(_14156_),
    .A1(\rvcpu.dp.rf.reg_file_arr[26][19] ),
    .S(_04985_),
    .X(_04988_));
 sky130_fd_sc_hd__clkbuf_1 _17443_ (.A(_04988_),
    .X(_01319_));
 sky130_fd_sc_hd__mux2_1 _17444_ (.A0(_14158_),
    .A1(\rvcpu.dp.rf.reg_file_arr[26][18] ),
    .S(_04985_),
    .X(_04989_));
 sky130_fd_sc_hd__clkbuf_1 _17445_ (.A(_04989_),
    .X(_01318_));
 sky130_fd_sc_hd__mux2_1 _17446_ (.A0(_14160_),
    .A1(\rvcpu.dp.rf.reg_file_arr[26][17] ),
    .S(_04985_),
    .X(_04990_));
 sky130_fd_sc_hd__clkbuf_1 _17447_ (.A(_04990_),
    .X(_01317_));
 sky130_fd_sc_hd__mux2_1 _17448_ (.A0(_14162_),
    .A1(\rvcpu.dp.rf.reg_file_arr[26][16] ),
    .S(_04985_),
    .X(_04991_));
 sky130_fd_sc_hd__clkbuf_1 _17449_ (.A(_04991_),
    .X(_01316_));
 sky130_fd_sc_hd__mux2_1 _17450_ (.A0(_14164_),
    .A1(\rvcpu.dp.rf.reg_file_arr[26][15] ),
    .S(_04985_),
    .X(_04992_));
 sky130_fd_sc_hd__clkbuf_1 _17451_ (.A(_04992_),
    .X(_01315_));
 sky130_fd_sc_hd__mux2_1 _17452_ (.A0(_14166_),
    .A1(\rvcpu.dp.rf.reg_file_arr[26][14] ),
    .S(_04985_),
    .X(_04993_));
 sky130_fd_sc_hd__clkbuf_1 _17453_ (.A(_04993_),
    .X(_01314_));
 sky130_fd_sc_hd__mux2_1 _17454_ (.A0(_14168_),
    .A1(\rvcpu.dp.rf.reg_file_arr[26][13] ),
    .S(_04985_),
    .X(_04994_));
 sky130_fd_sc_hd__clkbuf_1 _17455_ (.A(_04994_),
    .X(_01313_));
 sky130_fd_sc_hd__mux2_1 _17456_ (.A0(_14170_),
    .A1(\rvcpu.dp.rf.reg_file_arr[26][12] ),
    .S(_04985_),
    .X(_04995_));
 sky130_fd_sc_hd__clkbuf_1 _17457_ (.A(_04995_),
    .X(_01312_));
 sky130_fd_sc_hd__clkbuf_4 _17458_ (.A(_04973_),
    .X(_04996_));
 sky130_fd_sc_hd__mux2_1 _17459_ (.A0(_14172_),
    .A1(\rvcpu.dp.rf.reg_file_arr[26][11] ),
    .S(_04996_),
    .X(_04997_));
 sky130_fd_sc_hd__clkbuf_1 _17460_ (.A(_04997_),
    .X(_01311_));
 sky130_fd_sc_hd__mux2_1 _17461_ (.A0(_14175_),
    .A1(\rvcpu.dp.rf.reg_file_arr[26][10] ),
    .S(_04996_),
    .X(_04998_));
 sky130_fd_sc_hd__clkbuf_1 _17462_ (.A(_04998_),
    .X(_01310_));
 sky130_fd_sc_hd__mux2_1 _17463_ (.A0(_14177_),
    .A1(\rvcpu.dp.rf.reg_file_arr[26][9] ),
    .S(_04996_),
    .X(_04999_));
 sky130_fd_sc_hd__clkbuf_1 _17464_ (.A(_04999_),
    .X(_01309_));
 sky130_fd_sc_hd__mux2_1 _17465_ (.A0(_14179_),
    .A1(\rvcpu.dp.rf.reg_file_arr[26][8] ),
    .S(_04996_),
    .X(_05000_));
 sky130_fd_sc_hd__clkbuf_1 _17466_ (.A(_05000_),
    .X(_01308_));
 sky130_fd_sc_hd__mux2_1 _17467_ (.A0(_14181_),
    .A1(\rvcpu.dp.rf.reg_file_arr[26][7] ),
    .S(_04996_),
    .X(_05001_));
 sky130_fd_sc_hd__clkbuf_1 _17468_ (.A(_05001_),
    .X(_01307_));
 sky130_fd_sc_hd__mux2_1 _17469_ (.A0(_14183_),
    .A1(\rvcpu.dp.rf.reg_file_arr[26][6] ),
    .S(_04996_),
    .X(_05002_));
 sky130_fd_sc_hd__clkbuf_1 _17470_ (.A(_05002_),
    .X(_01306_));
 sky130_fd_sc_hd__mux2_1 _17471_ (.A0(_14185_),
    .A1(\rvcpu.dp.rf.reg_file_arr[26][5] ),
    .S(_04996_),
    .X(_05003_));
 sky130_fd_sc_hd__clkbuf_1 _17472_ (.A(_05003_),
    .X(_01305_));
 sky130_fd_sc_hd__mux2_1 _17473_ (.A0(_14187_),
    .A1(\rvcpu.dp.rf.reg_file_arr[26][4] ),
    .S(_04996_),
    .X(_05004_));
 sky130_fd_sc_hd__clkbuf_1 _17474_ (.A(_05004_),
    .X(_01304_));
 sky130_fd_sc_hd__mux2_1 _17475_ (.A0(_14189_),
    .A1(\rvcpu.dp.rf.reg_file_arr[26][3] ),
    .S(_04996_),
    .X(_05005_));
 sky130_fd_sc_hd__clkbuf_1 _17476_ (.A(_05005_),
    .X(_01303_));
 sky130_fd_sc_hd__mux2_1 _17477_ (.A0(_14191_),
    .A1(\rvcpu.dp.rf.reg_file_arr[26][2] ),
    .S(_04996_),
    .X(_05006_));
 sky130_fd_sc_hd__clkbuf_1 _17478_ (.A(_05006_),
    .X(_01302_));
 sky130_fd_sc_hd__mux2_1 _17479_ (.A0(_14193_),
    .A1(\rvcpu.dp.rf.reg_file_arr[26][1] ),
    .S(_04973_),
    .X(_05007_));
 sky130_fd_sc_hd__clkbuf_1 _17480_ (.A(_05007_),
    .X(_01301_));
 sky130_fd_sc_hd__mux2_1 _17481_ (.A0(_14195_),
    .A1(\rvcpu.dp.rf.reg_file_arr[26][0] ),
    .S(_04973_),
    .X(_05008_));
 sky130_fd_sc_hd__clkbuf_1 _17482_ (.A(_05008_),
    .X(_01300_));
 sky130_fd_sc_hd__nand2_2 _17483_ (.A(_14197_),
    .B(_04900_),
    .Y(_05009_));
 sky130_fd_sc_hd__clkbuf_4 _17484_ (.A(_05009_),
    .X(_05010_));
 sky130_fd_sc_hd__mux2_1 _17485_ (.A0(_13173_),
    .A1(\rvcpu.dp.rf.reg_file_arr[27][31] ),
    .S(_05010_),
    .X(_05011_));
 sky130_fd_sc_hd__clkbuf_1 _17486_ (.A(_05011_),
    .X(_01299_));
 sky130_fd_sc_hd__mux2_1 _17487_ (.A0(_13184_),
    .A1(\rvcpu.dp.rf.reg_file_arr[27][30] ),
    .S(_05010_),
    .X(_05012_));
 sky130_fd_sc_hd__clkbuf_1 _17488_ (.A(_05012_),
    .X(_01298_));
 sky130_fd_sc_hd__mux2_1 _17489_ (.A0(_13187_),
    .A1(\rvcpu.dp.rf.reg_file_arr[27][29] ),
    .S(_05010_),
    .X(_05013_));
 sky130_fd_sc_hd__clkbuf_1 _17490_ (.A(_05013_),
    .X(_01297_));
 sky130_fd_sc_hd__mux2_1 _17491_ (.A0(_13190_),
    .A1(\rvcpu.dp.rf.reg_file_arr[27][28] ),
    .S(_05010_),
    .X(_05014_));
 sky130_fd_sc_hd__clkbuf_1 _17492_ (.A(_05014_),
    .X(_01296_));
 sky130_fd_sc_hd__mux2_1 _17493_ (.A0(_13195_),
    .A1(\rvcpu.dp.rf.reg_file_arr[27][27] ),
    .S(_05010_),
    .X(_05015_));
 sky130_fd_sc_hd__clkbuf_1 _17494_ (.A(_05015_),
    .X(_01295_));
 sky130_fd_sc_hd__mux2_1 _17495_ (.A0(_13198_),
    .A1(\rvcpu.dp.rf.reg_file_arr[27][26] ),
    .S(_05010_),
    .X(_05016_));
 sky130_fd_sc_hd__clkbuf_1 _17496_ (.A(_05016_),
    .X(_01294_));
 sky130_fd_sc_hd__mux2_1 _17497_ (.A0(_13201_),
    .A1(\rvcpu.dp.rf.reg_file_arr[27][25] ),
    .S(_05010_),
    .X(_05017_));
 sky130_fd_sc_hd__clkbuf_1 _17498_ (.A(_05017_),
    .X(_01293_));
 sky130_fd_sc_hd__mux2_1 _17499_ (.A0(_13204_),
    .A1(\rvcpu.dp.rf.reg_file_arr[27][24] ),
    .S(_05010_),
    .X(_05018_));
 sky130_fd_sc_hd__clkbuf_1 _17500_ (.A(_05018_),
    .X(_01292_));
 sky130_fd_sc_hd__mux2_1 _17501_ (.A0(_13207_),
    .A1(\rvcpu.dp.rf.reg_file_arr[27][23] ),
    .S(_05010_),
    .X(_05019_));
 sky130_fd_sc_hd__clkbuf_1 _17502_ (.A(_05019_),
    .X(_01291_));
 sky130_fd_sc_hd__mux2_1 _17503_ (.A0(_13210_),
    .A1(\rvcpu.dp.rf.reg_file_arr[27][22] ),
    .S(_05010_),
    .X(_05020_));
 sky130_fd_sc_hd__clkbuf_1 _17504_ (.A(_05020_),
    .X(_01290_));
 sky130_fd_sc_hd__buf_4 _17505_ (.A(_05009_),
    .X(_05021_));
 sky130_fd_sc_hd__mux2_1 _17506_ (.A0(_13213_),
    .A1(\rvcpu.dp.rf.reg_file_arr[27][21] ),
    .S(_05021_),
    .X(_05022_));
 sky130_fd_sc_hd__clkbuf_1 _17507_ (.A(_05022_),
    .X(_01289_));
 sky130_fd_sc_hd__mux2_1 _17508_ (.A0(_13217_),
    .A1(\rvcpu.dp.rf.reg_file_arr[27][20] ),
    .S(_05021_),
    .X(_05023_));
 sky130_fd_sc_hd__clkbuf_1 _17509_ (.A(_05023_),
    .X(_01288_));
 sky130_fd_sc_hd__mux2_1 _17510_ (.A0(_13220_),
    .A1(\rvcpu.dp.rf.reg_file_arr[27][19] ),
    .S(_05021_),
    .X(_05024_));
 sky130_fd_sc_hd__clkbuf_1 _17511_ (.A(_05024_),
    .X(_01287_));
 sky130_fd_sc_hd__mux2_1 _17512_ (.A0(_13223_),
    .A1(\rvcpu.dp.rf.reg_file_arr[27][18] ),
    .S(_05021_),
    .X(_05025_));
 sky130_fd_sc_hd__clkbuf_1 _17513_ (.A(_05025_),
    .X(_01286_));
 sky130_fd_sc_hd__mux2_1 _17514_ (.A0(_13226_),
    .A1(\rvcpu.dp.rf.reg_file_arr[27][17] ),
    .S(_05021_),
    .X(_05026_));
 sky130_fd_sc_hd__clkbuf_1 _17515_ (.A(_05026_),
    .X(_01285_));
 sky130_fd_sc_hd__mux2_1 _17516_ (.A0(_13229_),
    .A1(\rvcpu.dp.rf.reg_file_arr[27][16] ),
    .S(_05021_),
    .X(_05027_));
 sky130_fd_sc_hd__clkbuf_1 _17517_ (.A(_05027_),
    .X(_01284_));
 sky130_fd_sc_hd__mux2_1 _17518_ (.A0(_13232_),
    .A1(\rvcpu.dp.rf.reg_file_arr[27][15] ),
    .S(_05021_),
    .X(_05028_));
 sky130_fd_sc_hd__clkbuf_1 _17519_ (.A(_05028_),
    .X(_01283_));
 sky130_fd_sc_hd__mux2_1 _17520_ (.A0(_13235_),
    .A1(\rvcpu.dp.rf.reg_file_arr[27][14] ),
    .S(_05021_),
    .X(_05029_));
 sky130_fd_sc_hd__clkbuf_1 _17521_ (.A(_05029_),
    .X(_01282_));
 sky130_fd_sc_hd__mux2_1 _17522_ (.A0(_13238_),
    .A1(\rvcpu.dp.rf.reg_file_arr[27][13] ),
    .S(_05021_),
    .X(_05030_));
 sky130_fd_sc_hd__clkbuf_1 _17523_ (.A(_05030_),
    .X(_01281_));
 sky130_fd_sc_hd__mux2_1 _17524_ (.A0(_13241_),
    .A1(\rvcpu.dp.rf.reg_file_arr[27][12] ),
    .S(_05021_),
    .X(_05031_));
 sky130_fd_sc_hd__clkbuf_1 _17525_ (.A(_05031_),
    .X(_01280_));
 sky130_fd_sc_hd__clkbuf_4 _17526_ (.A(_05009_),
    .X(_05032_));
 sky130_fd_sc_hd__mux2_1 _17527_ (.A0(_13244_),
    .A1(\rvcpu.dp.rf.reg_file_arr[27][11] ),
    .S(_05032_),
    .X(_05033_));
 sky130_fd_sc_hd__clkbuf_1 _17528_ (.A(_05033_),
    .X(_01279_));
 sky130_fd_sc_hd__mux2_1 _17529_ (.A0(_13248_),
    .A1(\rvcpu.dp.rf.reg_file_arr[27][10] ),
    .S(_05032_),
    .X(_05034_));
 sky130_fd_sc_hd__clkbuf_1 _17530_ (.A(_05034_),
    .X(_01278_));
 sky130_fd_sc_hd__mux2_1 _17531_ (.A0(_13251_),
    .A1(\rvcpu.dp.rf.reg_file_arr[27][9] ),
    .S(_05032_),
    .X(_05035_));
 sky130_fd_sc_hd__clkbuf_1 _17532_ (.A(_05035_),
    .X(_01277_));
 sky130_fd_sc_hd__mux2_1 _17533_ (.A0(_13254_),
    .A1(\rvcpu.dp.rf.reg_file_arr[27][8] ),
    .S(_05032_),
    .X(_05036_));
 sky130_fd_sc_hd__clkbuf_1 _17534_ (.A(_05036_),
    .X(_01276_));
 sky130_fd_sc_hd__mux2_1 _17535_ (.A0(_13257_),
    .A1(\rvcpu.dp.rf.reg_file_arr[27][7] ),
    .S(_05032_),
    .X(_05037_));
 sky130_fd_sc_hd__clkbuf_1 _17536_ (.A(_05037_),
    .X(_01275_));
 sky130_fd_sc_hd__mux2_1 _17537_ (.A0(_13260_),
    .A1(\rvcpu.dp.rf.reg_file_arr[27][6] ),
    .S(_05032_),
    .X(_05038_));
 sky130_fd_sc_hd__clkbuf_1 _17538_ (.A(_05038_),
    .X(_01274_));
 sky130_fd_sc_hd__mux2_1 _17539_ (.A0(_13263_),
    .A1(\rvcpu.dp.rf.reg_file_arr[27][5] ),
    .S(_05032_),
    .X(_05039_));
 sky130_fd_sc_hd__clkbuf_1 _17540_ (.A(_05039_),
    .X(_01273_));
 sky130_fd_sc_hd__mux2_1 _17541_ (.A0(_13266_),
    .A1(\rvcpu.dp.rf.reg_file_arr[27][4] ),
    .S(_05032_),
    .X(_05040_));
 sky130_fd_sc_hd__clkbuf_1 _17542_ (.A(_05040_),
    .X(_01272_));
 sky130_fd_sc_hd__mux2_1 _17543_ (.A0(_13269_),
    .A1(\rvcpu.dp.rf.reg_file_arr[27][3] ),
    .S(_05032_),
    .X(_05041_));
 sky130_fd_sc_hd__clkbuf_1 _17544_ (.A(_05041_),
    .X(_01271_));
 sky130_fd_sc_hd__mux2_1 _17545_ (.A0(_13272_),
    .A1(\rvcpu.dp.rf.reg_file_arr[27][2] ),
    .S(_05032_),
    .X(_05042_));
 sky130_fd_sc_hd__clkbuf_1 _17546_ (.A(_05042_),
    .X(_01270_));
 sky130_fd_sc_hd__mux2_1 _17547_ (.A0(_13275_),
    .A1(\rvcpu.dp.rf.reg_file_arr[27][1] ),
    .S(_05009_),
    .X(_05043_));
 sky130_fd_sc_hd__clkbuf_1 _17548_ (.A(_05043_),
    .X(_01269_));
 sky130_fd_sc_hd__mux2_1 _17549_ (.A0(_13278_),
    .A1(\rvcpu.dp.rf.reg_file_arr[27][0] ),
    .S(_05009_),
    .X(_05044_));
 sky130_fd_sc_hd__clkbuf_1 _17550_ (.A(_05044_),
    .X(_01268_));
 sky130_fd_sc_hd__nand2_2 _17551_ (.A(_14129_),
    .B(_04464_),
    .Y(_05045_));
 sky130_fd_sc_hd__clkbuf_4 _17552_ (.A(_05045_),
    .X(_05046_));
 sky130_fd_sc_hd__mux2_1 _17553_ (.A0(_13173_),
    .A1(\rvcpu.dp.rf.reg_file_arr[28][31] ),
    .S(_05046_),
    .X(_05047_));
 sky130_fd_sc_hd__clkbuf_1 _17554_ (.A(_05047_),
    .X(_01259_));
 sky130_fd_sc_hd__mux2_1 _17555_ (.A0(_13184_),
    .A1(\rvcpu.dp.rf.reg_file_arr[28][30] ),
    .S(_05046_),
    .X(_05048_));
 sky130_fd_sc_hd__clkbuf_1 _17556_ (.A(_05048_),
    .X(_01258_));
 sky130_fd_sc_hd__mux2_1 _17557_ (.A0(_13187_),
    .A1(\rvcpu.dp.rf.reg_file_arr[28][29] ),
    .S(_05046_),
    .X(_05049_));
 sky130_fd_sc_hd__clkbuf_1 _17558_ (.A(_05049_),
    .X(_01257_));
 sky130_fd_sc_hd__mux2_1 _17559_ (.A0(_13190_),
    .A1(\rvcpu.dp.rf.reg_file_arr[28][28] ),
    .S(_05046_),
    .X(_05050_));
 sky130_fd_sc_hd__clkbuf_1 _17560_ (.A(_05050_),
    .X(_01256_));
 sky130_fd_sc_hd__mux2_1 _17561_ (.A0(_13195_),
    .A1(\rvcpu.dp.rf.reg_file_arr[28][27] ),
    .S(_05046_),
    .X(_05051_));
 sky130_fd_sc_hd__clkbuf_1 _17562_ (.A(_05051_),
    .X(_01255_));
 sky130_fd_sc_hd__mux2_1 _17563_ (.A0(_13198_),
    .A1(\rvcpu.dp.rf.reg_file_arr[28][26] ),
    .S(_05046_),
    .X(_05052_));
 sky130_fd_sc_hd__clkbuf_1 _17564_ (.A(_05052_),
    .X(_01254_));
 sky130_fd_sc_hd__mux2_1 _17565_ (.A0(_13201_),
    .A1(\rvcpu.dp.rf.reg_file_arr[28][25] ),
    .S(_05046_),
    .X(_05053_));
 sky130_fd_sc_hd__clkbuf_1 _17566_ (.A(_05053_),
    .X(_01253_));
 sky130_fd_sc_hd__mux2_1 _17567_ (.A0(_13204_),
    .A1(\rvcpu.dp.rf.reg_file_arr[28][24] ),
    .S(_05046_),
    .X(_05054_));
 sky130_fd_sc_hd__clkbuf_1 _17568_ (.A(_05054_),
    .X(_01252_));
 sky130_fd_sc_hd__mux2_1 _17569_ (.A0(_13207_),
    .A1(\rvcpu.dp.rf.reg_file_arr[28][23] ),
    .S(_05046_),
    .X(_05055_));
 sky130_fd_sc_hd__clkbuf_1 _17570_ (.A(_05055_),
    .X(_01251_));
 sky130_fd_sc_hd__mux2_1 _17571_ (.A0(_13210_),
    .A1(\rvcpu.dp.rf.reg_file_arr[28][22] ),
    .S(_05046_),
    .X(_05056_));
 sky130_fd_sc_hd__clkbuf_1 _17572_ (.A(_05056_),
    .X(_01250_));
 sky130_fd_sc_hd__clkbuf_4 _17573_ (.A(_05045_),
    .X(_05057_));
 sky130_fd_sc_hd__mux2_1 _17574_ (.A0(_13213_),
    .A1(\rvcpu.dp.rf.reg_file_arr[28][21] ),
    .S(_05057_),
    .X(_05058_));
 sky130_fd_sc_hd__clkbuf_1 _17575_ (.A(_05058_),
    .X(_01249_));
 sky130_fd_sc_hd__mux2_1 _17576_ (.A0(_13217_),
    .A1(\rvcpu.dp.rf.reg_file_arr[28][20] ),
    .S(_05057_),
    .X(_05059_));
 sky130_fd_sc_hd__clkbuf_1 _17577_ (.A(_05059_),
    .X(_01248_));
 sky130_fd_sc_hd__mux2_1 _17578_ (.A0(_13220_),
    .A1(\rvcpu.dp.rf.reg_file_arr[28][19] ),
    .S(_05057_),
    .X(_05060_));
 sky130_fd_sc_hd__clkbuf_1 _17579_ (.A(_05060_),
    .X(_01247_));
 sky130_fd_sc_hd__mux2_1 _17580_ (.A0(_13223_),
    .A1(\rvcpu.dp.rf.reg_file_arr[28][18] ),
    .S(_05057_),
    .X(_05061_));
 sky130_fd_sc_hd__clkbuf_1 _17581_ (.A(_05061_),
    .X(_01246_));
 sky130_fd_sc_hd__mux2_1 _17582_ (.A0(_13226_),
    .A1(\rvcpu.dp.rf.reg_file_arr[28][17] ),
    .S(_05057_),
    .X(_05062_));
 sky130_fd_sc_hd__clkbuf_1 _17583_ (.A(_05062_),
    .X(_01245_));
 sky130_fd_sc_hd__mux2_1 _17584_ (.A0(_13229_),
    .A1(\rvcpu.dp.rf.reg_file_arr[28][16] ),
    .S(_05057_),
    .X(_05063_));
 sky130_fd_sc_hd__clkbuf_1 _17585_ (.A(_05063_),
    .X(_01244_));
 sky130_fd_sc_hd__mux2_1 _17586_ (.A0(_13232_),
    .A1(\rvcpu.dp.rf.reg_file_arr[28][15] ),
    .S(_05057_),
    .X(_05064_));
 sky130_fd_sc_hd__clkbuf_1 _17587_ (.A(_05064_),
    .X(_01243_));
 sky130_fd_sc_hd__mux2_1 _17588_ (.A0(_13235_),
    .A1(\rvcpu.dp.rf.reg_file_arr[28][14] ),
    .S(_05057_),
    .X(_05065_));
 sky130_fd_sc_hd__clkbuf_1 _17589_ (.A(_05065_),
    .X(_01242_));
 sky130_fd_sc_hd__mux2_1 _17590_ (.A0(_13238_),
    .A1(\rvcpu.dp.rf.reg_file_arr[28][13] ),
    .S(_05057_),
    .X(_05066_));
 sky130_fd_sc_hd__clkbuf_1 _17591_ (.A(_05066_),
    .X(_01241_));
 sky130_fd_sc_hd__mux2_1 _17592_ (.A0(_13241_),
    .A1(\rvcpu.dp.rf.reg_file_arr[28][12] ),
    .S(_05057_),
    .X(_05067_));
 sky130_fd_sc_hd__clkbuf_1 _17593_ (.A(_05067_),
    .X(_01240_));
 sky130_fd_sc_hd__buf_4 _17594_ (.A(_05045_),
    .X(_05068_));
 sky130_fd_sc_hd__mux2_1 _17595_ (.A0(_13244_),
    .A1(\rvcpu.dp.rf.reg_file_arr[28][11] ),
    .S(_05068_),
    .X(_05069_));
 sky130_fd_sc_hd__clkbuf_1 _17596_ (.A(_05069_),
    .X(_01239_));
 sky130_fd_sc_hd__mux2_1 _17597_ (.A0(_13248_),
    .A1(\rvcpu.dp.rf.reg_file_arr[28][10] ),
    .S(_05068_),
    .X(_05070_));
 sky130_fd_sc_hd__clkbuf_1 _17598_ (.A(_05070_),
    .X(_01238_));
 sky130_fd_sc_hd__mux2_1 _17599_ (.A0(_13251_),
    .A1(\rvcpu.dp.rf.reg_file_arr[28][9] ),
    .S(_05068_),
    .X(_05071_));
 sky130_fd_sc_hd__clkbuf_1 _17600_ (.A(_05071_),
    .X(_01237_));
 sky130_fd_sc_hd__mux2_1 _17601_ (.A0(_13254_),
    .A1(\rvcpu.dp.rf.reg_file_arr[28][8] ),
    .S(_05068_),
    .X(_05072_));
 sky130_fd_sc_hd__clkbuf_1 _17602_ (.A(_05072_),
    .X(_01236_));
 sky130_fd_sc_hd__mux2_1 _17603_ (.A0(_13257_),
    .A1(\rvcpu.dp.rf.reg_file_arr[28][7] ),
    .S(_05068_),
    .X(_05073_));
 sky130_fd_sc_hd__clkbuf_1 _17604_ (.A(_05073_),
    .X(_01235_));
 sky130_fd_sc_hd__mux2_1 _17605_ (.A0(_13260_),
    .A1(\rvcpu.dp.rf.reg_file_arr[28][6] ),
    .S(_05068_),
    .X(_05074_));
 sky130_fd_sc_hd__clkbuf_1 _17606_ (.A(_05074_),
    .X(_01234_));
 sky130_fd_sc_hd__mux2_1 _17607_ (.A0(_13263_),
    .A1(\rvcpu.dp.rf.reg_file_arr[28][5] ),
    .S(_05068_),
    .X(_05075_));
 sky130_fd_sc_hd__clkbuf_1 _17608_ (.A(_05075_),
    .X(_01233_));
 sky130_fd_sc_hd__mux2_1 _17609_ (.A0(_13266_),
    .A1(\rvcpu.dp.rf.reg_file_arr[28][4] ),
    .S(_05068_),
    .X(_05076_));
 sky130_fd_sc_hd__clkbuf_1 _17610_ (.A(_05076_),
    .X(_01232_));
 sky130_fd_sc_hd__mux2_1 _17611_ (.A0(_13269_),
    .A1(\rvcpu.dp.rf.reg_file_arr[28][3] ),
    .S(_05068_),
    .X(_05077_));
 sky130_fd_sc_hd__clkbuf_1 _17612_ (.A(_05077_),
    .X(_01231_));
 sky130_fd_sc_hd__mux2_1 _17613_ (.A0(_13272_),
    .A1(\rvcpu.dp.rf.reg_file_arr[28][2] ),
    .S(_05068_),
    .X(_05078_));
 sky130_fd_sc_hd__clkbuf_1 _17614_ (.A(_05078_),
    .X(_01230_));
 sky130_fd_sc_hd__mux2_1 _17615_ (.A0(_13275_),
    .A1(\rvcpu.dp.rf.reg_file_arr[28][1] ),
    .S(_05045_),
    .X(_05079_));
 sky130_fd_sc_hd__clkbuf_1 _17616_ (.A(_05079_),
    .X(_01229_));
 sky130_fd_sc_hd__mux2_1 _17617_ (.A0(_13278_),
    .A1(\rvcpu.dp.rf.reg_file_arr[28][0] ),
    .S(_05045_),
    .X(_05080_));
 sky130_fd_sc_hd__clkbuf_1 _17618_ (.A(_05080_),
    .X(_01228_));
 sky130_fd_sc_hd__nor2_2 _17619_ (.A(_14234_),
    .B(_14347_),
    .Y(_05081_));
 sky130_fd_sc_hd__buf_4 _17620_ (.A(_05081_),
    .X(_05082_));
 sky130_fd_sc_hd__mux2_1 _17621_ (.A0(\rvcpu.dp.rf.reg_file_arr[2][31] ),
    .A1(_13172_),
    .S(_05082_),
    .X(_05083_));
 sky130_fd_sc_hd__clkbuf_1 _17622_ (.A(_05083_),
    .X(_01227_));
 sky130_fd_sc_hd__mux2_1 _17623_ (.A0(\rvcpu.dp.rf.reg_file_arr[2][30] ),
    .A1(_13183_),
    .S(_05082_),
    .X(_05084_));
 sky130_fd_sc_hd__clkbuf_1 _17624_ (.A(_05084_),
    .X(_01226_));
 sky130_fd_sc_hd__mux2_1 _17625_ (.A0(\rvcpu.dp.rf.reg_file_arr[2][29] ),
    .A1(_13186_),
    .S(_05082_),
    .X(_05085_));
 sky130_fd_sc_hd__clkbuf_1 _17626_ (.A(_05085_),
    .X(_01225_));
 sky130_fd_sc_hd__mux2_1 _17627_ (.A0(\rvcpu.dp.rf.reg_file_arr[2][28] ),
    .A1(_13189_),
    .S(_05082_),
    .X(_05086_));
 sky130_fd_sc_hd__clkbuf_1 _17628_ (.A(_05086_),
    .X(_01224_));
 sky130_fd_sc_hd__mux2_1 _17629_ (.A0(\rvcpu.dp.rf.reg_file_arr[2][27] ),
    .A1(_13194_),
    .S(_05082_),
    .X(_05087_));
 sky130_fd_sc_hd__clkbuf_1 _17630_ (.A(_05087_),
    .X(_01223_));
 sky130_fd_sc_hd__mux2_1 _17631_ (.A0(\rvcpu.dp.rf.reg_file_arr[2][26] ),
    .A1(_13197_),
    .S(_05082_),
    .X(_05088_));
 sky130_fd_sc_hd__clkbuf_1 _17632_ (.A(_05088_),
    .X(_01222_));
 sky130_fd_sc_hd__mux2_1 _17633_ (.A0(\rvcpu.dp.rf.reg_file_arr[2][25] ),
    .A1(_13200_),
    .S(_05082_),
    .X(_05089_));
 sky130_fd_sc_hd__clkbuf_1 _17634_ (.A(_05089_),
    .X(_01221_));
 sky130_fd_sc_hd__mux2_1 _17635_ (.A0(\rvcpu.dp.rf.reg_file_arr[2][24] ),
    .A1(_13203_),
    .S(_05082_),
    .X(_05090_));
 sky130_fd_sc_hd__clkbuf_1 _17636_ (.A(_05090_),
    .X(_01220_));
 sky130_fd_sc_hd__mux2_1 _17637_ (.A0(\rvcpu.dp.rf.reg_file_arr[2][23] ),
    .A1(_13206_),
    .S(_05082_),
    .X(_05091_));
 sky130_fd_sc_hd__clkbuf_1 _17638_ (.A(_05091_),
    .X(_01219_));
 sky130_fd_sc_hd__mux2_1 _17639_ (.A0(\rvcpu.dp.rf.reg_file_arr[2][22] ),
    .A1(_13209_),
    .S(_05082_),
    .X(_05092_));
 sky130_fd_sc_hd__clkbuf_1 _17640_ (.A(_05092_),
    .X(_01218_));
 sky130_fd_sc_hd__buf_4 _17641_ (.A(_05081_),
    .X(_05093_));
 sky130_fd_sc_hd__mux2_1 _17642_ (.A0(\rvcpu.dp.rf.reg_file_arr[2][21] ),
    .A1(_13212_),
    .S(_05093_),
    .X(_05094_));
 sky130_fd_sc_hd__clkbuf_1 _17643_ (.A(_05094_),
    .X(_01217_));
 sky130_fd_sc_hd__mux2_1 _17644_ (.A0(\rvcpu.dp.rf.reg_file_arr[2][20] ),
    .A1(_13216_),
    .S(_05093_),
    .X(_05095_));
 sky130_fd_sc_hd__clkbuf_1 _17645_ (.A(_05095_),
    .X(_01216_));
 sky130_fd_sc_hd__mux2_1 _17646_ (.A0(\rvcpu.dp.rf.reg_file_arr[2][19] ),
    .A1(_13219_),
    .S(_05093_),
    .X(_05096_));
 sky130_fd_sc_hd__clkbuf_1 _17647_ (.A(_05096_),
    .X(_01215_));
 sky130_fd_sc_hd__mux2_1 _17648_ (.A0(\rvcpu.dp.rf.reg_file_arr[2][18] ),
    .A1(_13222_),
    .S(_05093_),
    .X(_05097_));
 sky130_fd_sc_hd__clkbuf_1 _17649_ (.A(_05097_),
    .X(_01214_));
 sky130_fd_sc_hd__mux2_1 _17650_ (.A0(\rvcpu.dp.rf.reg_file_arr[2][17] ),
    .A1(_13225_),
    .S(_05093_),
    .X(_05098_));
 sky130_fd_sc_hd__clkbuf_1 _17651_ (.A(_05098_),
    .X(_01213_));
 sky130_fd_sc_hd__mux2_1 _17652_ (.A0(\rvcpu.dp.rf.reg_file_arr[2][16] ),
    .A1(_13228_),
    .S(_05093_),
    .X(_05099_));
 sky130_fd_sc_hd__clkbuf_1 _17653_ (.A(_05099_),
    .X(_01212_));
 sky130_fd_sc_hd__mux2_1 _17654_ (.A0(\rvcpu.dp.rf.reg_file_arr[2][15] ),
    .A1(_13231_),
    .S(_05093_),
    .X(_05100_));
 sky130_fd_sc_hd__clkbuf_1 _17655_ (.A(_05100_),
    .X(_01211_));
 sky130_fd_sc_hd__mux2_1 _17656_ (.A0(\rvcpu.dp.rf.reg_file_arr[2][14] ),
    .A1(_13234_),
    .S(_05093_),
    .X(_05101_));
 sky130_fd_sc_hd__clkbuf_1 _17657_ (.A(_05101_),
    .X(_01210_));
 sky130_fd_sc_hd__mux2_1 _17658_ (.A0(\rvcpu.dp.rf.reg_file_arr[2][13] ),
    .A1(_13237_),
    .S(_05093_),
    .X(_05102_));
 sky130_fd_sc_hd__clkbuf_1 _17659_ (.A(_05102_),
    .X(_01209_));
 sky130_fd_sc_hd__mux2_1 _17660_ (.A0(\rvcpu.dp.rf.reg_file_arr[2][12] ),
    .A1(_13240_),
    .S(_05093_),
    .X(_05103_));
 sky130_fd_sc_hd__clkbuf_1 _17661_ (.A(_05103_),
    .X(_01208_));
 sky130_fd_sc_hd__clkbuf_4 _17662_ (.A(_05081_),
    .X(_05104_));
 sky130_fd_sc_hd__mux2_1 _17663_ (.A0(\rvcpu.dp.rf.reg_file_arr[2][11] ),
    .A1(_13243_),
    .S(_05104_),
    .X(_05105_));
 sky130_fd_sc_hd__clkbuf_1 _17664_ (.A(_05105_),
    .X(_01207_));
 sky130_fd_sc_hd__mux2_1 _17665_ (.A0(\rvcpu.dp.rf.reg_file_arr[2][10] ),
    .A1(_13247_),
    .S(_05104_),
    .X(_05106_));
 sky130_fd_sc_hd__clkbuf_1 _17666_ (.A(_05106_),
    .X(_01206_));
 sky130_fd_sc_hd__mux2_1 _17667_ (.A0(\rvcpu.dp.rf.reg_file_arr[2][9] ),
    .A1(_13250_),
    .S(_05104_),
    .X(_05107_));
 sky130_fd_sc_hd__clkbuf_1 _17668_ (.A(_05107_),
    .X(_01205_));
 sky130_fd_sc_hd__mux2_1 _17669_ (.A0(\rvcpu.dp.rf.reg_file_arr[2][8] ),
    .A1(_13253_),
    .S(_05104_),
    .X(_05108_));
 sky130_fd_sc_hd__clkbuf_1 _17670_ (.A(_05108_),
    .X(_01204_));
 sky130_fd_sc_hd__mux2_1 _17671_ (.A0(\rvcpu.dp.rf.reg_file_arr[2][7] ),
    .A1(_13256_),
    .S(_05104_),
    .X(_05109_));
 sky130_fd_sc_hd__clkbuf_1 _17672_ (.A(_05109_),
    .X(_01203_));
 sky130_fd_sc_hd__mux2_1 _17673_ (.A0(\rvcpu.dp.rf.reg_file_arr[2][6] ),
    .A1(_13259_),
    .S(_05104_),
    .X(_05110_));
 sky130_fd_sc_hd__clkbuf_1 _17674_ (.A(_05110_),
    .X(_01202_));
 sky130_fd_sc_hd__mux2_1 _17675_ (.A0(\rvcpu.dp.rf.reg_file_arr[2][5] ),
    .A1(_13262_),
    .S(_05104_),
    .X(_05111_));
 sky130_fd_sc_hd__clkbuf_1 _17676_ (.A(_05111_),
    .X(_01201_));
 sky130_fd_sc_hd__mux2_1 _17677_ (.A0(\rvcpu.dp.rf.reg_file_arr[2][4] ),
    .A1(_13265_),
    .S(_05104_),
    .X(_05112_));
 sky130_fd_sc_hd__clkbuf_1 _17678_ (.A(_05112_),
    .X(_01200_));
 sky130_fd_sc_hd__mux2_1 _17679_ (.A0(\rvcpu.dp.rf.reg_file_arr[2][3] ),
    .A1(_13268_),
    .S(_05104_),
    .X(_05113_));
 sky130_fd_sc_hd__clkbuf_1 _17680_ (.A(_05113_),
    .X(_01199_));
 sky130_fd_sc_hd__mux2_1 _17681_ (.A0(\rvcpu.dp.rf.reg_file_arr[2][2] ),
    .A1(_13271_),
    .S(_05104_),
    .X(_05114_));
 sky130_fd_sc_hd__clkbuf_1 _17682_ (.A(_05114_),
    .X(_01198_));
 sky130_fd_sc_hd__mux2_1 _17683_ (.A0(\rvcpu.dp.rf.reg_file_arr[2][1] ),
    .A1(_13274_),
    .S(_05081_),
    .X(_05115_));
 sky130_fd_sc_hd__clkbuf_1 _17684_ (.A(_05115_),
    .X(_01197_));
 sky130_fd_sc_hd__mux2_1 _17685_ (.A0(\rvcpu.dp.rf.reg_file_arr[2][0] ),
    .A1(_13277_),
    .S(_05081_),
    .X(_05116_));
 sky130_fd_sc_hd__clkbuf_1 _17686_ (.A(_05116_),
    .X(_01196_));
 sky130_fd_sc_hd__nand2_2 _17687_ (.A(_14129_),
    .B(_04538_),
    .Y(_05117_));
 sky130_fd_sc_hd__clkbuf_4 _17688_ (.A(_05117_),
    .X(_05118_));
 sky130_fd_sc_hd__mux2_1 _17689_ (.A0(_13173_),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][31] ),
    .S(_05118_),
    .X(_05119_));
 sky130_fd_sc_hd__clkbuf_1 _17690_ (.A(_05119_),
    .X(_01195_));
 sky130_fd_sc_hd__mux2_1 _17691_ (.A0(_13184_),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][30] ),
    .S(_05118_),
    .X(_05120_));
 sky130_fd_sc_hd__clkbuf_1 _17692_ (.A(_05120_),
    .X(_01194_));
 sky130_fd_sc_hd__mux2_1 _17693_ (.A0(_13187_),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][29] ),
    .S(_05118_),
    .X(_05121_));
 sky130_fd_sc_hd__clkbuf_1 _17694_ (.A(_05121_),
    .X(_01193_));
 sky130_fd_sc_hd__mux2_1 _17695_ (.A0(_13190_),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][28] ),
    .S(_05118_),
    .X(_05122_));
 sky130_fd_sc_hd__clkbuf_1 _17696_ (.A(_05122_),
    .X(_01192_));
 sky130_fd_sc_hd__mux2_1 _17697_ (.A0(_13195_),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][27] ),
    .S(_05118_),
    .X(_05123_));
 sky130_fd_sc_hd__clkbuf_1 _17698_ (.A(_05123_),
    .X(_01191_));
 sky130_fd_sc_hd__mux2_1 _17699_ (.A0(_13198_),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][26] ),
    .S(_05118_),
    .X(_05124_));
 sky130_fd_sc_hd__clkbuf_1 _17700_ (.A(_05124_),
    .X(_01190_));
 sky130_fd_sc_hd__mux2_1 _17701_ (.A0(_13201_),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][25] ),
    .S(_05118_),
    .X(_05125_));
 sky130_fd_sc_hd__clkbuf_1 _17702_ (.A(_05125_),
    .X(_01189_));
 sky130_fd_sc_hd__mux2_1 _17703_ (.A0(_13204_),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][24] ),
    .S(_05118_),
    .X(_05126_));
 sky130_fd_sc_hd__clkbuf_1 _17704_ (.A(_05126_),
    .X(_01188_));
 sky130_fd_sc_hd__mux2_1 _17705_ (.A0(_13207_),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][23] ),
    .S(_05118_),
    .X(_05127_));
 sky130_fd_sc_hd__clkbuf_1 _17706_ (.A(_05127_),
    .X(_01187_));
 sky130_fd_sc_hd__mux2_1 _17707_ (.A0(_13210_),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][22] ),
    .S(_05118_),
    .X(_05128_));
 sky130_fd_sc_hd__clkbuf_1 _17708_ (.A(_05128_),
    .X(_01186_));
 sky130_fd_sc_hd__clkbuf_4 _17709_ (.A(_05117_),
    .X(_05129_));
 sky130_fd_sc_hd__mux2_1 _17710_ (.A0(_13213_),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][21] ),
    .S(_05129_),
    .X(_05130_));
 sky130_fd_sc_hd__clkbuf_1 _17711_ (.A(_05130_),
    .X(_01185_));
 sky130_fd_sc_hd__mux2_1 _17712_ (.A0(_13217_),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][20] ),
    .S(_05129_),
    .X(_05131_));
 sky130_fd_sc_hd__clkbuf_1 _17713_ (.A(_05131_),
    .X(_01184_));
 sky130_fd_sc_hd__mux2_1 _17714_ (.A0(_13220_),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][19] ),
    .S(_05129_),
    .X(_05132_));
 sky130_fd_sc_hd__clkbuf_1 _17715_ (.A(_05132_),
    .X(_01183_));
 sky130_fd_sc_hd__mux2_1 _17716_ (.A0(_13223_),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][18] ),
    .S(_05129_),
    .X(_05133_));
 sky130_fd_sc_hd__clkbuf_1 _17717_ (.A(_05133_),
    .X(_01182_));
 sky130_fd_sc_hd__mux2_1 _17718_ (.A0(_13226_),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][17] ),
    .S(_05129_),
    .X(_05134_));
 sky130_fd_sc_hd__clkbuf_1 _17719_ (.A(_05134_),
    .X(_01181_));
 sky130_fd_sc_hd__mux2_1 _17720_ (.A0(_13229_),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][16] ),
    .S(_05129_),
    .X(_05135_));
 sky130_fd_sc_hd__clkbuf_1 _17721_ (.A(_05135_),
    .X(_01180_));
 sky130_fd_sc_hd__mux2_1 _17722_ (.A0(_13232_),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][15] ),
    .S(_05129_),
    .X(_05136_));
 sky130_fd_sc_hd__clkbuf_1 _17723_ (.A(_05136_),
    .X(_01179_));
 sky130_fd_sc_hd__mux2_1 _17724_ (.A0(_13235_),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][14] ),
    .S(_05129_),
    .X(_05137_));
 sky130_fd_sc_hd__clkbuf_1 _17725_ (.A(_05137_),
    .X(_01178_));
 sky130_fd_sc_hd__mux2_1 _17726_ (.A0(_13238_),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][13] ),
    .S(_05129_),
    .X(_05138_));
 sky130_fd_sc_hd__clkbuf_1 _17727_ (.A(_05138_),
    .X(_01177_));
 sky130_fd_sc_hd__mux2_1 _17728_ (.A0(_13241_),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][12] ),
    .S(_05129_),
    .X(_05139_));
 sky130_fd_sc_hd__clkbuf_1 _17729_ (.A(_05139_),
    .X(_01176_));
 sky130_fd_sc_hd__buf_4 _17730_ (.A(_05117_),
    .X(_05140_));
 sky130_fd_sc_hd__mux2_1 _17731_ (.A0(_13244_),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][11] ),
    .S(_05140_),
    .X(_05141_));
 sky130_fd_sc_hd__clkbuf_1 _17732_ (.A(_05141_),
    .X(_01175_));
 sky130_fd_sc_hd__mux2_1 _17733_ (.A0(_13248_),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][10] ),
    .S(_05140_),
    .X(_05142_));
 sky130_fd_sc_hd__clkbuf_1 _17734_ (.A(_05142_),
    .X(_01174_));
 sky130_fd_sc_hd__mux2_1 _17735_ (.A0(_13251_),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][9] ),
    .S(_05140_),
    .X(_05143_));
 sky130_fd_sc_hd__clkbuf_1 _17736_ (.A(_05143_),
    .X(_01173_));
 sky130_fd_sc_hd__mux2_1 _17737_ (.A0(_13254_),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][8] ),
    .S(_05140_),
    .X(_05144_));
 sky130_fd_sc_hd__clkbuf_1 _17738_ (.A(_05144_),
    .X(_01172_));
 sky130_fd_sc_hd__mux2_1 _17739_ (.A0(_13257_),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][7] ),
    .S(_05140_),
    .X(_05145_));
 sky130_fd_sc_hd__clkbuf_1 _17740_ (.A(_05145_),
    .X(_01171_));
 sky130_fd_sc_hd__mux2_1 _17741_ (.A0(_13260_),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][6] ),
    .S(_05140_),
    .X(_05146_));
 sky130_fd_sc_hd__clkbuf_1 _17742_ (.A(_05146_),
    .X(_01170_));
 sky130_fd_sc_hd__mux2_1 _17743_ (.A0(_13263_),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][5] ),
    .S(_05140_),
    .X(_05147_));
 sky130_fd_sc_hd__clkbuf_1 _17744_ (.A(_05147_),
    .X(_01169_));
 sky130_fd_sc_hd__mux2_1 _17745_ (.A0(_13266_),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][4] ),
    .S(_05140_),
    .X(_05148_));
 sky130_fd_sc_hd__clkbuf_1 _17746_ (.A(_05148_),
    .X(_01168_));
 sky130_fd_sc_hd__mux2_1 _17747_ (.A0(_13269_),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][3] ),
    .S(_05140_),
    .X(_05149_));
 sky130_fd_sc_hd__clkbuf_1 _17748_ (.A(_05149_),
    .X(_01167_));
 sky130_fd_sc_hd__mux2_1 _17749_ (.A0(_13272_),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][2] ),
    .S(_05140_),
    .X(_05150_));
 sky130_fd_sc_hd__clkbuf_1 _17750_ (.A(_05150_),
    .X(_01166_));
 sky130_fd_sc_hd__mux2_1 _17751_ (.A0(_13275_),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][1] ),
    .S(_05117_),
    .X(_05151_));
 sky130_fd_sc_hd__clkbuf_1 _17752_ (.A(_05151_),
    .X(_01165_));
 sky130_fd_sc_hd__mux2_1 _17753_ (.A0(_13278_),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][0] ),
    .S(_05117_),
    .X(_05152_));
 sky130_fd_sc_hd__clkbuf_1 _17754_ (.A(_05152_),
    .X(_01164_));
 sky130_fd_sc_hd__xnor2_1 _17755_ (.A(_13176_),
    .B(\rvcpu.dp.plde.Rs2E[4] ),
    .Y(_05153_));
 sky130_fd_sc_hd__o21a_2 _17756_ (.A1(_13175_),
    .A2(\rvcpu.dp.plde.Rs2E[3] ),
    .B1(_05153_),
    .X(_05154_));
 sky130_fd_sc_hd__xor2_1 _17757_ (.A(\rvcpu.dp.plmw.RdW[1] ),
    .B(\rvcpu.dp.plde.Rs2E[1] ),
    .X(_05155_));
 sky130_fd_sc_hd__a221o_1 _17758_ (.A1(_14346_),
    .A2(\rvcpu.dp.plde.Rs2E[0] ),
    .B1(\rvcpu.dp.plde.Rs2E[3] ),
    .B2(_13175_),
    .C1(_05155_),
    .X(_05156_));
 sky130_fd_sc_hd__or4_1 _17759_ (.A(\rvcpu.dp.plde.Rs2E[1] ),
    .B(\rvcpu.dp.plde.Rs2E[0] ),
    .C(\rvcpu.dp.plde.Rs2E[2] ),
    .D(\rvcpu.dp.plde.Rs2E[4] ),
    .X(_05157_));
 sky130_fd_sc_hd__nor2_1 _17760_ (.A(\rvcpu.dp.plde.Rs2E[3] ),
    .B(_05157_),
    .Y(_05158_));
 sky130_fd_sc_hd__xnor2_1 _17761_ (.A(_13174_),
    .B(\rvcpu.dp.plde.Rs2E[2] ),
    .Y(_05159_));
 sky130_fd_sc_hd__o21a_1 _17762_ (.A1(_14346_),
    .A2(\rvcpu.dp.plde.Rs2E[0] ),
    .B1(\rvcpu.dp.plmw.RegWriteW ),
    .X(_05160_));
 sky130_fd_sc_hd__and4bb_4 _17763_ (.A_N(_05156_),
    .B_N(_05158_),
    .C(_05159_),
    .D(_05160_),
    .X(_05161_));
 sky130_fd_sc_hd__inv_2 _17764_ (.A(\rvcpu.dp.plem.RdM[0] ),
    .Y(_05162_));
 sky130_fd_sc_hd__xnor2_1 _17765_ (.A(\rvcpu.dp.plem.RdM[4] ),
    .B(\rvcpu.dp.plde.Rs2E[4] ),
    .Y(_05163_));
 sky130_fd_sc_hd__o21ai_1 _17766_ (.A1(_05162_),
    .A2(\rvcpu.dp.plde.Rs2E[0] ),
    .B1(_05163_),
    .Y(_05164_));
 sky130_fd_sc_hd__inv_2 _17767_ (.A(\rvcpu.dp.plde.Rs2E[1] ),
    .Y(_05165_));
 sky130_fd_sc_hd__xor2_1 _17768_ (.A(\rvcpu.dp.plem.RdM[2] ),
    .B(\rvcpu.dp.plde.Rs2E[2] ),
    .X(_05166_));
 sky130_fd_sc_hd__a221o_1 _17769_ (.A1(\rvcpu.dp.plem.RdM[1] ),
    .A2(_05165_),
    .B1(\rvcpu.dp.plde.Rs2E[0] ),
    .B2(_05162_),
    .C1(_05166_),
    .X(_05167_));
 sky130_fd_sc_hd__and2_1 _17770_ (.A(\rvcpu.dp.plem.RdM[3] ),
    .B(\rvcpu.dp.plde.Rs2E[3] ),
    .X(_05168_));
 sky130_fd_sc_hd__nor2_1 _17771_ (.A(\rvcpu.dp.plem.RdM[3] ),
    .B(\rvcpu.dp.plde.Rs2E[3] ),
    .Y(_05169_));
 sky130_fd_sc_hd__o221a_1 _17772_ (.A1(\rvcpu.dp.plem.RdM[1] ),
    .A2(_05165_),
    .B1(_05168_),
    .B2(_05169_),
    .C1(\rvcpu.dp.plem.RegWriteM ),
    .X(_05170_));
 sky130_fd_sc_hd__nor4b_1 _17773_ (.A(_05158_),
    .B(_05164_),
    .C(_05167_),
    .D_N(_05170_),
    .Y(_05171_));
 sky130_fd_sc_hd__a31oi_1 _17774_ (.A1(_13277_),
    .A2(_05154_),
    .A3(_05161_),
    .B1(net115),
    .Y(_05172_));
 sky130_fd_sc_hd__a21bo_1 _17775_ (.A1(_05154_),
    .A2(_05161_),
    .B1_N(\rvcpu.dp.plde.RD2E[0] ),
    .X(_05173_));
 sky130_fd_sc_hd__or4b_2 _17776_ (.A(_05158_),
    .B(_05164_),
    .C(_05167_),
    .D_N(_05170_),
    .X(_05174_));
 sky130_fd_sc_hd__clkbuf_4 _17777_ (.A(_05174_),
    .X(_05175_));
 sky130_fd_sc_hd__clkbuf_4 _17778_ (.A(_05175_),
    .X(_05176_));
 sky130_fd_sc_hd__clkbuf_4 _17779_ (.A(_05176_),
    .X(_05177_));
 sky130_fd_sc_hd__clkbuf_4 _17780_ (.A(_05177_),
    .X(_05178_));
 sky130_fd_sc_hd__o2bb2a_1 _17781_ (.A1_N(_05172_),
    .A2_N(_05173_),
    .B1(_05178_),
    .B2(\rvcpu.dp.plem.ALUResultM[0] ),
    .X(\rvcpu.dp.SrcBFW_Mux.y[0] ));
 sky130_fd_sc_hd__buf_2 _17782_ (.A(_05154_),
    .X(_05179_));
 sky130_fd_sc_hd__buf_2 _17783_ (.A(_05161_),
    .X(_05180_));
 sky130_fd_sc_hd__a21boi_2 _17784_ (.A1(_05179_),
    .A2(_05180_),
    .B1_N(\rvcpu.dp.plde.RD2E[1] ),
    .Y(_05181_));
 sky130_fd_sc_hd__a31o_1 _17785_ (.A1(_13274_),
    .A2(_05154_),
    .A3(_05161_),
    .B1(net114),
    .X(_05182_));
 sky130_fd_sc_hd__o22a_1 _17786_ (.A1(\rvcpu.dp.plem.ALUResultM[1] ),
    .A2(_05178_),
    .B1(_05181_),
    .B2(_05182_),
    .X(\rvcpu.dp.SrcBFW_Mux.y[1] ));
 sky130_fd_sc_hd__nand3b_1 _17787_ (.A_N(_13271_),
    .B(_05179_),
    .C(_05180_),
    .Y(_05183_));
 sky130_fd_sc_hd__a21o_1 _17788_ (.A1(_05154_),
    .A2(_05161_),
    .B1(\rvcpu.dp.plde.RD2E[2] ),
    .X(_05184_));
 sky130_fd_sc_hd__inv_2 _17789_ (.A(net122),
    .Y(_05185_));
 sky130_fd_sc_hd__nor2_1 _17790_ (.A(_05185_),
    .B(_05175_),
    .Y(_05186_));
 sky130_fd_sc_hd__a31o_1 _17791_ (.A1(_05175_),
    .A2(_05183_),
    .A3(_05184_),
    .B1(_05186_),
    .X(_05187_));
 sky130_fd_sc_hd__buf_1 _17792_ (.A(_05187_),
    .X(\rvcpu.dp.SrcBFW_Mux.y[2] ));
 sky130_fd_sc_hd__a21boi_1 _17793_ (.A1(_05179_),
    .A2(_05180_),
    .B1_N(\rvcpu.dp.plde.RD2E[3] ),
    .Y(_05188_));
 sky130_fd_sc_hd__a31o_1 _17794_ (.A1(_13268_),
    .A2(_05154_),
    .A3(_05161_),
    .B1(net114),
    .X(_05189_));
 sky130_fd_sc_hd__o22a_1 _17795_ (.A1(\rvcpu.dp.plem.ALUResultM[3] ),
    .A2(_05175_),
    .B1(_05188_),
    .B2(_05189_),
    .X(_05190_));
 sky130_fd_sc_hd__buf_1 _17796_ (.A(_05190_),
    .X(\rvcpu.dp.SrcBFW_Mux.y[3] ));
 sky130_fd_sc_hd__a21boi_1 _17797_ (.A1(_05179_),
    .A2(_05180_),
    .B1_N(\rvcpu.dp.plde.RD2E[4] ),
    .Y(_05191_));
 sky130_fd_sc_hd__a31o_1 _17798_ (.A1(_13265_),
    .A2(_05179_),
    .A3(_05180_),
    .B1(net114),
    .X(_05192_));
 sky130_fd_sc_hd__o22a_1 _17799_ (.A1(\rvcpu.dp.plem.ALUResultM[4] ),
    .A2(_05175_),
    .B1(_05191_),
    .B2(_05192_),
    .X(_05193_));
 sky130_fd_sc_hd__clkbuf_2 _17800_ (.A(_05193_),
    .X(\rvcpu.dp.SrcBFW_Mux.y[4] ));
 sky130_fd_sc_hd__nand2_2 _17801_ (.A(_05154_),
    .B(_05161_),
    .Y(_05194_));
 sky130_fd_sc_hd__clkbuf_4 _17802_ (.A(_05194_),
    .X(_05195_));
 sky130_fd_sc_hd__clkbuf_4 _17803_ (.A(_05195_),
    .X(_05196_));
 sky130_fd_sc_hd__mux2_1 _17804_ (.A0(_13172_),
    .A1(\rvcpu.dp.plde.RD2E[31] ),
    .S(_05196_),
    .X(_05197_));
 sky130_fd_sc_hd__mux2_1 _17805_ (.A0(\rvcpu.dp.plem.ALUResultM[31] ),
    .A1(_05197_),
    .S(_05178_),
    .X(_05198_));
 sky130_fd_sc_hd__clkbuf_2 _17806_ (.A(_05198_),
    .X(\rvcpu.dp.SrcBFW_Mux.y[31] ));
 sky130_fd_sc_hd__mux2_1 _17807_ (.A0(_13183_),
    .A1(\rvcpu.dp.plde.RD2E[30] ),
    .S(_05196_),
    .X(_05199_));
 sky130_fd_sc_hd__mux2_1 _17808_ (.A0(\rvcpu.dp.plem.ALUResultM[30] ),
    .A1(_05199_),
    .S(_05178_),
    .X(_05200_));
 sky130_fd_sc_hd__clkbuf_2 _17809_ (.A(_05200_),
    .X(\rvcpu.dp.SrcBFW_Mux.y[30] ));
 sky130_fd_sc_hd__mux2_1 _17810_ (.A0(_13186_),
    .A1(\rvcpu.dp.plde.RD2E[29] ),
    .S(_05196_),
    .X(_05201_));
 sky130_fd_sc_hd__mux2_1 _17811_ (.A0(\rvcpu.dp.plem.ALUResultM[29] ),
    .A1(_05201_),
    .S(_05178_),
    .X(_05202_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17812_ (.A(_05202_),
    .X(\rvcpu.dp.SrcBFW_Mux.y[29] ));
 sky130_fd_sc_hd__mux2_1 _17813_ (.A0(_13189_),
    .A1(\rvcpu.dp.plde.RD2E[28] ),
    .S(_05196_),
    .X(_05203_));
 sky130_fd_sc_hd__mux2_1 _17814_ (.A0(\rvcpu.dp.plem.ALUResultM[28] ),
    .A1(_05203_),
    .S(_05178_),
    .X(_05204_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17815_ (.A(_05204_),
    .X(\rvcpu.dp.SrcBFW_Mux.y[28] ));
 sky130_fd_sc_hd__mux2_1 _17816_ (.A0(_13194_),
    .A1(\rvcpu.dp.plde.RD2E[27] ),
    .S(_05196_),
    .X(_05205_));
 sky130_fd_sc_hd__mux2_1 _17817_ (.A0(\rvcpu.dp.plem.ALUResultM[27] ),
    .A1(_05205_),
    .S(_05178_),
    .X(_05206_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17818_ (.A(_05206_),
    .X(\rvcpu.dp.SrcBFW_Mux.y[27] ));
 sky130_fd_sc_hd__mux2_1 _17819_ (.A0(_13197_),
    .A1(\rvcpu.dp.plde.RD2E[26] ),
    .S(_05196_),
    .X(_05207_));
 sky130_fd_sc_hd__mux2_1 _17820_ (.A0(\rvcpu.dp.plem.ALUResultM[26] ),
    .A1(_05207_),
    .S(_05178_),
    .X(_05208_));
 sky130_fd_sc_hd__buf_1 _17821_ (.A(_05208_),
    .X(\rvcpu.dp.SrcBFW_Mux.y[26] ));
 sky130_fd_sc_hd__mux2_1 _17822_ (.A0(_13200_),
    .A1(\rvcpu.dp.plde.RD2E[25] ),
    .S(_05196_),
    .X(_05209_));
 sky130_fd_sc_hd__mux2_1 _17823_ (.A0(\rvcpu.dp.plem.ALUResultM[25] ),
    .A1(_05209_),
    .S(_05178_),
    .X(_05210_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17824_ (.A(_05210_),
    .X(\rvcpu.dp.SrcBFW_Mux.y[25] ));
 sky130_fd_sc_hd__mux2_1 _17825_ (.A0(_13203_),
    .A1(\rvcpu.dp.plde.RD2E[24] ),
    .S(_05196_),
    .X(_05211_));
 sky130_fd_sc_hd__mux2_1 _17826_ (.A0(\rvcpu.dp.plem.ALUResultM[24] ),
    .A1(_05211_),
    .S(_05178_),
    .X(_05212_));
 sky130_fd_sc_hd__clkbuf_2 _17827_ (.A(_05212_),
    .X(\rvcpu.dp.SrcBFW_Mux.y[24] ));
 sky130_fd_sc_hd__mux2_1 _17828_ (.A0(_13206_),
    .A1(\rvcpu.dp.plde.RD2E[23] ),
    .S(_05195_),
    .X(_05213_));
 sky130_fd_sc_hd__mux2_1 _17829_ (.A0(\rvcpu.dp.plem.ALUResultM[23] ),
    .A1(_05213_),
    .S(_05177_),
    .X(_05214_));
 sky130_fd_sc_hd__clkbuf_2 _17830_ (.A(_05214_),
    .X(\rvcpu.dp.SrcBFW_Mux.y[23] ));
 sky130_fd_sc_hd__mux2_1 _17831_ (.A0(_13209_),
    .A1(\rvcpu.dp.plde.RD2E[22] ),
    .S(_05196_),
    .X(_05215_));
 sky130_fd_sc_hd__mux2_1 _17832_ (.A0(\rvcpu.dp.plem.ALUResultM[22] ),
    .A1(_05215_),
    .S(_05177_),
    .X(_05216_));
 sky130_fd_sc_hd__clkbuf_2 _17833_ (.A(_05216_),
    .X(\rvcpu.dp.SrcBFW_Mux.y[22] ));
 sky130_fd_sc_hd__mux2_1 _17834_ (.A0(_13212_),
    .A1(\rvcpu.dp.plde.RD2E[21] ),
    .S(_05195_),
    .X(_05217_));
 sky130_fd_sc_hd__mux2_1 _17835_ (.A0(\rvcpu.dp.plem.ALUResultM[21] ),
    .A1(_05217_),
    .S(_05177_),
    .X(_05218_));
 sky130_fd_sc_hd__clkbuf_2 _17836_ (.A(_05218_),
    .X(\rvcpu.dp.SrcBFW_Mux.y[21] ));
 sky130_fd_sc_hd__mux2_1 _17837_ (.A0(_13219_),
    .A1(\rvcpu.dp.plde.RD2E[19] ),
    .S(_05195_),
    .X(_05219_));
 sky130_fd_sc_hd__mux2_1 _17838_ (.A0(\rvcpu.dp.plem.ALUResultM[19] ),
    .A1(_05219_),
    .S(_05177_),
    .X(_05220_));
 sky130_fd_sc_hd__clkbuf_2 _17839_ (.A(_05220_),
    .X(\rvcpu.dp.SrcBFW_Mux.y[19] ));
 sky130_fd_sc_hd__mux2_1 _17840_ (.A0(_13225_),
    .A1(\rvcpu.dp.plde.RD2E[17] ),
    .S(_05195_),
    .X(_05221_));
 sky130_fd_sc_hd__mux2_1 _17841_ (.A0(\rvcpu.dp.plem.ALUResultM[17] ),
    .A1(_05221_),
    .S(_05177_),
    .X(_05222_));
 sky130_fd_sc_hd__buf_1 _17842_ (.A(_05222_),
    .X(\rvcpu.dp.SrcBFW_Mux.y[17] ));
 sky130_fd_sc_hd__mux2_1 _17843_ (.A0(_13231_),
    .A1(\rvcpu.dp.plde.RD2E[15] ),
    .S(_05194_),
    .X(_05223_));
 sky130_fd_sc_hd__mux2_1 _17844_ (.A0(\rvcpu.dp.plem.ALUResultM[15] ),
    .A1(_05223_),
    .S(_05175_),
    .X(_05224_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17845_ (.A(_05224_),
    .X(\rvcpu.dp.SrcBFW_Mux.y[15] ));
 sky130_fd_sc_hd__a31o_1 _17846_ (.A1(_13237_),
    .A2(_05179_),
    .A3(_05180_),
    .B1(net114),
    .X(_05225_));
 sky130_fd_sc_hd__a21oi_2 _17847_ (.A1(\rvcpu.dp.plde.RD2E[13] ),
    .A2(_05195_),
    .B1(_05225_),
    .Y(_05226_));
 sky130_fd_sc_hd__nor2_1 _17848_ (.A(\rvcpu.dp.plem.ALUResultM[13] ),
    .B(_05177_),
    .Y(_05227_));
 sky130_fd_sc_hd__nor2_1 _17849_ (.A(_05226_),
    .B(_05227_),
    .Y(\rvcpu.dp.SrcBFW_Mux.y[13] ));
 sky130_fd_sc_hd__mux2_1 _17850_ (.A0(_13243_),
    .A1(\rvcpu.dp.plde.RD2E[11] ),
    .S(_05194_),
    .X(_05228_));
 sky130_fd_sc_hd__mux2_1 _17851_ (.A0(\rvcpu.dp.plem.ALUResultM[11] ),
    .A1(_05228_),
    .S(_05176_),
    .X(_05229_));
 sky130_fd_sc_hd__buf_1 _17852_ (.A(_05229_),
    .X(\rvcpu.dp.SrcBFW_Mux.y[11] ));
 sky130_fd_sc_hd__mux2_1 _17853_ (.A0(_13250_),
    .A1(\rvcpu.dp.plde.RD2E[9] ),
    .S(_05194_),
    .X(_05230_));
 sky130_fd_sc_hd__mux2_1 _17854_ (.A0(\rvcpu.dp.plem.ALUResultM[9] ),
    .A1(_05230_),
    .S(_05176_),
    .X(_05231_));
 sky130_fd_sc_hd__buf_1 _17855_ (.A(_05231_),
    .X(\rvcpu.dp.SrcBFW_Mux.y[9] ));
 sky130_fd_sc_hd__mux2_1 _17856_ (.A0(_13256_),
    .A1(\rvcpu.dp.plde.RD2E[7] ),
    .S(_05195_),
    .X(_05232_));
 sky130_fd_sc_hd__mux2_1 _17857_ (.A0(\rvcpu.dp.plem.ALUResultM[7] ),
    .A1(_05232_),
    .S(_05176_),
    .X(_05233_));
 sky130_fd_sc_hd__buf_1 _17858_ (.A(_05233_),
    .X(\rvcpu.dp.SrcBFW_Mux.y[7] ));
 sky130_fd_sc_hd__a21boi_1 _17859_ (.A1(_05179_),
    .A2(_05180_),
    .B1_N(\rvcpu.dp.plde.RD2E[5] ),
    .Y(_05234_));
 sky130_fd_sc_hd__a31o_1 _17860_ (.A1(_13262_),
    .A2(_05179_),
    .A3(_05180_),
    .B1(net114),
    .X(_05235_));
 sky130_fd_sc_hd__o22a_1 _17861_ (.A1(\rvcpu.dp.plem.ALUResultM[5] ),
    .A2(_05176_),
    .B1(_05234_),
    .B2(_05235_),
    .X(\rvcpu.dp.SrcBFW_Mux.y[5] ));
 sky130_fd_sc_hd__or2_1 _17862_ (.A(\rvcpu.dp.plde.ALUControlE[3] ),
    .B(\rvcpu.dp.plde.ALUControlE[2] ),
    .X(_05236_));
 sky130_fd_sc_hd__or2_1 _17863_ (.A(\rvcpu.dp.plde.ALUControlE[1] ),
    .B(_05236_),
    .X(_05237_));
 sky130_fd_sc_hd__buf_2 _17864_ (.A(_05237_),
    .X(_00003_));
 sky130_fd_sc_hd__nor2_1 _17865_ (.A(\rvcpu.dp.plde.ALUControlE[0] ),
    .B(_00003_),
    .Y(_05238_));
 sky130_fd_sc_hd__clkbuf_4 _17866_ (.A(_05238_),
    .X(_05239_));
 sky130_fd_sc_hd__clkbuf_4 _17867_ (.A(_05239_),
    .X(_05240_));
 sky130_fd_sc_hd__inv_2 _17868_ (.A(\rvcpu.dp.plde.Rs1E[0] ),
    .Y(_05241_));
 sky130_fd_sc_hd__or4_1 _17869_ (.A(\rvcpu.dp.plde.Rs1E[1] ),
    .B(\rvcpu.dp.plde.Rs1E[0] ),
    .C(\rvcpu.dp.plde.Rs1E[2] ),
    .D(\rvcpu.dp.plde.Rs1E[4] ),
    .X(_05242_));
 sky130_fd_sc_hd__xnor2_1 _17870_ (.A(\rvcpu.dp.plde.Rs1E[4] ),
    .B(\rvcpu.dp.plem.RdM[4] ),
    .Y(_05243_));
 sky130_fd_sc_hd__o221a_1 _17871_ (.A1(_05241_),
    .A2(\rvcpu.dp.plem.RdM[0] ),
    .B1(_05242_),
    .B2(\rvcpu.dp.plde.Rs1E[3] ),
    .C1(_05243_),
    .X(_05244_));
 sky130_fd_sc_hd__inv_2 _17872_ (.A(\rvcpu.dp.plem.RdM[3] ),
    .Y(_05245_));
 sky130_fd_sc_hd__xnor2_1 _17873_ (.A(\rvcpu.dp.plde.Rs1E[2] ),
    .B(\rvcpu.dp.plem.RdM[2] ),
    .Y(_05246_));
 sky130_fd_sc_hd__o221a_1 _17874_ (.A1(\rvcpu.dp.plde.Rs1E[0] ),
    .A2(_05162_),
    .B1(_05245_),
    .B2(\rvcpu.dp.plde.Rs1E[3] ),
    .C1(_05246_),
    .X(_05247_));
 sky130_fd_sc_hd__inv_2 _17875_ (.A(\rvcpu.dp.plde.Rs1E[3] ),
    .Y(_05248_));
 sky130_fd_sc_hd__and2_1 _17876_ (.A(\rvcpu.dp.plde.Rs1E[1] ),
    .B(\rvcpu.dp.plem.RdM[1] ),
    .X(_05249_));
 sky130_fd_sc_hd__nor2_1 _17877_ (.A(\rvcpu.dp.plde.Rs1E[1] ),
    .B(\rvcpu.dp.plem.RdM[1] ),
    .Y(_05250_));
 sky130_fd_sc_hd__o221a_1 _17878_ (.A1(_05248_),
    .A2(\rvcpu.dp.plem.RdM[3] ),
    .B1(_05249_),
    .B2(_05250_),
    .C1(\rvcpu.dp.plem.RegWriteM ),
    .X(_05251_));
 sky130_fd_sc_hd__nand3_2 _17879_ (.A(_05244_),
    .B(_05247_),
    .C(_05251_),
    .Y(_05252_));
 sky130_fd_sc_hd__xor2_1 _17880_ (.A(\rvcpu.dp.plde.Rs1E[3] ),
    .B(\rvcpu.dp.plmw.RdW[3] ),
    .X(_05253_));
 sky130_fd_sc_hd__or2b_1 _17881_ (.A(\rvcpu.dp.plde.Rs1E[0] ),
    .B_N(\rvcpu.dp.plmw.RegWriteW ),
    .X(_05254_));
 sky130_fd_sc_hd__and2b_1 _17882_ (.A_N(\rvcpu.dp.plmw.RdW[4] ),
    .B(\rvcpu.dp.plde.Rs1E[4] ),
    .X(_05255_));
 sky130_fd_sc_hd__xor2_1 _17883_ (.A(\rvcpu.dp.plde.Rs1E[1] ),
    .B(\rvcpu.dp.plmw.RdW[1] ),
    .X(_05256_));
 sky130_fd_sc_hd__and2b_1 _17884_ (.A_N(\rvcpu.dp.plde.Rs1E[2] ),
    .B(_13174_),
    .X(_05257_));
 sky130_fd_sc_hd__a2111o_1 _17885_ (.A1(_13178_),
    .A2(_05254_),
    .B1(_05255_),
    .C1(_05256_),
    .D1(_05257_),
    .X(_05258_));
 sky130_fd_sc_hd__or2b_1 _17886_ (.A(\rvcpu.dp.plmw.RdW[2] ),
    .B_N(\rvcpu.dp.plde.Rs1E[2] ),
    .X(_05259_));
 sky130_fd_sc_hd__or2b_1 _17887_ (.A(\rvcpu.dp.plde.Rs1E[4] ),
    .B_N(_13176_),
    .X(_05260_));
 sky130_fd_sc_hd__or2b_1 _17888_ (.A(\rvcpu.dp.plde.Rs1E[0] ),
    .B_N(\rvcpu.dp.plmw.RdW[0] ),
    .X(_05261_));
 sky130_fd_sc_hd__o2111a_1 _17889_ (.A1(\rvcpu.dp.plde.Rs1E[3] ),
    .A2(_05242_),
    .B1(_05259_),
    .C1(_05260_),
    .D1(_05261_),
    .X(_05262_));
 sky130_fd_sc_hd__or3b_4 _17890_ (.A(_05253_),
    .B(_05258_),
    .C_N(_05262_),
    .X(_05263_));
 sky130_fd_sc_hd__and2_1 _17891_ (.A(_05252_),
    .B(_05263_),
    .X(_05264_));
 sky130_fd_sc_hd__clkbuf_4 _17892_ (.A(_05264_),
    .X(_05265_));
 sky130_fd_sc_hd__buf_4 _17893_ (.A(_05265_),
    .X(_05266_));
 sky130_fd_sc_hd__buf_4 _17894_ (.A(_05266_),
    .X(_05267_));
 sky130_fd_sc_hd__and3_4 _17895_ (.A(_05244_),
    .B(_05247_),
    .C(_05251_),
    .X(_05268_));
 sky130_fd_sc_hd__nor2_4 _17896_ (.A(_05268_),
    .B(_05263_),
    .Y(_05269_));
 sky130_fd_sc_hd__clkbuf_4 _17897_ (.A(_05269_),
    .X(_05270_));
 sky130_fd_sc_hd__buf_4 _17898_ (.A(_05270_),
    .X(_05271_));
 sky130_fd_sc_hd__buf_2 _17899_ (.A(_05268_),
    .X(_05272_));
 sky130_fd_sc_hd__and2_1 _17900_ (.A(\rvcpu.dp.plem.ALUResultM[31] ),
    .B(_05272_),
    .X(_05273_));
 sky130_fd_sc_hd__a221o_1 _17901_ (.A1(\rvcpu.dp.plde.RD1E[31] ),
    .A2(_05267_),
    .B1(_05271_),
    .B2(_13172_),
    .C1(_05273_),
    .X(_05274_));
 sky130_fd_sc_hd__buf_2 _17902_ (.A(_05274_),
    .X(_05275_));
 sky130_fd_sc_hd__inv_2 _17903_ (.A(\rvcpu.dp.plde.ALUSrcE ),
    .Y(_05276_));
 sky130_fd_sc_hd__clkbuf_4 _17904_ (.A(_05276_),
    .X(_05277_));
 sky130_fd_sc_hd__clkbuf_4 _17905_ (.A(_05277_),
    .X(_05278_));
 sky130_fd_sc_hd__clkbuf_4 _17906_ (.A(_05278_),
    .X(_05279_));
 sky130_fd_sc_hd__mux2_1 _17907_ (.A0(\rvcpu.dp.plde.ImmExtE[31] ),
    .A1(\rvcpu.dp.SrcBFW_Mux.y[31] ),
    .S(_05279_),
    .X(_05280_));
 sky130_fd_sc_hd__or2_1 _17908_ (.A(_05275_),
    .B(_05280_),
    .X(_05281_));
 sky130_fd_sc_hd__nand2_1 _17909_ (.A(_05275_),
    .B(_05280_),
    .Y(_05282_));
 sky130_fd_sc_hd__and2_1 _17910_ (.A(_05281_),
    .B(_05282_),
    .X(_05283_));
 sky130_fd_sc_hd__inv_2 _17911_ (.A(_05283_),
    .Y(_05284_));
 sky130_fd_sc_hd__and2_1 _17912_ (.A(\rvcpu.dp.plem.ALUResultM[30] ),
    .B(_05268_),
    .X(_05285_));
 sky130_fd_sc_hd__a221o_2 _17913_ (.A1(\rvcpu.dp.plde.RD1E[30] ),
    .A2(_05265_),
    .B1(_05269_),
    .B2(_13183_),
    .C1(_05285_),
    .X(_05286_));
 sky130_fd_sc_hd__mux2_1 _17914_ (.A0(\rvcpu.dp.plde.ImmExtE[30] ),
    .A1(\rvcpu.dp.SrcBFW_Mux.y[30] ),
    .S(_05279_),
    .X(_05287_));
 sky130_fd_sc_hd__nand2_1 _17915_ (.A(_05286_),
    .B(_05287_),
    .Y(_05288_));
 sky130_fd_sc_hd__or2_1 _17916_ (.A(_05286_),
    .B(_05287_),
    .X(_05289_));
 sky130_fd_sc_hd__nand2_2 _17917_ (.A(_05288_),
    .B(_05289_),
    .Y(_05290_));
 sky130_fd_sc_hd__nand2_4 _17918_ (.A(_05252_),
    .B(_05263_),
    .Y(_05291_));
 sky130_fd_sc_hd__clkbuf_4 _17919_ (.A(_05291_),
    .X(_05292_));
 sky130_fd_sc_hd__clkbuf_4 _17920_ (.A(_05252_),
    .X(_05293_));
 sky130_fd_sc_hd__or2_2 _17921_ (.A(_05268_),
    .B(_05263_),
    .X(_05294_));
 sky130_fd_sc_hd__o22a_1 _17922_ (.A1(\rvcpu.dp.plem.ALUResultM[29] ),
    .A2(_05293_),
    .B1(_05294_),
    .B2(_13186_),
    .X(_05295_));
 sky130_fd_sc_hd__o21a_1 _17923_ (.A1(\rvcpu.dp.plde.RD1E[29] ),
    .A2(_05292_),
    .B1(_05295_),
    .X(_05296_));
 sky130_fd_sc_hd__mux2_1 _17924_ (.A0(\rvcpu.dp.plde.ImmExtE[29] ),
    .A1(\rvcpu.dp.SrcBFW_Mux.y[29] ),
    .S(_05279_),
    .X(_05297_));
 sky130_fd_sc_hd__nor2_2 _17925_ (.A(_05296_),
    .B(_05297_),
    .Y(_05298_));
 sky130_fd_sc_hd__or2_1 _17926_ (.A(\rvcpu.dp.plem.ALUResultM[28] ),
    .B(_05252_),
    .X(_05299_));
 sky130_fd_sc_hd__o221a_2 _17927_ (.A1(\rvcpu.dp.plde.RD1E[28] ),
    .A2(_05291_),
    .B1(_05294_),
    .B2(_13189_),
    .C1(_05299_),
    .X(_05300_));
 sky130_fd_sc_hd__mux2_1 _17928_ (.A0(\rvcpu.dp.plde.ImmExtE[28] ),
    .A1(\rvcpu.dp.SrcBFW_Mux.y[28] ),
    .S(_05279_),
    .X(_05301_));
 sky130_fd_sc_hd__and2_1 _17929_ (.A(_05300_),
    .B(_05301_),
    .X(_05302_));
 sky130_fd_sc_hd__nor2_1 _17930_ (.A(_05300_),
    .B(_05301_),
    .Y(_05303_));
 sky130_fd_sc_hd__or2_1 _17931_ (.A(_05302_),
    .B(_05303_),
    .X(_05304_));
 sky130_fd_sc_hd__buf_2 _17932_ (.A(_05304_),
    .X(_05305_));
 sky130_fd_sc_hd__and3_1 _17933_ (.A(\rvcpu.dp.plde.RD1E[14] ),
    .B(_05293_),
    .C(_05263_),
    .X(_05306_));
 sky130_fd_sc_hd__a221oi_2 _17934_ (.A1(\rvcpu.dp.plem.ALUResultM[14] ),
    .A2(_05272_),
    .B1(_05270_),
    .B2(_13234_),
    .C1(_05306_),
    .Y(_05307_));
 sky130_fd_sc_hd__mux2_1 _17935_ (.A0(_13234_),
    .A1(\rvcpu.dp.plde.RD2E[14] ),
    .S(_05194_),
    .X(_05308_));
 sky130_fd_sc_hd__mux2_1 _17936_ (.A0(\rvcpu.dp.plem.ALUResultM[14] ),
    .A1(_05308_),
    .S(_05176_),
    .X(_05309_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17937_ (.A(_05309_),
    .X(\rvcpu.dp.SrcBFW_Mux.y[14] ));
 sky130_fd_sc_hd__mux2_2 _17938_ (.A0(\rvcpu.dp.plde.ImmExtE[14] ),
    .A1(\rvcpu.dp.SrcBFW_Mux.y[14] ),
    .S(_05277_),
    .X(_05310_));
 sky130_fd_sc_hd__xnor2_4 _17939_ (.A(net105),
    .B(_05310_),
    .Y(_05311_));
 sky130_fd_sc_hd__and2_1 _17940_ (.A(\rvcpu.dp.plem.ALUResultM[15] ),
    .B(_05272_),
    .X(_05312_));
 sky130_fd_sc_hd__a221o_2 _17941_ (.A1(\rvcpu.dp.plde.RD1E[15] ),
    .A2(_05267_),
    .B1(_05271_),
    .B2(_13231_),
    .C1(_05312_),
    .X(_05313_));
 sky130_fd_sc_hd__mux2_1 _17942_ (.A0(\rvcpu.dp.plde.ImmExtE[15] ),
    .A1(\rvcpu.dp.SrcBFW_Mux.y[15] ),
    .S(_05277_),
    .X(_05314_));
 sky130_fd_sc_hd__nand2_1 _17943_ (.A(_05313_),
    .B(_05314_),
    .Y(_05315_));
 sky130_fd_sc_hd__or2_1 _17944_ (.A(_05313_),
    .B(_05314_),
    .X(_05316_));
 sky130_fd_sc_hd__and2_1 _17945_ (.A(_05315_),
    .B(_05316_),
    .X(_05317_));
 sky130_fd_sc_hd__clkbuf_2 _17946_ (.A(_05317_),
    .X(_05318_));
 sky130_fd_sc_hd__and2_1 _17947_ (.A(\rvcpu.dp.plem.ALUResultM[13] ),
    .B(_05268_),
    .X(_05319_));
 sky130_fd_sc_hd__a221o_2 _17948_ (.A1(\rvcpu.dp.plde.RD1E[13] ),
    .A2(_05266_),
    .B1(_05270_),
    .B2(_13237_),
    .C1(_05319_),
    .X(_05320_));
 sky130_fd_sc_hd__buf_4 _17949_ (.A(\rvcpu.dp.plde.ALUSrcE ),
    .X(_05321_));
 sky130_fd_sc_hd__nand2_1 _17950_ (.A(_05321_),
    .B(\rvcpu.dp.plde.ImmExtE[13] ),
    .Y(_05322_));
 sky130_fd_sc_hd__o31ai_4 _17951_ (.A1(_05321_),
    .A2(_05226_),
    .A3(_05227_),
    .B1(_05322_),
    .Y(_05323_));
 sky130_fd_sc_hd__nor2_1 _17952_ (.A(_05320_),
    .B(_05323_),
    .Y(_05324_));
 sky130_fd_sc_hd__inv_2 _17953_ (.A(_05324_),
    .Y(_05325_));
 sky130_fd_sc_hd__and2_1 _17954_ (.A(\rvcpu.dp.plem.ALUResultM[12] ),
    .B(_05268_),
    .X(_05326_));
 sky130_fd_sc_hd__a221o_2 _17955_ (.A1(\rvcpu.dp.plde.RD1E[12] ),
    .A2(_05265_),
    .B1(_05269_),
    .B2(_13240_),
    .C1(_05326_),
    .X(_05327_));
 sky130_fd_sc_hd__mux2_1 _17956_ (.A0(_13240_),
    .A1(\rvcpu.dp.plde.RD2E[12] ),
    .S(_05194_),
    .X(_05328_));
 sky130_fd_sc_hd__mux2_1 _17957_ (.A0(\rvcpu.dp.plem.ALUResultM[12] ),
    .A1(_05328_),
    .S(_05175_),
    .X(_05329_));
 sky130_fd_sc_hd__buf_1 _17958_ (.A(_05329_),
    .X(\rvcpu.dp.SrcBFW_Mux.y[12] ));
 sky130_fd_sc_hd__mux2_1 _17959_ (.A0(\rvcpu.dp.plde.ImmExtE[12] ),
    .A1(\rvcpu.dp.SrcBFW_Mux.y[12] ),
    .S(_05277_),
    .X(_05330_));
 sky130_fd_sc_hd__and2_1 _17960_ (.A(_05327_),
    .B(_05330_),
    .X(_05331_));
 sky130_fd_sc_hd__and2_1 _17961_ (.A(_05320_),
    .B(_05323_),
    .X(_05332_));
 sky130_fd_sc_hd__a21o_1 _17962_ (.A1(_05325_),
    .A2(_05331_),
    .B1(_05332_),
    .X(_05333_));
 sky130_fd_sc_hd__a221o_2 _17963_ (.A1(\rvcpu.dp.plem.ALUResultM[14] ),
    .A2(_05272_),
    .B1(_05270_),
    .B2(_13234_),
    .C1(_05306_),
    .X(_05334_));
 sky130_fd_sc_hd__and2_1 _17964_ (.A(_05334_),
    .B(_05310_),
    .X(_05335_));
 sky130_fd_sc_hd__a21bo_1 _17965_ (.A1(_05335_),
    .A2(_05316_),
    .B1_N(_05315_),
    .X(_05336_));
 sky130_fd_sc_hd__a31oi_1 _17966_ (.A1(_05311_),
    .A2(_05318_),
    .A3(_05333_),
    .B1(_05336_),
    .Y(_05337_));
 sky130_fd_sc_hd__inv_2 _17967_ (.A(_05337_),
    .Y(_05338_));
 sky130_fd_sc_hd__buf_2 _17968_ (.A(_05293_),
    .X(_05339_));
 sky130_fd_sc_hd__clkbuf_4 _17969_ (.A(_05294_),
    .X(_05340_));
 sky130_fd_sc_hd__o22a_1 _17970_ (.A1(\rvcpu.dp.plem.ALUResultM[7] ),
    .A2(_05339_),
    .B1(_05340_),
    .B2(_13256_),
    .X(_05341_));
 sky130_fd_sc_hd__o21a_2 _17971_ (.A1(\rvcpu.dp.plde.RD1E[7] ),
    .A2(_05292_),
    .B1(_05341_),
    .X(_05342_));
 sky130_fd_sc_hd__mux2_1 _17972_ (.A0(\rvcpu.dp.plde.ImmExtE[7] ),
    .A1(\rvcpu.dp.SrcBFW_Mux.y[7] ),
    .S(_05278_),
    .X(_05343_));
 sky130_fd_sc_hd__and2_1 _17973_ (.A(_05342_),
    .B(_05343_),
    .X(_05344_));
 sky130_fd_sc_hd__nor2_1 _17974_ (.A(_05342_),
    .B(_05343_),
    .Y(_05345_));
 sky130_fd_sc_hd__nor2_2 _17975_ (.A(_05344_),
    .B(_05345_),
    .Y(_05346_));
 sky130_fd_sc_hd__inv_6 _17976_ (.A(\rvcpu.dp.plem.ALUResultM[6] ),
    .Y(_05347_));
 sky130_fd_sc_hd__nor2_1 _17977_ (.A(_05347_),
    .B(_05339_),
    .Y(_05348_));
 sky130_fd_sc_hd__a221o_4 _17978_ (.A1(\rvcpu.dp.plde.RD1E[6] ),
    .A2(_05267_),
    .B1(_05271_),
    .B2(_13259_),
    .C1(_05348_),
    .X(_05349_));
 sky130_fd_sc_hd__nand3b_1 _17979_ (.A_N(_13259_),
    .B(_05179_),
    .C(_05180_),
    .Y(_05350_));
 sky130_fd_sc_hd__a21o_1 _17980_ (.A1(_05179_),
    .A2(_05180_),
    .B1(\rvcpu.dp.plde.RD2E[6] ),
    .X(_05351_));
 sky130_fd_sc_hd__nor2_1 _17981_ (.A(_05347_),
    .B(_05176_),
    .Y(_05352_));
 sky130_fd_sc_hd__a31o_1 _17982_ (.A1(_05176_),
    .A2(_05350_),
    .A3(_05351_),
    .B1(_05352_),
    .X(\rvcpu.dp.SrcBFW_Mux.y[6] ));
 sky130_fd_sc_hd__mux2_1 _17983_ (.A0(\rvcpu.dp.plde.ImmExtE[6] ),
    .A1(\rvcpu.dp.SrcBFW_Mux.y[6] ),
    .S(_05277_),
    .X(_05353_));
 sky130_fd_sc_hd__and2_1 _17984_ (.A(_05349_),
    .B(_05353_),
    .X(_05354_));
 sky130_fd_sc_hd__nor2_1 _17985_ (.A(_05349_),
    .B(_05353_),
    .Y(_05355_));
 sky130_fd_sc_hd__nor2_2 _17986_ (.A(_05354_),
    .B(_05355_),
    .Y(_05356_));
 sky130_fd_sc_hd__and2_1 _17987_ (.A(\rvcpu.dp.plem.ALUResultM[5] ),
    .B(_05272_),
    .X(_05357_));
 sky130_fd_sc_hd__a221o_4 _17988_ (.A1(\rvcpu.dp.plde.RD1E[5] ),
    .A2(_05266_),
    .B1(_05270_),
    .B2(_13262_),
    .C1(_05357_),
    .X(_05358_));
 sky130_fd_sc_hd__mux2_2 _17989_ (.A0(\rvcpu.dp.plde.ImmExtE[5] ),
    .A1(\rvcpu.dp.SrcBFW_Mux.y[5] ),
    .S(_05277_),
    .X(_05359_));
 sky130_fd_sc_hd__nor2_1 _17990_ (.A(_05358_),
    .B(_05359_),
    .Y(_05360_));
 sky130_fd_sc_hd__inv_2 _17991_ (.A(_05360_),
    .Y(_05361_));
 sky130_fd_sc_hd__or2_1 _17992_ (.A(_05277_),
    .B(\rvcpu.dp.plde.ImmExtE[4] ),
    .X(_05362_));
 sky130_fd_sc_hd__o21ai_4 _17993_ (.A1(_05321_),
    .A2(\rvcpu.dp.SrcBFW_Mux.y[4] ),
    .B1(_05362_),
    .Y(_05363_));
 sky130_fd_sc_hd__o22a_1 _17994_ (.A1(\rvcpu.dp.plem.ALUResultM[4] ),
    .A2(_05339_),
    .B1(_05340_),
    .B2(_13265_),
    .X(_05364_));
 sky130_fd_sc_hd__o21ai_4 _17995_ (.A1(\rvcpu.dp.plde.RD1E[4] ),
    .A2(_05291_),
    .B1(_05364_),
    .Y(_05365_));
 sky130_fd_sc_hd__nor2_1 _17996_ (.A(_05363_),
    .B(_05365_),
    .Y(_05366_));
 sky130_fd_sc_hd__nand2_1 _17997_ (.A(_05363_),
    .B(_05365_),
    .Y(_05367_));
 sky130_fd_sc_hd__nor2b_2 _17998_ (.A(_05366_),
    .B_N(_05367_),
    .Y(_05368_));
 sky130_fd_sc_hd__or2_1 _17999_ (.A(_05276_),
    .B(\rvcpu.dp.plde.ImmExtE[3] ),
    .X(_05369_));
 sky130_fd_sc_hd__o21a_2 _18000_ (.A1(_05321_),
    .A2(\rvcpu.dp.SrcBFW_Mux.y[3] ),
    .B1(_05369_),
    .X(_05370_));
 sky130_fd_sc_hd__inv_4 _18001_ (.A(\rvcpu.dp.plem.ALUResultM[3] ),
    .Y(_05371_));
 sky130_fd_sc_hd__nor2_1 _18002_ (.A(_05371_),
    .B(_05293_),
    .Y(_05372_));
 sky130_fd_sc_hd__a221o_2 _18003_ (.A1(\rvcpu.dp.plde.RD1E[3] ),
    .A2(_05265_),
    .B1(_05269_),
    .B2(_13268_),
    .C1(_05372_),
    .X(_05373_));
 sky130_fd_sc_hd__nand2_1 _18004_ (.A(_05370_),
    .B(_05373_),
    .Y(_05374_));
 sky130_fd_sc_hd__o21ai_4 _18005_ (.A1(_05321_),
    .A2(\rvcpu.dp.SrcBFW_Mux.y[3] ),
    .B1(_05369_),
    .Y(_05375_));
 sky130_fd_sc_hd__inv_2 _18006_ (.A(_05373_),
    .Y(_05376_));
 sky130_fd_sc_hd__nand2_1 _18007_ (.A(_05375_),
    .B(_05376_),
    .Y(_05377_));
 sky130_fd_sc_hd__and2_1 _18008_ (.A(_05374_),
    .B(_05377_),
    .X(_05378_));
 sky130_fd_sc_hd__or2_1 _18009_ (.A(_05277_),
    .B(\rvcpu.dp.plde.ImmExtE[2] ),
    .X(_05379_));
 sky130_fd_sc_hd__o21a_2 _18010_ (.A1(_05321_),
    .A2(\rvcpu.dp.SrcBFW_Mux.y[2] ),
    .B1(_05379_),
    .X(_05380_));
 sky130_fd_sc_hd__a22o_1 _18011_ (.A1(net122),
    .A2(_05268_),
    .B1(_05269_),
    .B2(_13271_),
    .X(_05381_));
 sky130_fd_sc_hd__a21oi_4 _18012_ (.A1(\rvcpu.dp.plde.RD1E[2] ),
    .A2(_05266_),
    .B1(_05381_),
    .Y(_05382_));
 sky130_fd_sc_hd__xnor2_2 _18013_ (.A(_05380_),
    .B(_05382_),
    .Y(_05383_));
 sky130_fd_sc_hd__nand2_1 _18014_ (.A(_05321_),
    .B(\rvcpu.dp.plde.ImmExtE[1] ),
    .Y(_05384_));
 sky130_fd_sc_hd__o221ai_4 _18015_ (.A1(\rvcpu.dp.plem.ALUResultM[1] ),
    .A2(_05175_),
    .B1(_05181_),
    .B2(_05182_),
    .C1(_05276_),
    .Y(_05385_));
 sky130_fd_sc_hd__inv_2 _18016_ (.A(\rvcpu.dp.plem.ALUResultM[1] ),
    .Y(_05386_));
 sky130_fd_sc_hd__nor2_1 _18017_ (.A(_05386_),
    .B(_05293_),
    .Y(_05387_));
 sky130_fd_sc_hd__a221oi_4 _18018_ (.A1(\rvcpu.dp.plde.RD1E[1] ),
    .A2(_05265_),
    .B1(_05269_),
    .B2(_13274_),
    .C1(_05387_),
    .Y(_05388_));
 sky130_fd_sc_hd__nand3_1 _18019_ (.A(_05384_),
    .B(_05385_),
    .C(_05388_),
    .Y(_05389_));
 sky130_fd_sc_hd__nand2_1 _18020_ (.A(\rvcpu.dp.plde.ImmExtE[0] ),
    .B(_05321_),
    .Y(_05390_));
 sky130_fd_sc_hd__inv_2 _18021_ (.A(\rvcpu.dp.plem.ALUResultM[0] ),
    .Y(_05391_));
 sky130_fd_sc_hd__a221o_1 _18022_ (.A1(_05391_),
    .A2(net115),
    .B1(_05173_),
    .B2(_05172_),
    .C1(\rvcpu.dp.plde.ALUSrcE ),
    .X(_05392_));
 sky130_fd_sc_hd__nor2_1 _18023_ (.A(_05391_),
    .B(_05293_),
    .Y(_05393_));
 sky130_fd_sc_hd__a221oi_4 _18024_ (.A1(\rvcpu.dp.plde.RD1E[0] ),
    .A2(_05265_),
    .B1(_05269_),
    .B2(_13277_),
    .C1(_05393_),
    .Y(_05394_));
 sky130_fd_sc_hd__a21oi_2 _18025_ (.A1(_05390_),
    .A2(_05392_),
    .B1(_05394_),
    .Y(_05395_));
 sky130_fd_sc_hd__a21oi_1 _18026_ (.A1(_05384_),
    .A2(_05385_),
    .B1(_05388_),
    .Y(_05396_));
 sky130_fd_sc_hd__a21o_1 _18027_ (.A1(_05389_),
    .A2(_05395_),
    .B1(_05396_),
    .X(_05397_));
 sky130_fd_sc_hd__o21ai_2 _18028_ (.A1(_05321_),
    .A2(\rvcpu.dp.SrcBFW_Mux.y[2] ),
    .B1(_05379_),
    .Y(_05398_));
 sky130_fd_sc_hd__nor2_1 _18029_ (.A(_05398_),
    .B(_05382_),
    .Y(_05399_));
 sky130_fd_sc_hd__a21o_1 _18030_ (.A1(_05383_),
    .A2(_05397_),
    .B1(_05399_),
    .X(_05400_));
 sky130_fd_sc_hd__a21bo_1 _18031_ (.A1(_05378_),
    .A2(_05400_),
    .B1_N(_05374_),
    .X(_05401_));
 sky130_fd_sc_hd__nand2_1 _18032_ (.A(_05358_),
    .B(_05359_),
    .Y(_05402_));
 sky130_fd_sc_hd__inv_2 _18033_ (.A(_05402_),
    .Y(_05403_));
 sky130_fd_sc_hd__a211o_1 _18034_ (.A1(_05368_),
    .A2(_05401_),
    .B1(_05403_),
    .C1(_05366_),
    .X(_05404_));
 sky130_fd_sc_hd__a31o_1 _18035_ (.A1(_05356_),
    .A2(_05361_),
    .A3(_05404_),
    .B1(_05354_),
    .X(_05405_));
 sky130_fd_sc_hd__a21o_1 _18036_ (.A1(_05346_),
    .A2(_05405_),
    .B1(_05344_),
    .X(_05406_));
 sky130_fd_sc_hd__and2_1 _18037_ (.A(\rvcpu.dp.plem.ALUResultM[11] ),
    .B(_05272_),
    .X(_05407_));
 sky130_fd_sc_hd__a221oi_4 _18038_ (.A1(\rvcpu.dp.plde.RD1E[11] ),
    .A2(_05267_),
    .B1(_05271_),
    .B2(_13243_),
    .C1(_05407_),
    .Y(_05408_));
 sky130_fd_sc_hd__mux2_2 _18039_ (.A0(\rvcpu.dp.plde.ImmExtE[11] ),
    .A1(\rvcpu.dp.SrcBFW_Mux.y[11] ),
    .S(_05277_),
    .X(_05409_));
 sky130_fd_sc_hd__xnor2_4 _18040_ (.A(net103),
    .B(_05409_),
    .Y(_05410_));
 sky130_fd_sc_hd__and2_1 _18041_ (.A(\rvcpu.dp.plem.ALUResultM[10] ),
    .B(_05272_),
    .X(_05411_));
 sky130_fd_sc_hd__a221o_2 _18042_ (.A1(\rvcpu.dp.plde.RD1E[10] ),
    .A2(_05267_),
    .B1(_05271_),
    .B2(_13247_),
    .C1(_05411_),
    .X(_05412_));
 sky130_fd_sc_hd__mux2_1 _18043_ (.A0(_13247_),
    .A1(\rvcpu.dp.plde.RD2E[10] ),
    .S(_05195_),
    .X(_05413_));
 sky130_fd_sc_hd__mux2_1 _18044_ (.A0(\rvcpu.dp.plem.ALUResultM[10] ),
    .A1(_05413_),
    .S(_05176_),
    .X(_05414_));
 sky130_fd_sc_hd__buf_1 _18045_ (.A(_05414_),
    .X(\rvcpu.dp.SrcBFW_Mux.y[10] ));
 sky130_fd_sc_hd__mux2_1 _18046_ (.A0(\rvcpu.dp.plde.ImmExtE[10] ),
    .A1(\rvcpu.dp.SrcBFW_Mux.y[10] ),
    .S(_05278_),
    .X(_05415_));
 sky130_fd_sc_hd__and2_1 _18047_ (.A(_05412_),
    .B(_05415_),
    .X(_05416_));
 sky130_fd_sc_hd__nor2_1 _18048_ (.A(_05412_),
    .B(_05415_),
    .Y(_05417_));
 sky130_fd_sc_hd__nor2_1 _18049_ (.A(_05416_),
    .B(_05417_),
    .Y(_05418_));
 sky130_fd_sc_hd__buf_2 _18050_ (.A(_05418_),
    .X(_05419_));
 sky130_fd_sc_hd__and2_1 _18051_ (.A(_13253_),
    .B(_05271_),
    .X(_05420_));
 sky130_fd_sc_hd__a221o_2 _18052_ (.A1(\rvcpu.dp.plem.ALUResultM[8] ),
    .A2(_05272_),
    .B1(_05267_),
    .B2(\rvcpu.dp.plde.RD1E[8] ),
    .C1(_05420_),
    .X(_05421_));
 sky130_fd_sc_hd__mux2_1 _18053_ (.A0(_13253_),
    .A1(\rvcpu.dp.plde.RD2E[8] ),
    .S(_05195_),
    .X(_05422_));
 sky130_fd_sc_hd__mux2_1 _18054_ (.A0(\rvcpu.dp.plem.ALUResultM[8] ),
    .A1(_05422_),
    .S(_05177_),
    .X(_05423_));
 sky130_fd_sc_hd__buf_1 _18055_ (.A(_05423_),
    .X(\rvcpu.dp.SrcBFW_Mux.y[8] ));
 sky130_fd_sc_hd__mux2_1 _18056_ (.A0(\rvcpu.dp.plde.ImmExtE[8] ),
    .A1(\rvcpu.dp.SrcBFW_Mux.y[8] ),
    .S(_05278_),
    .X(_05424_));
 sky130_fd_sc_hd__and2_1 _18057_ (.A(_05421_),
    .B(_05424_),
    .X(_05425_));
 sky130_fd_sc_hd__nor2_1 _18058_ (.A(_05421_),
    .B(_05424_),
    .Y(_05426_));
 sky130_fd_sc_hd__nor2_1 _18059_ (.A(_05425_),
    .B(_05426_),
    .Y(_05427_));
 sky130_fd_sc_hd__and2_1 _18060_ (.A(\rvcpu.dp.plem.ALUResultM[9] ),
    .B(_05272_),
    .X(_05428_));
 sky130_fd_sc_hd__a221oi_2 _18061_ (.A1(\rvcpu.dp.plde.RD1E[9] ),
    .A2(_05267_),
    .B1(_05271_),
    .B2(_13250_),
    .C1(_05428_),
    .Y(_05429_));
 sky130_fd_sc_hd__mux2_2 _18062_ (.A0(\rvcpu.dp.plde.ImmExtE[9] ),
    .A1(\rvcpu.dp.SrcBFW_Mux.y[9] ),
    .S(_05277_),
    .X(_05430_));
 sky130_fd_sc_hd__xnor2_2 _18063_ (.A(net102),
    .B(_05430_),
    .Y(_05431_));
 sky130_fd_sc_hd__nand4_1 _18064_ (.A(_05410_),
    .B(_05419_),
    .C(_05427_),
    .D(_05431_),
    .Y(_05432_));
 sky130_fd_sc_hd__inv_2 _18065_ (.A(_05432_),
    .Y(_05433_));
 sky130_fd_sc_hd__or2_1 _18066_ (.A(_05327_),
    .B(_05330_),
    .X(_05434_));
 sky130_fd_sc_hd__and2b_1 _18067_ (.A_N(_05331_),
    .B(_05434_),
    .X(_05435_));
 sky130_fd_sc_hd__buf_2 _18068_ (.A(_05435_),
    .X(_05436_));
 sky130_fd_sc_hd__a221oi_4 _18069_ (.A1(\rvcpu.dp.plde.RD1E[13] ),
    .A2(_05266_),
    .B1(_05270_),
    .B2(_13237_),
    .C1(_05319_),
    .Y(_05437_));
 sky130_fd_sc_hd__xnor2_2 _18070_ (.A(_05437_),
    .B(_05323_),
    .Y(_05438_));
 sky130_fd_sc_hd__nand4_1 _18071_ (.A(_05311_),
    .B(_05318_),
    .C(_05436_),
    .D(_05438_),
    .Y(_05439_));
 sky130_fd_sc_hd__inv_2 _18072_ (.A(_05439_),
    .Y(_05440_));
 sky130_fd_sc_hd__a221o_2 _18073_ (.A1(\rvcpu.dp.plde.RD1E[9] ),
    .A2(_05267_),
    .B1(_05271_),
    .B2(_13250_),
    .C1(_05428_),
    .X(_05441_));
 sky130_fd_sc_hd__nor2_1 _18074_ (.A(_05441_),
    .B(_05430_),
    .Y(_05442_));
 sky130_fd_sc_hd__inv_2 _18075_ (.A(_05425_),
    .Y(_05443_));
 sky130_fd_sc_hd__and2_1 _18076_ (.A(_05441_),
    .B(_05430_),
    .X(_05444_));
 sky130_fd_sc_hd__o21bai_1 _18077_ (.A1(_05442_),
    .A2(_05443_),
    .B1_N(_05444_),
    .Y(_05445_));
 sky130_fd_sc_hd__a221o_2 _18078_ (.A1(\rvcpu.dp.plde.RD1E[11] ),
    .A2(_05266_),
    .B1(_05270_),
    .B2(_13243_),
    .C1(_05407_),
    .X(_05446_));
 sky130_fd_sc_hd__nor2_1 _18079_ (.A(_05446_),
    .B(_05409_),
    .Y(_05447_));
 sky130_fd_sc_hd__inv_2 _18080_ (.A(_05416_),
    .Y(_05448_));
 sky130_fd_sc_hd__nand2_1 _18081_ (.A(_05446_),
    .B(_05409_),
    .Y(_05449_));
 sky130_fd_sc_hd__o21ai_1 _18082_ (.A1(_05447_),
    .A2(_05448_),
    .B1(_05449_),
    .Y(_05450_));
 sky130_fd_sc_hd__a31o_1 _18083_ (.A1(_05410_),
    .A2(_05419_),
    .A3(_05445_),
    .B1(_05450_),
    .X(_05451_));
 sky130_fd_sc_hd__and2_1 _18084_ (.A(_05451_),
    .B(_05440_),
    .X(_05452_));
 sky130_fd_sc_hd__a31o_1 _18085_ (.A1(_05406_),
    .A2(_05433_),
    .A3(_05440_),
    .B1(_05452_),
    .X(_05453_));
 sky130_fd_sc_hd__or2_2 _18086_ (.A(_05338_),
    .B(_05453_),
    .X(_05454_));
 sky130_fd_sc_hd__o22a_1 _18087_ (.A1(\rvcpu.dp.plem.ALUResultM[23] ),
    .A2(_05339_),
    .B1(_05340_),
    .B2(_13206_),
    .X(_05455_));
 sky130_fd_sc_hd__o21a_2 _18088_ (.A1(\rvcpu.dp.plde.RD1E[23] ),
    .A2(_05292_),
    .B1(_05455_),
    .X(_05456_));
 sky130_fd_sc_hd__mux2_1 _18089_ (.A0(\rvcpu.dp.plde.ImmExtE[23] ),
    .A1(\rvcpu.dp.SrcBFW_Mux.y[23] ),
    .S(_05278_),
    .X(_05457_));
 sky130_fd_sc_hd__or2_1 _18090_ (.A(_05456_),
    .B(_05457_),
    .X(_05458_));
 sky130_fd_sc_hd__nand2_1 _18091_ (.A(_05456_),
    .B(_05457_),
    .Y(_05459_));
 sky130_fd_sc_hd__and2_1 _18092_ (.A(_05458_),
    .B(_05459_),
    .X(_05460_));
 sky130_fd_sc_hd__buf_2 _18093_ (.A(_05460_),
    .X(_05461_));
 sky130_fd_sc_hd__o22a_1 _18094_ (.A1(\rvcpu.dp.plem.ALUResultM[22] ),
    .A2(_05339_),
    .B1(_05340_),
    .B2(_13209_),
    .X(_05462_));
 sky130_fd_sc_hd__o21a_2 _18095_ (.A1(\rvcpu.dp.plde.RD1E[22] ),
    .A2(_05292_),
    .B1(_05462_),
    .X(_05463_));
 sky130_fd_sc_hd__mux2_1 _18096_ (.A0(\rvcpu.dp.plde.ImmExtE[22] ),
    .A1(\rvcpu.dp.SrcBFW_Mux.y[22] ),
    .S(_05279_),
    .X(_05464_));
 sky130_fd_sc_hd__nor2_1 _18097_ (.A(_05463_),
    .B(_05464_),
    .Y(_05465_));
 sky130_fd_sc_hd__and2_1 _18098_ (.A(_05463_),
    .B(_05464_),
    .X(_05466_));
 sky130_fd_sc_hd__nor2_2 _18099_ (.A(_05465_),
    .B(_05466_),
    .Y(_05467_));
 sky130_fd_sc_hd__o22a_1 _18100_ (.A1(\rvcpu.dp.plem.ALUResultM[21] ),
    .A2(_05339_),
    .B1(_05340_),
    .B2(_13212_),
    .X(_05468_));
 sky130_fd_sc_hd__o21a_2 _18101_ (.A1(\rvcpu.dp.plde.RD1E[21] ),
    .A2(_05292_),
    .B1(_05468_),
    .X(_05469_));
 sky130_fd_sc_hd__mux2_1 _18102_ (.A0(\rvcpu.dp.plde.ImmExtE[21] ),
    .A1(\rvcpu.dp.SrcBFW_Mux.y[21] ),
    .S(_05278_),
    .X(_05470_));
 sky130_fd_sc_hd__nor2_1 _18103_ (.A(_05469_),
    .B(_05470_),
    .Y(_05471_));
 sky130_fd_sc_hd__and2_1 _18104_ (.A(_05469_),
    .B(_05470_),
    .X(_05472_));
 sky130_fd_sc_hd__nor2_2 _18105_ (.A(_05471_),
    .B(_05472_),
    .Y(_05473_));
 sky130_fd_sc_hd__o22a_1 _18106_ (.A1(\rvcpu.dp.plem.ALUResultM[20] ),
    .A2(_05339_),
    .B1(_05340_),
    .B2(_13216_),
    .X(_05474_));
 sky130_fd_sc_hd__o21a_2 _18107_ (.A1(\rvcpu.dp.plde.RD1E[20] ),
    .A2(_05292_),
    .B1(_05474_),
    .X(_05475_));
 sky130_fd_sc_hd__mux2_1 _18108_ (.A0(_13216_),
    .A1(\rvcpu.dp.plde.RD2E[20] ),
    .S(_05196_),
    .X(_05476_));
 sky130_fd_sc_hd__mux2_1 _18109_ (.A0(\rvcpu.dp.plem.ALUResultM[20] ),
    .A1(_05476_),
    .S(_05177_),
    .X(_05477_));
 sky130_fd_sc_hd__clkbuf_2 _18110_ (.A(_05477_),
    .X(\rvcpu.dp.SrcBFW_Mux.y[20] ));
 sky130_fd_sc_hd__mux2_1 _18111_ (.A0(\rvcpu.dp.plde.ImmExtE[20] ),
    .A1(\rvcpu.dp.SrcBFW_Mux.y[20] ),
    .S(_05279_),
    .X(_05478_));
 sky130_fd_sc_hd__and2_1 _18112_ (.A(_05475_),
    .B(_05478_),
    .X(_05479_));
 sky130_fd_sc_hd__nor2_1 _18113_ (.A(_05475_),
    .B(_05478_),
    .Y(_05480_));
 sky130_fd_sc_hd__nor2_2 _18114_ (.A(_05479_),
    .B(_05480_),
    .Y(_05481_));
 sky130_fd_sc_hd__and4_1 _18115_ (.A(_05461_),
    .B(_05467_),
    .C(_05473_),
    .D(_05481_),
    .X(_05482_));
 sky130_fd_sc_hd__o22a_1 _18116_ (.A1(\rvcpu.dp.plem.ALUResultM[19] ),
    .A2(_05339_),
    .B1(_05340_),
    .B2(_13219_),
    .X(_05483_));
 sky130_fd_sc_hd__o21a_2 _18117_ (.A1(\rvcpu.dp.plde.RD1E[19] ),
    .A2(_05292_),
    .B1(_05483_),
    .X(_05484_));
 sky130_fd_sc_hd__mux2_1 _18118_ (.A0(\rvcpu.dp.plde.ImmExtE[19] ),
    .A1(\rvcpu.dp.SrcBFW_Mux.y[19] ),
    .S(_05278_),
    .X(_05485_));
 sky130_fd_sc_hd__nor2_1 _18119_ (.A(_05484_),
    .B(_05485_),
    .Y(_05486_));
 sky130_fd_sc_hd__nand2_1 _18120_ (.A(_05484_),
    .B(_05485_),
    .Y(_05487_));
 sky130_fd_sc_hd__and2b_1 _18121_ (.A_N(_05486_),
    .B(_05487_),
    .X(_05488_));
 sky130_fd_sc_hd__o22a_1 _18122_ (.A1(\rvcpu.dp.plem.ALUResultM[18] ),
    .A2(_05339_),
    .B1(_05340_),
    .B2(_13222_),
    .X(_05489_));
 sky130_fd_sc_hd__o21a_2 _18123_ (.A1(\rvcpu.dp.plde.RD1E[18] ),
    .A2(_05292_),
    .B1(_05489_),
    .X(_05490_));
 sky130_fd_sc_hd__mux2_1 _18124_ (.A0(_13222_),
    .A1(\rvcpu.dp.plde.RD2E[18] ),
    .S(_05194_),
    .X(_05491_));
 sky130_fd_sc_hd__mux2_1 _18125_ (.A0(\rvcpu.dp.plem.ALUResultM[18] ),
    .A1(_05491_),
    .S(_05176_),
    .X(_05492_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _18126_ (.A(_05492_),
    .X(\rvcpu.dp.SrcBFW_Mux.y[18] ));
 sky130_fd_sc_hd__mux2_1 _18127_ (.A0(\rvcpu.dp.plde.ImmExtE[18] ),
    .A1(\rvcpu.dp.SrcBFW_Mux.y[18] ),
    .S(_05278_),
    .X(_05493_));
 sky130_fd_sc_hd__nand2_1 _18128_ (.A(_05490_),
    .B(_05493_),
    .Y(_05494_));
 sky130_fd_sc_hd__or2_1 _18129_ (.A(_05490_),
    .B(_05493_),
    .X(_05495_));
 sky130_fd_sc_hd__and2_1 _18130_ (.A(_05494_),
    .B(_05495_),
    .X(_05496_));
 sky130_fd_sc_hd__clkbuf_2 _18131_ (.A(_05496_),
    .X(_05497_));
 sky130_fd_sc_hd__and2_1 _18132_ (.A(_05488_),
    .B(_05497_),
    .X(_05498_));
 sky130_fd_sc_hd__o22a_1 _18133_ (.A1(\rvcpu.dp.plem.ALUResultM[17] ),
    .A2(_05339_),
    .B1(_05340_),
    .B2(_13225_),
    .X(_05499_));
 sky130_fd_sc_hd__o21a_2 _18134_ (.A1(\rvcpu.dp.plde.RD1E[17] ),
    .A2(_05292_),
    .B1(_05499_),
    .X(_05500_));
 sky130_fd_sc_hd__mux2_1 _18135_ (.A0(\rvcpu.dp.plde.ImmExtE[17] ),
    .A1(\rvcpu.dp.SrcBFW_Mux.y[17] ),
    .S(_05278_),
    .X(_05501_));
 sky130_fd_sc_hd__and2_1 _18136_ (.A(_05500_),
    .B(_05501_),
    .X(_05502_));
 sky130_fd_sc_hd__nor2_1 _18137_ (.A(_05500_),
    .B(_05501_),
    .Y(_05503_));
 sky130_fd_sc_hd__nor2_2 _18138_ (.A(_05502_),
    .B(_05503_),
    .Y(_05504_));
 sky130_fd_sc_hd__and2_1 _18139_ (.A(\rvcpu.dp.plem.ALUResultM[16] ),
    .B(_05268_),
    .X(_05505_));
 sky130_fd_sc_hd__a221o_4 _18140_ (.A1(\rvcpu.dp.plde.RD1E[16] ),
    .A2(_05265_),
    .B1(_05269_),
    .B2(_13228_),
    .C1(_05505_),
    .X(_05506_));
 sky130_fd_sc_hd__mux2_1 _18141_ (.A0(_13228_),
    .A1(\rvcpu.dp.plde.RD2E[16] ),
    .S(_05195_),
    .X(_05507_));
 sky130_fd_sc_hd__mux2_1 _18142_ (.A0(\rvcpu.dp.plem.ALUResultM[16] ),
    .A1(_05507_),
    .S(_05177_),
    .X(_05508_));
 sky130_fd_sc_hd__buf_1 _18143_ (.A(_05508_),
    .X(\rvcpu.dp.SrcBFW_Mux.y[16] ));
 sky130_fd_sc_hd__mux2_1 _18144_ (.A0(\rvcpu.dp.plde.ImmExtE[16] ),
    .A1(\rvcpu.dp.SrcBFW_Mux.y[16] ),
    .S(_05278_),
    .X(_05509_));
 sky130_fd_sc_hd__and2_1 _18145_ (.A(_05506_),
    .B(_05509_),
    .X(_05510_));
 sky130_fd_sc_hd__nor2_1 _18146_ (.A(_05506_),
    .B(_05509_),
    .Y(_05511_));
 sky130_fd_sc_hd__nor2_1 _18147_ (.A(_05510_),
    .B(_05511_),
    .Y(_05512_));
 sky130_fd_sc_hd__buf_2 _18148_ (.A(_05512_),
    .X(_05513_));
 sky130_fd_sc_hd__and3_1 _18149_ (.A(_05498_),
    .B(_05504_),
    .C(_05513_),
    .X(_05514_));
 sky130_fd_sc_hd__nor2_1 _18150_ (.A(_05502_),
    .B(_05510_),
    .Y(_05515_));
 sky130_fd_sc_hd__nor2_1 _18151_ (.A(_05503_),
    .B(_05515_),
    .Y(_05516_));
 sky130_fd_sc_hd__nand2_1 _18152_ (.A(_05498_),
    .B(_05516_),
    .Y(_05517_));
 sky130_fd_sc_hd__o211a_1 _18153_ (.A1(_05486_),
    .A2(_05494_),
    .B1(_05517_),
    .C1(_05487_),
    .X(_05518_));
 sky130_fd_sc_hd__inv_2 _18154_ (.A(_05518_),
    .Y(_05519_));
 sky130_fd_sc_hd__or2_1 _18155_ (.A(_05469_),
    .B(_05470_),
    .X(_05520_));
 sky130_fd_sc_hd__a21o_1 _18156_ (.A1(_05520_),
    .A2(_05479_),
    .B1(_05472_),
    .X(_05521_));
 sky130_fd_sc_hd__a21bo_1 _18157_ (.A1(_05458_),
    .A2(_05466_),
    .B1_N(_05459_),
    .X(_05522_));
 sky130_fd_sc_hd__a31o_1 _18158_ (.A1(_05461_),
    .A2(_05467_),
    .A3(_05521_),
    .B1(_05522_),
    .X(_05523_));
 sky130_fd_sc_hd__a21o_1 _18159_ (.A1(_05482_),
    .A2(_05519_),
    .B1(_05523_),
    .X(_05524_));
 sky130_fd_sc_hd__a31o_2 _18160_ (.A1(_05454_),
    .A2(_05482_),
    .A3(_05514_),
    .B1(_05524_),
    .X(_05525_));
 sky130_fd_sc_hd__o22a_1 _18161_ (.A1(\rvcpu.dp.plem.ALUResultM[25] ),
    .A2(_05293_),
    .B1(_05340_),
    .B2(_13200_),
    .X(_05526_));
 sky130_fd_sc_hd__o21a_1 _18162_ (.A1(\rvcpu.dp.plde.RD1E[25] ),
    .A2(_05291_),
    .B1(_05526_),
    .X(_05527_));
 sky130_fd_sc_hd__mux2_1 _18163_ (.A0(\rvcpu.dp.plde.ImmExtE[25] ),
    .A1(\rvcpu.dp.SrcBFW_Mux.y[25] ),
    .S(_05279_),
    .X(_05528_));
 sky130_fd_sc_hd__and2_1 _18164_ (.A(_05527_),
    .B(_05528_),
    .X(_05529_));
 sky130_fd_sc_hd__nor2_1 _18165_ (.A(_05527_),
    .B(_05528_),
    .Y(_05530_));
 sky130_fd_sc_hd__nor2_2 _18166_ (.A(_05529_),
    .B(_05530_),
    .Y(_05531_));
 sky130_fd_sc_hd__o22a_1 _18167_ (.A1(\rvcpu.dp.plem.ALUResultM[24] ),
    .A2(_05293_),
    .B1(_05294_),
    .B2(_13203_),
    .X(_05532_));
 sky130_fd_sc_hd__o21a_1 _18168_ (.A1(\rvcpu.dp.plde.RD1E[24] ),
    .A2(_05291_),
    .B1(_05532_),
    .X(_05533_));
 sky130_fd_sc_hd__mux2_1 _18169_ (.A0(\rvcpu.dp.plde.ImmExtE[24] ),
    .A1(\rvcpu.dp.SrcBFW_Mux.y[24] ),
    .S(_05279_),
    .X(_05534_));
 sky130_fd_sc_hd__and2_1 _18170_ (.A(_05533_),
    .B(_05534_),
    .X(_05535_));
 sky130_fd_sc_hd__nor2_1 _18171_ (.A(_05533_),
    .B(_05534_),
    .Y(_05536_));
 sky130_fd_sc_hd__nor2_2 _18172_ (.A(_05535_),
    .B(_05536_),
    .Y(_05537_));
 sky130_fd_sc_hd__o22a_1 _18173_ (.A1(\rvcpu.dp.plem.ALUResultM[27] ),
    .A2(_05293_),
    .B1(_05294_),
    .B2(_13194_),
    .X(_05538_));
 sky130_fd_sc_hd__o21a_1 _18174_ (.A1(\rvcpu.dp.plde.RD1E[27] ),
    .A2(_05291_),
    .B1(_05538_),
    .X(_05539_));
 sky130_fd_sc_hd__mux2_1 _18175_ (.A0(\rvcpu.dp.plde.ImmExtE[27] ),
    .A1(\rvcpu.dp.SrcBFW_Mux.y[27] ),
    .S(_05279_),
    .X(_05540_));
 sky130_fd_sc_hd__nor2_1 _18176_ (.A(_05539_),
    .B(_05540_),
    .Y(_05541_));
 sky130_fd_sc_hd__and2_1 _18177_ (.A(_05539_),
    .B(_05540_),
    .X(_05542_));
 sky130_fd_sc_hd__nor2_2 _18178_ (.A(_05541_),
    .B(_05542_),
    .Y(_05543_));
 sky130_fd_sc_hd__o22a_1 _18179_ (.A1(\rvcpu.dp.plem.ALUResultM[26] ),
    .A2(_05293_),
    .B1(_05294_),
    .B2(_13197_),
    .X(_05544_));
 sky130_fd_sc_hd__o21a_1 _18180_ (.A1(\rvcpu.dp.plde.RD1E[26] ),
    .A2(_05291_),
    .B1(_05544_),
    .X(_05545_));
 sky130_fd_sc_hd__mux2_1 _18181_ (.A0(\rvcpu.dp.plde.ImmExtE[26] ),
    .A1(\rvcpu.dp.SrcBFW_Mux.y[26] ),
    .S(_05279_),
    .X(_05546_));
 sky130_fd_sc_hd__and2_1 _18182_ (.A(_05545_),
    .B(_05546_),
    .X(_05547_));
 sky130_fd_sc_hd__nor2_1 _18183_ (.A(_05545_),
    .B(_05546_),
    .Y(_05548_));
 sky130_fd_sc_hd__nor2_2 _18184_ (.A(_05547_),
    .B(_05548_),
    .Y(_05549_));
 sky130_fd_sc_hd__and4_1 _18185_ (.A(_05531_),
    .B(_05537_),
    .C(_05543_),
    .D(_05549_),
    .X(_05550_));
 sky130_fd_sc_hd__inv_2 _18186_ (.A(_05530_),
    .Y(_05551_));
 sky130_fd_sc_hd__a21o_1 _18187_ (.A1(_05551_),
    .A2(_05535_),
    .B1(_05529_),
    .X(_05552_));
 sky130_fd_sc_hd__a211o_1 _18188_ (.A1(_05549_),
    .A2(_05552_),
    .B1(_05542_),
    .C1(_05547_),
    .X(_05553_));
 sky130_fd_sc_hd__or2_1 _18189_ (.A(_05539_),
    .B(_05540_),
    .X(_05554_));
 sky130_fd_sc_hd__a22oi_2 _18190_ (.A1(_05525_),
    .A2(_05550_),
    .B1(_05553_),
    .B2(_05554_),
    .Y(_05555_));
 sky130_fd_sc_hd__and2_1 _18191_ (.A(_05296_),
    .B(_05297_),
    .X(_05556_));
 sky130_fd_sc_hd__nor2_1 _18192_ (.A(_05302_),
    .B(_05556_),
    .Y(_05557_));
 sky130_fd_sc_hd__o21a_1 _18193_ (.A1(_05305_),
    .A2(_05555_),
    .B1(_05557_),
    .X(_05558_));
 sky130_fd_sc_hd__o31ai_2 _18194_ (.A1(_05290_),
    .A2(_05298_),
    .A3(_05558_),
    .B1(_05288_),
    .Y(_05559_));
 sky130_fd_sc_hd__xnor2_1 _18195_ (.A(_05284_),
    .B(_05559_),
    .Y(_05560_));
 sky130_fd_sc_hd__nor2_2 _18196_ (.A(_05298_),
    .B(_05556_),
    .Y(_05561_));
 sky130_fd_sc_hd__inv_2 _18197_ (.A(_05561_),
    .Y(_05562_));
 sky130_fd_sc_hd__or2b_1 _18198_ (.A(_05486_),
    .B_N(_05487_),
    .X(_05563_));
 sky130_fd_sc_hd__clkbuf_4 _18199_ (.A(_05291_),
    .X(_05564_));
 sky130_fd_sc_hd__o21ai_2 _18200_ (.A1(\rvcpu.dp.plde.RD1E[17] ),
    .A2(_05564_),
    .B1(_05499_),
    .Y(_05565_));
 sky130_fd_sc_hd__inv_2 _18201_ (.A(_05506_),
    .Y(_05566_));
 sky130_fd_sc_hd__or2_1 _18202_ (.A(_05566_),
    .B(_05509_),
    .X(_05567_));
 sky130_fd_sc_hd__or2_1 _18203_ (.A(_05504_),
    .B(_05567_),
    .X(_05568_));
 sky130_fd_sc_hd__o21a_1 _18204_ (.A1(_05565_),
    .A2(_05501_),
    .B1(_05568_),
    .X(_05569_));
 sky130_fd_sc_hd__o21ai_2 _18205_ (.A1(\rvcpu.dp.plde.RD1E[18] ),
    .A2(_05564_),
    .B1(_05489_),
    .Y(_05570_));
 sky130_fd_sc_hd__or2_1 _18206_ (.A(_05570_),
    .B(_05493_),
    .X(_05571_));
 sky130_fd_sc_hd__o21ai_1 _18207_ (.A1(_05497_),
    .A2(_05569_),
    .B1(_05571_),
    .Y(_05572_));
 sky130_fd_sc_hd__nand2_1 _18208_ (.A(_05563_),
    .B(_05572_),
    .Y(_05573_));
 sky130_fd_sc_hd__o21ai_2 _18209_ (.A1(\rvcpu.dp.plde.RD1E[19] ),
    .A2(_05564_),
    .B1(_05483_),
    .Y(_05574_));
 sky130_fd_sc_hd__a21o_1 _18210_ (.A1(_05384_),
    .A2(_05385_),
    .B1(_05388_),
    .X(_05575_));
 sky130_fd_sc_hd__nand2_1 _18211_ (.A(_05390_),
    .B(_05392_),
    .Y(_05576_));
 sky130_fd_sc_hd__a22o_1 _18212_ (.A1(_05575_),
    .A2(_05389_),
    .B1(_05576_),
    .B2(_05394_),
    .X(_05577_));
 sky130_fd_sc_hd__and2_1 _18213_ (.A(_05384_),
    .B(_05385_),
    .X(_05578_));
 sky130_fd_sc_hd__clkbuf_4 _18214_ (.A(_05578_),
    .X(_05579_));
 sky130_fd_sc_hd__a221o_1 _18215_ (.A1(\rvcpu.dp.plde.RD1E[1] ),
    .A2(_05266_),
    .B1(_05270_),
    .B2(_13274_),
    .C1(_05387_),
    .X(_05580_));
 sky130_fd_sc_hd__nand2_1 _18216_ (.A(_05579_),
    .B(_05580_),
    .Y(_05581_));
 sky130_fd_sc_hd__a21oi_1 _18217_ (.A1(_05577_),
    .A2(_05581_),
    .B1(_05383_),
    .Y(_05582_));
 sky130_fd_sc_hd__nor2_1 _18218_ (.A(_05380_),
    .B(_05382_),
    .Y(_05583_));
 sky130_fd_sc_hd__nand2_1 _18219_ (.A(_05374_),
    .B(_05377_),
    .Y(_05584_));
 sky130_fd_sc_hd__o21ai_1 _18220_ (.A1(_05582_),
    .A2(_05583_),
    .B1(_05584_),
    .Y(_05585_));
 sky130_fd_sc_hd__nand2_1 _18221_ (.A(_05375_),
    .B(_05373_),
    .Y(_05586_));
 sky130_fd_sc_hd__inv_2 _18222_ (.A(_05358_),
    .Y(_05587_));
 sky130_fd_sc_hd__xnor2_4 _18223_ (.A(_05587_),
    .B(_05359_),
    .Y(_05588_));
 sky130_fd_sc_hd__a211o_1 _18224_ (.A1(_05585_),
    .A2(_05586_),
    .B1(_05368_),
    .C1(_05588_),
    .X(_05589_));
 sky130_fd_sc_hd__o21a_4 _18225_ (.A1(_05321_),
    .A2(\rvcpu.dp.SrcBFW_Mux.y[4] ),
    .B1(_05362_),
    .X(_05590_));
 sky130_fd_sc_hd__or2_1 _18226_ (.A(_05590_),
    .B(_05365_),
    .X(_05591_));
 sky130_fd_sc_hd__nor2_1 _18227_ (.A(_05587_),
    .B(_05359_),
    .Y(_05592_));
 sky130_fd_sc_hd__o21ba_1 _18228_ (.A1(_05588_),
    .A2(_05591_),
    .B1_N(_05592_),
    .X(_05593_));
 sky130_fd_sc_hd__or2b_1 _18229_ (.A(_05353_),
    .B_N(_05349_),
    .X(_05594_));
 sky130_fd_sc_hd__o21a_1 _18230_ (.A1(_05356_),
    .A2(_05593_),
    .B1(_05594_),
    .X(_05595_));
 sky130_fd_sc_hd__o21ai_2 _18231_ (.A1(\rvcpu.dp.plde.RD1E[7] ),
    .A2(_05292_),
    .B1(_05341_),
    .Y(_05596_));
 sky130_fd_sc_hd__or2_1 _18232_ (.A(_05596_),
    .B(_05343_),
    .X(_05597_));
 sky130_fd_sc_hd__o21a_1 _18233_ (.A1(_05346_),
    .A2(_05595_),
    .B1(_05597_),
    .X(_05598_));
 sky130_fd_sc_hd__o31ai_4 _18234_ (.A1(_05346_),
    .A2(_05356_),
    .A3(_05589_),
    .B1(_05598_),
    .Y(_05599_));
 sky130_fd_sc_hd__or4_1 _18235_ (.A(_05311_),
    .B(_05318_),
    .C(_05436_),
    .D(_05438_),
    .X(_05600_));
 sky130_fd_sc_hd__nor2_1 _18236_ (.A(_05427_),
    .B(_05431_),
    .Y(_05601_));
 sky130_fd_sc_hd__nor4b_1 _18237_ (.A(_05410_),
    .B(_05600_),
    .C(_05419_),
    .D_N(_05601_),
    .Y(_05602_));
 sky130_fd_sc_hd__a221oi_4 _18238_ (.A1(\rvcpu.dp.plde.RD1E[15] ),
    .A2(_05266_),
    .B1(_05271_),
    .B2(_13231_),
    .C1(_05312_),
    .Y(_05603_));
 sky130_fd_sc_hd__a221oi_4 _18239_ (.A1(\rvcpu.dp.plem.ALUResultM[8] ),
    .A2(_05272_),
    .B1(_05267_),
    .B2(\rvcpu.dp.plde.RD1E[8] ),
    .C1(_05420_),
    .Y(_05604_));
 sky130_fd_sc_hd__o32a_1 _18240_ (.A1(_05604_),
    .A2(_05424_),
    .A3(_05431_),
    .B1(_05430_),
    .B2(net102),
    .X(_05605_));
 sky130_fd_sc_hd__a221oi_4 _18241_ (.A1(\rvcpu.dp.plde.RD1E[10] ),
    .A2(_05267_),
    .B1(_05271_),
    .B2(_13247_),
    .C1(_05411_),
    .Y(_05606_));
 sky130_fd_sc_hd__or2_1 _18242_ (.A(_05606_),
    .B(_05415_),
    .X(_05607_));
 sky130_fd_sc_hd__o22a_1 _18243_ (.A1(net103),
    .A2(_05409_),
    .B1(_05410_),
    .B2(_05607_),
    .X(_05608_));
 sky130_fd_sc_hd__o31a_1 _18244_ (.A1(_05410_),
    .A2(_05418_),
    .A3(_05605_),
    .B1(_05608_),
    .X(_05609_));
 sky130_fd_sc_hd__inv_2 _18245_ (.A(_05327_),
    .Y(_05610_));
 sky130_fd_sc_hd__o32a_1 _18246_ (.A1(_05610_),
    .A2(_05330_),
    .A3(_05438_),
    .B1(_05323_),
    .B2(_05437_),
    .X(_05611_));
 sky130_fd_sc_hd__or2_1 _18247_ (.A(net105),
    .B(_05310_),
    .X(_05612_));
 sky130_fd_sc_hd__o21a_1 _18248_ (.A1(_05311_),
    .A2(_05611_),
    .B1(_05612_),
    .X(_05613_));
 sky130_fd_sc_hd__or2_1 _18249_ (.A(_05318_),
    .B(_05613_),
    .X(_05614_));
 sky130_fd_sc_hd__o221a_1 _18250_ (.A1(_05603_),
    .A2(_05314_),
    .B1(_05600_),
    .B2(_05609_),
    .C1(_05614_),
    .X(_05615_));
 sky130_fd_sc_hd__a21boi_2 _18251_ (.A1(_05599_),
    .A2(_05602_),
    .B1_N(_05615_),
    .Y(_05616_));
 sky130_fd_sc_hd__or4_1 _18252_ (.A(_05488_),
    .B(_05497_),
    .C(_05504_),
    .D(_05512_),
    .X(_05617_));
 sky130_fd_sc_hd__o22a_1 _18253_ (.A1(_05574_),
    .A2(_05485_),
    .B1(_05616_),
    .B2(_05617_),
    .X(_05618_));
 sky130_fd_sc_hd__a21oi_2 _18254_ (.A1(_05573_),
    .A2(_05618_),
    .B1(_05481_),
    .Y(_05619_));
 sky130_fd_sc_hd__nor3_1 _18255_ (.A(_05461_),
    .B(_05467_),
    .C(_05473_),
    .Y(_05620_));
 sky130_fd_sc_hd__o21ai_2 _18256_ (.A1(\rvcpu.dp.plde.RD1E[21] ),
    .A2(_05564_),
    .B1(_05468_),
    .Y(_05621_));
 sky130_fd_sc_hd__o21ai_2 _18257_ (.A1(\rvcpu.dp.plde.RD1E[20] ),
    .A2(_05564_),
    .B1(_05474_),
    .Y(_05622_));
 sky130_fd_sc_hd__or3_1 _18258_ (.A(_05473_),
    .B(_05622_),
    .C(_05478_),
    .X(_05623_));
 sky130_fd_sc_hd__o21a_1 _18259_ (.A1(_05621_),
    .A2(_05470_),
    .B1(_05623_),
    .X(_05624_));
 sky130_fd_sc_hd__o21ai_2 _18260_ (.A1(\rvcpu.dp.plde.RD1E[23] ),
    .A2(_05564_),
    .B1(_05455_),
    .Y(_05625_));
 sky130_fd_sc_hd__o21ai_2 _18261_ (.A1(\rvcpu.dp.plde.RD1E[22] ),
    .A2(_05564_),
    .B1(_05462_),
    .Y(_05626_));
 sky130_fd_sc_hd__or2_1 _18262_ (.A(_05626_),
    .B(_05464_),
    .X(_05627_));
 sky130_fd_sc_hd__o22a_1 _18263_ (.A1(_05625_),
    .A2(_05457_),
    .B1(_05461_),
    .B2(_05627_),
    .X(_05628_));
 sky130_fd_sc_hd__o31ai_2 _18264_ (.A1(_05461_),
    .A2(_05467_),
    .A3(_05624_),
    .B1(_05628_),
    .Y(_05629_));
 sky130_fd_sc_hd__a21o_1 _18265_ (.A1(_05619_),
    .A2(_05620_),
    .B1(_05629_),
    .X(_05630_));
 sky130_fd_sc_hd__nor4_1 _18266_ (.A(_05531_),
    .B(_05537_),
    .C(_05543_),
    .D(_05549_),
    .Y(_05631_));
 sky130_fd_sc_hd__o21ai_1 _18267_ (.A1(\rvcpu.dp.plde.RD1E[25] ),
    .A2(_05564_),
    .B1(_05526_),
    .Y(_05632_));
 sky130_fd_sc_hd__o21ai_2 _18268_ (.A1(\rvcpu.dp.plde.RD1E[24] ),
    .A2(_05291_),
    .B1(_05532_),
    .Y(_05633_));
 sky130_fd_sc_hd__or3_1 _18269_ (.A(_05531_),
    .B(_05633_),
    .C(_05534_),
    .X(_05634_));
 sky130_fd_sc_hd__o21a_1 _18270_ (.A1(_05632_),
    .A2(_05528_),
    .B1(_05634_),
    .X(_05635_));
 sky130_fd_sc_hd__o21ai_1 _18271_ (.A1(\rvcpu.dp.plde.RD1E[27] ),
    .A2(_05564_),
    .B1(_05538_),
    .Y(_05636_));
 sky130_fd_sc_hd__o21ai_1 _18272_ (.A1(\rvcpu.dp.plde.RD1E[26] ),
    .A2(_05564_),
    .B1(_05544_),
    .Y(_05637_));
 sky130_fd_sc_hd__or2_1 _18273_ (.A(_05637_),
    .B(_05546_),
    .X(_05638_));
 sky130_fd_sc_hd__o22a_1 _18274_ (.A1(_05636_),
    .A2(_05540_),
    .B1(_05543_),
    .B2(_05638_),
    .X(_05639_));
 sky130_fd_sc_hd__o31ai_1 _18275_ (.A1(_05543_),
    .A2(_05549_),
    .A3(_05635_),
    .B1(_05639_),
    .Y(_05640_));
 sky130_fd_sc_hd__a21o_1 _18276_ (.A1(_05630_),
    .A2(_05631_),
    .B1(_05640_),
    .X(_05641_));
 sky130_fd_sc_hd__o21ai_2 _18277_ (.A1(\rvcpu.dp.plde.RD1E[29] ),
    .A2(_05291_),
    .B1(_05295_),
    .Y(_05642_));
 sky130_fd_sc_hd__inv_2 _18278_ (.A(_05300_),
    .Y(_05643_));
 sky130_fd_sc_hd__or2_1 _18279_ (.A(_05643_),
    .B(_05301_),
    .X(_05644_));
 sky130_fd_sc_hd__or2_1 _18280_ (.A(_05561_),
    .B(_05644_),
    .X(_05645_));
 sky130_fd_sc_hd__o21ai_1 _18281_ (.A1(_05642_),
    .A2(_05297_),
    .B1(_05645_),
    .Y(_05646_));
 sky130_fd_sc_hd__a31o_1 _18282_ (.A1(_05305_),
    .A2(_05562_),
    .A3(_05641_),
    .B1(_05646_),
    .X(_05647_));
 sky130_fd_sc_hd__inv_2 _18283_ (.A(_05286_),
    .Y(_05648_));
 sky130_fd_sc_hd__or2_1 _18284_ (.A(_05648_),
    .B(_05287_),
    .X(_05649_));
 sky130_fd_sc_hd__nand2_1 _18285_ (.A(_05283_),
    .B(_05649_),
    .Y(_05650_));
 sky130_fd_sc_hd__a21oi_1 _18286_ (.A1(_05290_),
    .A2(_05647_),
    .B1(_05650_),
    .Y(_05651_));
 sky130_fd_sc_hd__inv_2 _18287_ (.A(\rvcpu.dp.plde.ALUControlE[0] ),
    .Y(_05652_));
 sky130_fd_sc_hd__or2_1 _18288_ (.A(_05652_),
    .B(_00003_),
    .X(_05653_));
 sky130_fd_sc_hd__buf_2 _18289_ (.A(_05653_),
    .X(_05654_));
 sky130_fd_sc_hd__clkbuf_4 _18290_ (.A(_05654_),
    .X(_05655_));
 sky130_fd_sc_hd__nor2_1 _18291_ (.A(_05283_),
    .B(_05649_),
    .Y(_05656_));
 sky130_fd_sc_hd__a311o_1 _18292_ (.A1(_05284_),
    .A2(_05290_),
    .A3(_05647_),
    .B1(_05655_),
    .C1(_05656_),
    .X(_05657_));
 sky130_fd_sc_hd__clkbuf_4 _18293_ (.A(_05363_),
    .X(_05658_));
 sky130_fd_sc_hd__nand2_1 _18294_ (.A(\rvcpu.dp.plde.ALUControlE[0] ),
    .B(\rvcpu.dp.plde.ALUControlE[1] ),
    .Y(_05659_));
 sky130_fd_sc_hd__or3b_4 _18295_ (.A(\rvcpu.dp.plde.ALUControlE[2] ),
    .B(_05659_),
    .C_N(\rvcpu.dp.plde.ALUControlE[3] ),
    .X(_05660_));
 sky130_fd_sc_hd__nor2_2 _18296_ (.A(_05658_),
    .B(_05660_),
    .Y(_05661_));
 sky130_fd_sc_hd__clkbuf_4 _18297_ (.A(_05576_),
    .X(_05662_));
 sky130_fd_sc_hd__clkbuf_4 _18298_ (.A(_05662_),
    .X(_05663_));
 sky130_fd_sc_hd__clkbuf_4 _18299_ (.A(_05663_),
    .X(_05664_));
 sky130_fd_sc_hd__clkbuf_4 _18300_ (.A(_05664_),
    .X(_05665_));
 sky130_fd_sc_hd__clkbuf_4 _18301_ (.A(_05665_),
    .X(_05666_));
 sky130_fd_sc_hd__nand2_2 _18302_ (.A(_05384_),
    .B(_05385_),
    .Y(_05667_));
 sky130_fd_sc_hd__clkbuf_4 _18303_ (.A(_05667_),
    .X(_05668_));
 sky130_fd_sc_hd__clkbuf_4 _18304_ (.A(_05668_),
    .X(_05669_));
 sky130_fd_sc_hd__clkbuf_4 _18305_ (.A(_05669_),
    .X(_05670_));
 sky130_fd_sc_hd__clkbuf_4 _18306_ (.A(_05670_),
    .X(_05671_));
 sky130_fd_sc_hd__mux4_1 _18307_ (.A0(_05313_),
    .A1(_05334_),
    .A2(_05320_),
    .A3(_05327_),
    .S0(_05666_),
    .S1(_05671_),
    .X(_05672_));
 sky130_fd_sc_hd__mux4_1 _18308_ (.A0(_05446_),
    .A1(_05412_),
    .A2(_05441_),
    .A3(_05421_),
    .S0(_05665_),
    .S1(_05670_),
    .X(_05673_));
 sky130_fd_sc_hd__buf_2 _18309_ (.A(_05380_),
    .X(_05674_));
 sky130_fd_sc_hd__buf_2 _18310_ (.A(_05674_),
    .X(_05675_));
 sky130_fd_sc_hd__clkbuf_4 _18311_ (.A(_05675_),
    .X(_05676_));
 sky130_fd_sc_hd__clkbuf_4 _18312_ (.A(_05676_),
    .X(_05677_));
 sky130_fd_sc_hd__mux2_1 _18313_ (.A0(_05672_),
    .A1(_05673_),
    .S(_05677_),
    .X(_05678_));
 sky130_fd_sc_hd__inv_2 _18314_ (.A(_05365_),
    .Y(_05679_));
 sky130_fd_sc_hd__mux4_2 _18315_ (.A0(_05342_),
    .A1(_05349_),
    .A2(_05358_),
    .A3(_05679_),
    .S0(_05664_),
    .S1(_05669_),
    .X(_05680_));
 sky130_fd_sc_hd__and2_1 _18316_ (.A(_05390_),
    .B(_05392_),
    .X(_05681_));
 sky130_fd_sc_hd__buf_2 _18317_ (.A(_05681_),
    .X(_05682_));
 sky130_fd_sc_hd__clkbuf_4 _18318_ (.A(_05682_),
    .X(_05683_));
 sky130_fd_sc_hd__clkbuf_4 _18319_ (.A(_05683_),
    .X(_05684_));
 sky130_fd_sc_hd__a21o_1 _18320_ (.A1(_05580_),
    .A2(_05684_),
    .B1(_05395_),
    .X(_05685_));
 sky130_fd_sc_hd__nand2_1 _18321_ (.A(_05382_),
    .B(_05662_),
    .Y(_05686_));
 sky130_fd_sc_hd__o21a_1 _18322_ (.A1(_05373_),
    .A2(_05663_),
    .B1(_05686_),
    .X(_05687_));
 sky130_fd_sc_hd__clkbuf_4 _18323_ (.A(_05579_),
    .X(_05688_));
 sky130_fd_sc_hd__clkbuf_4 _18324_ (.A(_05688_),
    .X(_05689_));
 sky130_fd_sc_hd__mux2_1 _18325_ (.A0(_05685_),
    .A1(_05687_),
    .S(_05689_),
    .X(_05690_));
 sky130_fd_sc_hd__mux2_2 _18326_ (.A0(_05680_),
    .A1(_05690_),
    .S(_05676_),
    .X(_05691_));
 sky130_fd_sc_hd__buf_2 _18327_ (.A(_05370_),
    .X(_05692_));
 sky130_fd_sc_hd__buf_2 _18328_ (.A(_05692_),
    .X(_05693_));
 sky130_fd_sc_hd__buf_2 _18329_ (.A(_05693_),
    .X(_05694_));
 sky130_fd_sc_hd__mux2_1 _18330_ (.A0(_05678_),
    .A1(_05691_),
    .S(_05694_),
    .X(_05695_));
 sky130_fd_sc_hd__clkbuf_4 _18331_ (.A(_05375_),
    .X(_05696_));
 sky130_fd_sc_hd__clkbuf_4 _18332_ (.A(_05696_),
    .X(_05697_));
 sky130_fd_sc_hd__buf_2 _18333_ (.A(_05697_),
    .X(_05698_));
 sky130_fd_sc_hd__mux4_1 _18334_ (.A0(_05456_),
    .A1(_05463_),
    .A2(_05469_),
    .A3(_05475_),
    .S0(_05666_),
    .S1(_05671_),
    .X(_05699_));
 sky130_fd_sc_hd__mux4_1 _18335_ (.A0(_05484_),
    .A1(_05490_),
    .A2(_05500_),
    .A3(_05506_),
    .S0(_05666_),
    .S1(_05671_),
    .X(_05700_));
 sky130_fd_sc_hd__mux2_1 _18336_ (.A0(_05699_),
    .A1(_05700_),
    .S(_05677_),
    .X(_05701_));
 sky130_fd_sc_hd__nor2_4 _18337_ (.A(_05590_),
    .B(_05660_),
    .Y(_05702_));
 sky130_fd_sc_hd__buf_2 _18338_ (.A(_05702_),
    .X(_05703_));
 sky130_fd_sc_hd__buf_2 _18339_ (.A(_05398_),
    .X(_05704_));
 sky130_fd_sc_hd__clkbuf_4 _18340_ (.A(_05704_),
    .X(_05705_));
 sky130_fd_sc_hd__buf_2 _18341_ (.A(_05705_),
    .X(_05706_));
 sky130_fd_sc_hd__clkbuf_4 _18342_ (.A(_05706_),
    .X(_05707_));
 sky130_fd_sc_hd__mux2_1 _18343_ (.A0(_05296_),
    .A1(_05300_),
    .S(_05665_),
    .X(_05708_));
 sky130_fd_sc_hd__nand2_2 _18344_ (.A(_05688_),
    .B(_05663_),
    .Y(_05709_));
 sky130_fd_sc_hd__inv_2 _18345_ (.A(_05709_),
    .Y(_05710_));
 sky130_fd_sc_hd__and3_1 _18346_ (.A(_05274_),
    .B(_05688_),
    .C(_05684_),
    .X(_05711_));
 sky130_fd_sc_hd__a221o_1 _18347_ (.A1(_05671_),
    .A2(_05708_),
    .B1(_05710_),
    .B2(_05286_),
    .C1(_05711_),
    .X(_05712_));
 sky130_fd_sc_hd__mux2_1 _18348_ (.A0(_05539_),
    .A1(_05545_),
    .S(_05666_),
    .X(_05713_));
 sky130_fd_sc_hd__mux2_1 _18349_ (.A0(_05527_),
    .A1(_05533_),
    .S(_05665_),
    .X(_05714_));
 sky130_fd_sc_hd__mux2_1 _18350_ (.A0(_05713_),
    .A1(_05714_),
    .S(_05671_),
    .X(_05715_));
 sky130_fd_sc_hd__a21o_1 _18351_ (.A1(_05677_),
    .A2(_05715_),
    .B1(_05694_),
    .X(_05716_));
 sky130_fd_sc_hd__a21o_1 _18352_ (.A1(_05707_),
    .A2(_05712_),
    .B1(_05716_),
    .X(_05717_));
 sky130_fd_sc_hd__o211a_1 _18353_ (.A1(_05698_),
    .A2(_05701_),
    .B1(_05703_),
    .C1(_05717_),
    .X(_05718_));
 sky130_fd_sc_hd__or3_2 _18354_ (.A(_05380_),
    .B(_05668_),
    .C(_05662_),
    .X(_05719_));
 sky130_fd_sc_hd__nand2_2 _18355_ (.A(_05363_),
    .B(_05375_),
    .Y(_05720_));
 sky130_fd_sc_hd__nor2_1 _18356_ (.A(_05719_),
    .B(_05720_),
    .Y(_05721_));
 sky130_fd_sc_hd__or2b_1 _18357_ (.A(\rvcpu.dp.plde.ALUControlE[3] ),
    .B_N(\rvcpu.dp.plde.ALUControlE[2] ),
    .X(_05722_));
 sky130_fd_sc_hd__or3b_1 _18358_ (.A(\rvcpu.dp.plde.ALUControlE[0] ),
    .B(\rvcpu.dp.plde.ALUControlE[2] ),
    .C_N(\rvcpu.dp.plde.ALUControlE[3] ),
    .X(_05723_));
 sky130_fd_sc_hd__o21ai_2 _18359_ (.A1(_05659_),
    .A2(_05722_),
    .B1(_05723_),
    .Y(_05724_));
 sky130_fd_sc_hd__and3b_1 _18360_ (.A_N(_05722_),
    .B(_05652_),
    .C(\rvcpu.dp.plde.ALUControlE[1] ),
    .X(_05725_));
 sky130_fd_sc_hd__buf_2 _18361_ (.A(_05725_),
    .X(_05726_));
 sky130_fd_sc_hd__clkbuf_4 _18362_ (.A(_05726_),
    .X(_05727_));
 sky130_fd_sc_hd__clkbuf_4 _18363_ (.A(_05727_),
    .X(_05728_));
 sky130_fd_sc_hd__nor2_2 _18364_ (.A(_05236_),
    .B(_05659_),
    .Y(_05729_));
 sky130_fd_sc_hd__buf_2 _18365_ (.A(_05729_),
    .X(_05730_));
 sky130_fd_sc_hd__or3b_1 _18366_ (.A(_05236_),
    .B(\rvcpu.dp.plde.ALUControlE[0] ),
    .C_N(\rvcpu.dp.plde.ALUControlE[1] ),
    .X(_05731_));
 sky130_fd_sc_hd__clkbuf_4 _18367_ (.A(_05731_),
    .X(_05732_));
 sky130_fd_sc_hd__and4_2 _18368_ (.A(\rvcpu.dp.plde.ALUControlE[0] ),
    .B(\rvcpu.dp.plde.ALUControlE[1] ),
    .C(\rvcpu.dp.plde.ALUControlE[3] ),
    .D(\rvcpu.dp.plde.ALUControlE[2] ),
    .X(_05733_));
 sky130_fd_sc_hd__nand2_1 _18369_ (.A(_05275_),
    .B(_05733_),
    .Y(_05734_));
 sky130_fd_sc_hd__o21ai_1 _18370_ (.A1(_05282_),
    .A2(_05732_),
    .B1(_05734_),
    .Y(_05735_));
 sky130_fd_sc_hd__a221o_1 _18371_ (.A1(_05283_),
    .A2(_05728_),
    .B1(_05730_),
    .B2(_05281_),
    .C1(_05735_),
    .X(_05736_));
 sky130_fd_sc_hd__a31o_1 _18372_ (.A1(_05275_),
    .A2(_05721_),
    .A3(_05724_),
    .B1(_05736_),
    .X(_05737_));
 sky130_fd_sc_hd__a211o_1 _18373_ (.A1(_05661_),
    .A2(_05695_),
    .B1(_05718_),
    .C1(_05737_),
    .X(_05738_));
 sky130_fd_sc_hd__o21bai_1 _18374_ (.A1(_05651_),
    .A2(_05657_),
    .B1_N(_05738_),
    .Y(_05739_));
 sky130_fd_sc_hd__a21o_1 _18375_ (.A1(_05240_),
    .A2(_05560_),
    .B1(_05739_),
    .X(_05740_));
 sky130_fd_sc_hd__buf_1 _18376_ (.A(_05740_),
    .X(\rvcpu.ALUResultE[31] ));
 sky130_fd_sc_hd__a221oi_4 _18377_ (.A1(\rvcpu.dp.plde.RD1E[31] ),
    .A2(_05266_),
    .B1(_05270_),
    .B2(_13172_),
    .C1(_05273_),
    .Y(_05741_));
 sky130_fd_sc_hd__nor2_1 _18378_ (.A(_05741_),
    .B(_05280_),
    .Y(_05742_));
 sky130_fd_sc_hd__a311o_1 _18379_ (.A1(_05284_),
    .A2(_05290_),
    .A3(_05647_),
    .B1(_05656_),
    .C1(_05742_),
    .X(_05743_));
 sky130_fd_sc_hd__or2_1 _18380_ (.A(\rvcpu.dp.plde.unsignE ),
    .B(_05284_),
    .X(_05744_));
 sky130_fd_sc_hd__or2_1 _18381_ (.A(_05742_),
    .B(_05744_),
    .X(_05745_));
 sky130_fd_sc_hd__or4b_1 _18382_ (.A(_05652_),
    .B(\rvcpu.dp.plde.ALUControlE[1] ),
    .C(_05722_),
    .D_N(_05745_),
    .X(_05746_));
 sky130_fd_sc_hd__a21oi_1 _18383_ (.A1(_05743_),
    .A2(_05744_),
    .B1(_05746_),
    .Y(_05747_));
 sky130_fd_sc_hd__or2_1 _18384_ (.A(_05724_),
    .B(_05733_),
    .X(_05748_));
 sky130_fd_sc_hd__clkbuf_4 _18385_ (.A(_05748_),
    .X(_05749_));
 sky130_fd_sc_hd__nand2_2 _18386_ (.A(_05590_),
    .B(_05749_),
    .Y(_05750_));
 sky130_fd_sc_hd__mux4_1 _18387_ (.A0(_05574_),
    .A1(_05570_),
    .A2(_05565_),
    .A3(_05566_),
    .S0(_05683_),
    .S1(_05579_),
    .X(_05751_));
 sky130_fd_sc_hd__mux4_1 _18388_ (.A0(_05456_),
    .A1(_05463_),
    .A2(_05469_),
    .A3(_05475_),
    .S0(_05683_),
    .S1(_05688_),
    .X(_05752_));
 sky130_fd_sc_hd__inv_2 _18389_ (.A(_05752_),
    .Y(_05753_));
 sky130_fd_sc_hd__mux2_1 _18390_ (.A0(_05751_),
    .A1(_05753_),
    .S(_05676_),
    .X(_05754_));
 sky130_fd_sc_hd__nand2_1 _18391_ (.A(_05642_),
    .B(_05662_),
    .Y(_05755_));
 sky130_fd_sc_hd__o21ai_1 _18392_ (.A1(_05300_),
    .A2(_05663_),
    .B1(_05755_),
    .Y(_05756_));
 sky130_fd_sc_hd__nor2_1 _18393_ (.A(_05286_),
    .B(_05662_),
    .Y(_05757_));
 sky130_fd_sc_hd__a21o_1 _18394_ (.A1(_05741_),
    .A2(_05662_),
    .B1(_05757_),
    .X(_05758_));
 sky130_fd_sc_hd__mux2_1 _18395_ (.A0(_05756_),
    .A1(_05758_),
    .S(_05668_),
    .X(_05759_));
 sky130_fd_sc_hd__mux2_1 _18396_ (.A0(_05527_),
    .A1(_05533_),
    .S(_05683_),
    .X(_05760_));
 sky130_fd_sc_hd__mux2_1 _18397_ (.A0(_05539_),
    .A1(_05545_),
    .S(_05682_),
    .X(_05761_));
 sky130_fd_sc_hd__mux2_1 _18398_ (.A0(_05760_),
    .A1(_05761_),
    .S(_05668_),
    .X(_05762_));
 sky130_fd_sc_hd__nand2_1 _18399_ (.A(_05705_),
    .B(_05762_),
    .Y(_05763_));
 sky130_fd_sc_hd__o21a_1 _18400_ (.A1(_05705_),
    .A2(_05759_),
    .B1(_05763_),
    .X(_05764_));
 sky130_fd_sc_hd__mux2_1 _18401_ (.A0(_05754_),
    .A1(_05764_),
    .S(_05693_),
    .X(_05765_));
 sky130_fd_sc_hd__mux4_1 _18402_ (.A0(_05342_),
    .A1(_05349_),
    .A2(_05358_),
    .A3(_05679_),
    .S0(_05683_),
    .S1(_05688_),
    .X(_05766_));
 sky130_fd_sc_hd__inv_2 _18403_ (.A(_05766_),
    .Y(_05767_));
 sky130_fd_sc_hd__clkbuf_4 _18404_ (.A(_05689_),
    .X(_05768_));
 sky130_fd_sc_hd__clkbuf_4 _18405_ (.A(_05683_),
    .X(_05769_));
 sky130_fd_sc_hd__mux2_1 _18406_ (.A0(_05376_),
    .A1(_05382_),
    .S(_05769_),
    .X(_05770_));
 sky130_fd_sc_hd__a221o_2 _18407_ (.A1(\rvcpu.dp.plde.RD1E[0] ),
    .A2(_05266_),
    .B1(_05270_),
    .B2(_13277_),
    .C1(_05393_),
    .X(_05771_));
 sky130_fd_sc_hd__nor2_1 _18408_ (.A(_05666_),
    .B(_05771_),
    .Y(_05772_));
 sky130_fd_sc_hd__a211o_1 _18409_ (.A1(_05388_),
    .A2(_05666_),
    .B1(_05772_),
    .C1(_05671_),
    .X(_05773_));
 sky130_fd_sc_hd__o211a_1 _18410_ (.A1(_05768_),
    .A2(_05770_),
    .B1(_05773_),
    .C1(_05707_),
    .X(_05774_));
 sky130_fd_sc_hd__nor2_4 _18411_ (.A(_05590_),
    .B(_05370_),
    .Y(_05775_));
 sky130_fd_sc_hd__nand2_4 _18412_ (.A(_05775_),
    .B(_05749_),
    .Y(_05776_));
 sky130_fd_sc_hd__a211o_1 _18413_ (.A1(_05677_),
    .A2(_05767_),
    .B1(_05774_),
    .C1(_05776_),
    .X(_05777_));
 sky130_fd_sc_hd__mux4_1 _18414_ (.A0(_05408_),
    .A1(_05606_),
    .A2(net102),
    .A3(_05604_),
    .S0(_05684_),
    .S1(_05689_),
    .X(_05778_));
 sky130_fd_sc_hd__mux4_1 _18415_ (.A0(_05603_),
    .A1(_05307_),
    .A2(_05437_),
    .A3(_05610_),
    .S0(_05683_),
    .S1(_05579_),
    .X(_05779_));
 sky130_fd_sc_hd__mux2_1 _18416_ (.A0(_05778_),
    .A1(_05779_),
    .S(_05677_),
    .X(_05780_));
 sky130_fd_sc_hd__nor2_2 _18417_ (.A(_05590_),
    .B(_05375_),
    .Y(_05781_));
 sky130_fd_sc_hd__nand2_2 _18418_ (.A(_05749_),
    .B(_05781_),
    .Y(_05782_));
 sky130_fd_sc_hd__or2_1 _18419_ (.A(_05236_),
    .B(_05659_),
    .X(_05783_));
 sky130_fd_sc_hd__buf_2 _18420_ (.A(_05783_),
    .X(_05784_));
 sky130_fd_sc_hd__buf_2 _18421_ (.A(_05784_),
    .X(_05785_));
 sky130_fd_sc_hd__or3b_4 _18422_ (.A(_05722_),
    .B(\rvcpu.dp.plde.ALUControlE[0] ),
    .C_N(\rvcpu.dp.plde.ALUControlE[1] ),
    .X(_05786_));
 sky130_fd_sc_hd__a21o_1 _18423_ (.A1(_00003_),
    .A2(_05786_),
    .B1(_05395_),
    .X(_05787_));
 sky130_fd_sc_hd__a21o_1 _18424_ (.A1(_05785_),
    .A2(_05787_),
    .B1(_05772_),
    .X(_05788_));
 sky130_fd_sc_hd__and4b_1 _18425_ (.A_N(\rvcpu.dp.plde.ALUControlE[2] ),
    .B(\rvcpu.dp.plde.ALUControlE[3] ),
    .C(\rvcpu.dp.plde.ALUControlE[1] ),
    .D(\rvcpu.dp.plde.ALUControlE[0] ),
    .X(_05789_));
 sky130_fd_sc_hd__nand2_1 _18426_ (.A(_05789_),
    .B(_05775_),
    .Y(_05790_));
 sky130_fd_sc_hd__nand2_1 _18427_ (.A(_05576_),
    .B(_05771_),
    .Y(_05791_));
 sky130_fd_sc_hd__o32a_1 _18428_ (.A1(_05394_),
    .A2(_05719_),
    .A3(_05790_),
    .B1(_05732_),
    .B2(_05791_),
    .X(_05792_));
 sky130_fd_sc_hd__o211a_1 _18429_ (.A1(_05780_),
    .A2(_05782_),
    .B1(_05788_),
    .C1(_05792_),
    .X(_05793_));
 sky130_fd_sc_hd__o211ai_2 _18430_ (.A1(_05750_),
    .A2(_05765_),
    .B1(_05777_),
    .C1(_05793_),
    .Y(_05794_));
 sky130_fd_sc_hd__or2_1 _18431_ (.A(_05747_),
    .B(_05794_),
    .X(_05795_));
 sky130_fd_sc_hd__buf_1 _18432_ (.A(_05795_),
    .X(\rvcpu.ALUResultE[0] ));
 sky130_fd_sc_hd__nand2_1 _18433_ (.A(_05689_),
    .B(_05685_),
    .Y(_05796_));
 sky130_fd_sc_hd__or2_1 _18434_ (.A(_05674_),
    .B(_05796_),
    .X(_05797_));
 sky130_fd_sc_hd__inv_2 _18435_ (.A(_05797_),
    .Y(_05798_));
 sky130_fd_sc_hd__clkbuf_4 _18436_ (.A(_05704_),
    .X(_05799_));
 sky130_fd_sc_hd__mux4_1 _18437_ (.A0(_05421_),
    .A1(_05342_),
    .A2(_05349_),
    .A3(_05358_),
    .S0(_05769_),
    .S1(_05689_),
    .X(_05800_));
 sky130_fd_sc_hd__nand2_1 _18438_ (.A(_05581_),
    .B(_05709_),
    .Y(_05801_));
 sky130_fd_sc_hd__nand2_1 _18439_ (.A(_05365_),
    .B(_05662_),
    .Y(_05802_));
 sky130_fd_sc_hd__o21a_1 _18440_ (.A1(_05373_),
    .A2(_05663_),
    .B1(_05802_),
    .X(_05803_));
 sky130_fd_sc_hd__a221o_1 _18441_ (.A1(_05686_),
    .A2(_05801_),
    .B1(_05803_),
    .B2(_05669_),
    .C1(_05675_),
    .X(_05804_));
 sky130_fd_sc_hd__nor2_2 _18442_ (.A(_05724_),
    .B(_05733_),
    .Y(_05805_));
 sky130_fd_sc_hd__nor2_1 _18443_ (.A(_05720_),
    .B(_05805_),
    .Y(_05806_));
 sky130_fd_sc_hd__o211a_1 _18444_ (.A1(_05799_),
    .A2(_05800_),
    .B1(_05804_),
    .C1(_05806_),
    .X(_05807_));
 sky130_fd_sc_hd__and3b_2 _18445_ (.A_N(_05236_),
    .B(_05652_),
    .C(\rvcpu.dp.plde.ALUControlE[1] ),
    .X(_05808_));
 sky130_fd_sc_hd__nor2_4 _18446_ (.A(_05652_),
    .B(_00003_),
    .Y(_05809_));
 sky130_fd_sc_hd__nand2_1 _18447_ (.A(_05575_),
    .B(_05389_),
    .Y(_05810_));
 sky130_fd_sc_hd__or3_1 _18448_ (.A(_05810_),
    .B(_05684_),
    .C(_05771_),
    .X(_05811_));
 sky130_fd_sc_hd__or2_1 _18449_ (.A(\rvcpu.dp.plde.ALUControlE[0] ),
    .B(_00003_),
    .X(_05812_));
 sky130_fd_sc_hd__a21oi_1 _18450_ (.A1(_05810_),
    .A2(_05791_),
    .B1(_05812_),
    .Y(_05813_));
 sky130_fd_sc_hd__or2_1 _18451_ (.A(_05810_),
    .B(_05791_),
    .X(_05814_));
 sky130_fd_sc_hd__a2bb2o_1 _18452_ (.A1_N(_05810_),
    .A2_N(_05786_),
    .B1(_05813_),
    .B2(_05814_),
    .X(_05815_));
 sky130_fd_sc_hd__a31o_1 _18453_ (.A1(_05577_),
    .A2(_05809_),
    .A3(_05811_),
    .B1(_05815_),
    .X(_05816_));
 sky130_fd_sc_hd__a221o_1 _18454_ (.A1(_05389_),
    .A2(_05729_),
    .B1(_05808_),
    .B2(_05396_),
    .C1(_05816_),
    .X(_05817_));
 sky130_fd_sc_hd__a311o_1 _18455_ (.A1(_05696_),
    .A2(_05702_),
    .A3(_05798_),
    .B1(_05807_),
    .C1(_05817_),
    .X(_05818_));
 sky130_fd_sc_hd__o41a_2 _18456_ (.A1(_05370_),
    .A2(_05380_),
    .A3(_05667_),
    .A4(_05576_),
    .B1(_05590_),
    .X(_05819_));
 sky130_fd_sc_hd__and3_2 _18457_ (.A(_05274_),
    .B(_05733_),
    .C(_05819_),
    .X(_05820_));
 sky130_fd_sc_hd__and3_1 _18458_ (.A(_05370_),
    .B(_05674_),
    .C(_05820_),
    .X(_05821_));
 sky130_fd_sc_hd__mux4_1 _18459_ (.A0(_05622_),
    .A1(_05574_),
    .A2(_05570_),
    .A3(_05565_),
    .S0(_05682_),
    .S1(_05579_),
    .X(_05822_));
 sky130_fd_sc_hd__mux4_1 _18460_ (.A0(_05625_),
    .A1(_05621_),
    .A2(_05633_),
    .A3(_05626_),
    .S0(_05579_),
    .S1(_05662_),
    .X(_05823_));
 sky130_fd_sc_hd__mux2_1 _18461_ (.A0(_05822_),
    .A1(_05823_),
    .S(_05674_),
    .X(_05824_));
 sky130_fd_sc_hd__mux4_1 _18462_ (.A0(_05643_),
    .A1(_05636_),
    .A2(_05637_),
    .A3(_05632_),
    .S0(_05682_),
    .S1(_05579_),
    .X(_05825_));
 sky130_fd_sc_hd__nand2_1 _18463_ (.A(_05667_),
    .B(_05683_),
    .Y(_05826_));
 sky130_fd_sc_hd__mux2_1 _18464_ (.A0(_05648_),
    .A1(_05642_),
    .S(_05682_),
    .X(_05827_));
 sky130_fd_sc_hd__o22a_1 _18465_ (.A1(_05741_),
    .A2(_05826_),
    .B1(_05827_),
    .B2(_05667_),
    .X(_05828_));
 sky130_fd_sc_hd__mux2_1 _18466_ (.A0(_05825_),
    .A1(_05828_),
    .S(_05380_),
    .X(_05829_));
 sky130_fd_sc_hd__mux2_1 _18467_ (.A0(_05824_),
    .A1(_05829_),
    .S(_05370_),
    .X(_05830_));
 sky130_fd_sc_hd__mux4_1 _18468_ (.A0(_05327_),
    .A1(_05446_),
    .A2(_05412_),
    .A3(_05441_),
    .S0(_05683_),
    .S1(_05688_),
    .X(_05831_));
 sky130_fd_sc_hd__mux4_1 _18469_ (.A0(_05313_),
    .A1(_05320_),
    .A2(_05506_),
    .A3(_05334_),
    .S0(_05579_),
    .S1(_05663_),
    .X(_05832_));
 sky130_fd_sc_hd__mux2_1 _18470_ (.A0(_05831_),
    .A1(_05832_),
    .S(_05674_),
    .X(_05833_));
 sky130_fd_sc_hd__a2bb2o_1 _18471_ (.A1_N(_05363_),
    .A2_N(_05830_),
    .B1(_05833_),
    .B2(_05781_),
    .X(_05834_));
 sky130_fd_sc_hd__a32o_1 _18472_ (.A1(_05669_),
    .A2(_05665_),
    .A3(_05821_),
    .B1(_05834_),
    .B2(_05749_),
    .X(_05835_));
 sky130_fd_sc_hd__or2_1 _18473_ (.A(_05818_),
    .B(_05835_),
    .X(_05836_));
 sky130_fd_sc_hd__buf_1 _18474_ (.A(_05836_),
    .X(\rvcpu.ALUResultE[1] ));
 sky130_fd_sc_hd__inv_2 _18475_ (.A(_05750_),
    .Y(_05837_));
 sky130_fd_sc_hd__mux4_1 _18476_ (.A0(_05469_),
    .A1(_05475_),
    .A2(_05484_),
    .A3(_05490_),
    .S0(_05769_),
    .S1(_05689_),
    .X(_05838_));
 sky130_fd_sc_hd__mux2_1 _18477_ (.A0(_05456_),
    .A1(_05463_),
    .S(_05684_),
    .X(_05839_));
 sky130_fd_sc_hd__mux2_1 _18478_ (.A0(_05839_),
    .A1(_05760_),
    .S(_05668_),
    .X(_05840_));
 sky130_fd_sc_hd__mux2_1 _18479_ (.A0(_05838_),
    .A1(_05840_),
    .S(_05676_),
    .X(_05841_));
 sky130_fd_sc_hd__nand2_1 _18480_ (.A(_05768_),
    .B(_05761_),
    .Y(_05842_));
 sky130_fd_sc_hd__o21a_1 _18481_ (.A1(_05768_),
    .A2(_05756_),
    .B1(_05842_),
    .X(_05843_));
 sky130_fd_sc_hd__or3_1 _18482_ (.A(_05704_),
    .B(_05669_),
    .C(_05758_),
    .X(_05844_));
 sky130_fd_sc_hd__o21ai_2 _18483_ (.A1(_05676_),
    .A2(_05843_),
    .B1(_05844_),
    .Y(_05845_));
 sky130_fd_sc_hd__mux2_1 _18484_ (.A0(_05841_),
    .A1(_05845_),
    .S(_05692_),
    .X(_05846_));
 sky130_fd_sc_hd__mux2_1 _18485_ (.A0(_05441_),
    .A1(_05421_),
    .S(_05769_),
    .X(_05847_));
 sky130_fd_sc_hd__or2_1 _18486_ (.A(_05349_),
    .B(_05663_),
    .X(_05848_));
 sky130_fd_sc_hd__o211a_1 _18487_ (.A1(_05342_),
    .A2(_05769_),
    .B1(_05848_),
    .C1(_05689_),
    .X(_05849_));
 sky130_fd_sc_hd__a21oi_1 _18488_ (.A1(_05669_),
    .A2(_05847_),
    .B1(_05849_),
    .Y(_05850_));
 sky130_fd_sc_hd__nand2_1 _18489_ (.A(_05587_),
    .B(_05664_),
    .Y(_05851_));
 sky130_fd_sc_hd__o21ai_1 _18490_ (.A1(_05679_),
    .A2(_05664_),
    .B1(_05851_),
    .Y(_05852_));
 sky130_fd_sc_hd__mux2_1 _18491_ (.A0(_05852_),
    .A1(_05770_),
    .S(_05768_),
    .X(_05853_));
 sky130_fd_sc_hd__mux2_1 _18492_ (.A0(_05850_),
    .A1(_05853_),
    .S(_05799_),
    .X(_05854_));
 sky130_fd_sc_hd__mux4_1 _18493_ (.A0(_05320_),
    .A1(_05327_),
    .A2(_05446_),
    .A3(_05412_),
    .S0(_05769_),
    .S1(_05689_),
    .X(_05855_));
 sky130_fd_sc_hd__mux4_1 _18494_ (.A0(_05313_),
    .A1(_05334_),
    .A2(_05500_),
    .A3(_05506_),
    .S0(_05684_),
    .S1(_05668_),
    .X(_05856_));
 sky130_fd_sc_hd__mux2_1 _18495_ (.A0(_05855_),
    .A1(_05856_),
    .S(_05676_),
    .X(_05857_));
 sky130_fd_sc_hd__inv_2 _18496_ (.A(_05782_),
    .Y(_05858_));
 sky130_fd_sc_hd__a2bb2o_1 _18497_ (.A1_N(_05776_),
    .A2_N(_05854_),
    .B1(_05857_),
    .B2(_05858_),
    .X(_05859_));
 sky130_fd_sc_hd__nand2_1 _18498_ (.A(_05383_),
    .B(_05397_),
    .Y(_05860_));
 sky130_fd_sc_hd__o21a_1 _18499_ (.A1(_05383_),
    .A2(_05397_),
    .B1(_05238_),
    .X(_05861_));
 sky130_fd_sc_hd__and3_1 _18500_ (.A(_05398_),
    .B(_05688_),
    .C(_05684_),
    .X(_05862_));
 sky130_fd_sc_hd__a21oi_1 _18501_ (.A1(_05688_),
    .A2(_05684_),
    .B1(_05398_),
    .Y(_05863_));
 sky130_fd_sc_hd__or2_2 _18502_ (.A(_05862_),
    .B(_05863_),
    .X(_05864_));
 sky130_fd_sc_hd__and3_1 _18503_ (.A(_05275_),
    .B(_05709_),
    .C(_05864_),
    .X(_05865_));
 sky130_fd_sc_hd__buf_2 _18504_ (.A(_05590_),
    .X(_05866_));
 sky130_fd_sc_hd__and4_1 _18505_ (.A(_05866_),
    .B(_05692_),
    .C(_05719_),
    .D(_05733_),
    .X(_05867_));
 sky130_fd_sc_hd__a21oi_1 _18506_ (.A1(_05704_),
    .A2(_05382_),
    .B1(_05784_),
    .Y(_05868_));
 sky130_fd_sc_hd__a221o_1 _18507_ (.A1(_05383_),
    .A2(_05726_),
    .B1(_05808_),
    .B2(_05399_),
    .C1(_05868_),
    .X(_05869_));
 sky130_fd_sc_hd__mux2_1 _18508_ (.A0(_05382_),
    .A1(_05388_),
    .S(_05662_),
    .X(_05870_));
 sky130_fd_sc_hd__o22a_1 _18509_ (.A1(_05394_),
    .A2(_05826_),
    .B1(_05870_),
    .B2(_05668_),
    .X(_05871_));
 sky130_fd_sc_hd__nor2_1 _18510_ (.A(_05675_),
    .B(_05871_),
    .Y(_05872_));
 sky130_fd_sc_hd__and3_1 _18511_ (.A(_05789_),
    .B(_05775_),
    .C(_05872_),
    .X(_05873_));
 sky130_fd_sc_hd__a211o_1 _18512_ (.A1(_05865_),
    .A2(_05867_),
    .B1(_05869_),
    .C1(_05873_),
    .X(_05874_));
 sky130_fd_sc_hd__and3_1 _18513_ (.A(_05383_),
    .B(_05577_),
    .C(_05581_),
    .X(_05875_));
 sky130_fd_sc_hd__nor3_1 _18514_ (.A(_05582_),
    .B(_05654_),
    .C(_05875_),
    .Y(_05876_));
 sky130_fd_sc_hd__a211o_1 _18515_ (.A1(_05860_),
    .A2(_05861_),
    .B1(_05874_),
    .C1(_05876_),
    .X(_05877_));
 sky130_fd_sc_hd__a211o_2 _18516_ (.A1(_05837_),
    .A2(_05846_),
    .B1(_05859_),
    .C1(_05877_),
    .X(\rvcpu.ALUResultE[2] ));
 sky130_fd_sc_hd__and2_1 _18517_ (.A(_05704_),
    .B(_05690_),
    .X(_05878_));
 sky130_fd_sc_hd__and3_1 _18518_ (.A(_05370_),
    .B(_05719_),
    .C(_05820_),
    .X(_05879_));
 sky130_fd_sc_hd__a22o_1 _18519_ (.A1(_05378_),
    .A2(_05726_),
    .B1(_05729_),
    .B2(_05377_),
    .X(_05880_));
 sky130_fd_sc_hd__nor2_1 _18520_ (.A(_05374_),
    .B(_05732_),
    .Y(_05881_));
 sky130_fd_sc_hd__a211o_1 _18521_ (.A1(_05879_),
    .A2(_05864_),
    .B1(_05880_),
    .C1(_05881_),
    .X(_05882_));
 sky130_fd_sc_hd__a31o_1 _18522_ (.A1(_05375_),
    .A2(_05702_),
    .A3(_05878_),
    .B1(_05882_),
    .X(_05883_));
 sky130_fd_sc_hd__or3_1 _18523_ (.A(_05584_),
    .B(_05582_),
    .C(_05583_),
    .X(_05884_));
 sky130_fd_sc_hd__and3_1 _18524_ (.A(_05585_),
    .B(_05809_),
    .C(_05884_),
    .X(_05885_));
 sky130_fd_sc_hd__buf_4 _18525_ (.A(_05812_),
    .X(_05886_));
 sky130_fd_sc_hd__a21oi_1 _18526_ (.A1(_05378_),
    .A2(_05400_),
    .B1(_05886_),
    .Y(_05887_));
 sky130_fd_sc_hd__o21a_1 _18527_ (.A1(_05378_),
    .A2(_05400_),
    .B1(_05887_),
    .X(_05888_));
 sky130_fd_sc_hd__nor2_1 _18528_ (.A(_05866_),
    .B(_05805_),
    .Y(_05889_));
 sky130_fd_sc_hd__mux4_1 _18529_ (.A0(_05334_),
    .A1(_05320_),
    .A2(_05327_),
    .A3(_05446_),
    .S0(_05682_),
    .S1(_05579_),
    .X(_05890_));
 sky130_fd_sc_hd__inv_2 _18530_ (.A(_05890_),
    .Y(_05891_));
 sky130_fd_sc_hd__mux4_1 _18531_ (.A0(_05603_),
    .A1(_05565_),
    .A2(_05566_),
    .A3(_05570_),
    .S0(_05668_),
    .S1(_05663_),
    .X(_05892_));
 sky130_fd_sc_hd__mux2_1 _18532_ (.A0(_05891_),
    .A1(_05892_),
    .S(_05674_),
    .X(_05893_));
 sky130_fd_sc_hd__nand2_1 _18533_ (.A(_05692_),
    .B(_05893_),
    .Y(_05894_));
 sky130_fd_sc_hd__mux2_1 _18534_ (.A0(_05349_),
    .A1(_05358_),
    .S(_05684_),
    .X(_05895_));
 sky130_fd_sc_hd__mux2_1 _18535_ (.A0(_05803_),
    .A1(_05895_),
    .S(_05668_),
    .X(_05896_));
 sky130_fd_sc_hd__mux4_1 _18536_ (.A0(_05606_),
    .A1(net102),
    .A2(_05604_),
    .A3(_05596_),
    .S0(_05684_),
    .S1(_05689_),
    .X(_05897_));
 sky130_fd_sc_hd__nor2_1 _18537_ (.A(_05704_),
    .B(_05897_),
    .Y(_05898_));
 sky130_fd_sc_hd__a211o_1 _18538_ (.A1(_05704_),
    .A2(_05896_),
    .B1(_05898_),
    .C1(_05692_),
    .X(_05899_));
 sky130_fd_sc_hd__mux4_1 _18539_ (.A0(_05625_),
    .A1(_05632_),
    .A2(_05633_),
    .A3(_05637_),
    .S0(_05667_),
    .S1(_05663_),
    .X(_05900_));
 sky130_fd_sc_hd__mux4_1 _18540_ (.A0(_05626_),
    .A1(_05621_),
    .A2(_05622_),
    .A3(_05574_),
    .S0(_05682_),
    .S1(_05579_),
    .X(_05901_));
 sky130_fd_sc_hd__or2_1 _18541_ (.A(_05674_),
    .B(_05901_),
    .X(_05902_));
 sky130_fd_sc_hd__o21ai_1 _18542_ (.A1(_05704_),
    .A2(_05900_),
    .B1(_05902_),
    .Y(_05903_));
 sky130_fd_sc_hd__mux4_2 _18543_ (.A0(_05648_),
    .A1(_05642_),
    .A2(_05643_),
    .A3(_05636_),
    .S0(_05683_),
    .S1(_05688_),
    .X(_05904_));
 sky130_fd_sc_hd__nor2_1 _18544_ (.A(_05704_),
    .B(_05711_),
    .Y(_05905_));
 sky130_fd_sc_hd__a21oi_2 _18545_ (.A1(_05704_),
    .A2(_05904_),
    .B1(_05905_),
    .Y(_05906_));
 sky130_fd_sc_hd__mux2_1 _18546_ (.A0(_05903_),
    .A1(_05906_),
    .S(_05370_),
    .X(_05907_));
 sky130_fd_sc_hd__a32o_1 _18547_ (.A1(_05889_),
    .A2(_05894_),
    .A3(_05899_),
    .B1(_05837_),
    .B2(_05907_),
    .X(_05908_));
 sky130_fd_sc_hd__or4_1 _18548_ (.A(_05883_),
    .B(_05885_),
    .C(_05888_),
    .D(_05908_),
    .X(_05909_));
 sky130_fd_sc_hd__clkbuf_2 _18549_ (.A(_05909_),
    .X(\rvcpu.ALUResultE[3] ));
 sky130_fd_sc_hd__a21o_1 _18550_ (.A1(_05585_),
    .A2(_05586_),
    .B1(_05368_),
    .X(_05910_));
 sky130_fd_sc_hd__a31oi_1 _18551_ (.A1(_05368_),
    .A2(_05585_),
    .A3(_05586_),
    .B1(_05654_),
    .Y(_05911_));
 sky130_fd_sc_hd__nor2_1 _18552_ (.A(_05368_),
    .B(_05401_),
    .Y(_05912_));
 sky130_fd_sc_hd__a21o_1 _18553_ (.A1(_05368_),
    .A2(_05401_),
    .B1(_05886_),
    .X(_05913_));
 sky130_fd_sc_hd__mux2_1 _18554_ (.A0(_05365_),
    .A1(_05376_),
    .S(_05662_),
    .X(_05914_));
 sky130_fd_sc_hd__mux2_1 _18555_ (.A0(_05870_),
    .A1(_05914_),
    .S(_05688_),
    .X(_05915_));
 sky130_fd_sc_hd__or4_1 _18556_ (.A(_05398_),
    .B(_05668_),
    .C(_05663_),
    .D(_05394_),
    .X(_05916_));
 sky130_fd_sc_hd__o21a_1 _18557_ (.A1(_05675_),
    .A2(_05915_),
    .B1(_05916_),
    .X(_05917_));
 sky130_fd_sc_hd__a22o_1 _18558_ (.A1(_05367_),
    .A2(_05729_),
    .B1(_05808_),
    .B2(_05366_),
    .X(_05918_));
 sky130_fd_sc_hd__a211oi_1 _18559_ (.A1(_05368_),
    .A2(_05726_),
    .B1(_05821_),
    .C1(_05918_),
    .Y(_05919_));
 sky130_fd_sc_hd__nor2_1 _18560_ (.A(_05674_),
    .B(_05766_),
    .Y(_05920_));
 sky130_fd_sc_hd__a211o_1 _18561_ (.A1(_05675_),
    .A2(_05778_),
    .B1(_05920_),
    .C1(_05776_),
    .X(_05921_));
 sky130_fd_sc_hd__mux2_1 _18562_ (.A0(_05779_),
    .A1(_05751_),
    .S(_05674_),
    .X(_05922_));
 sky130_fd_sc_hd__or2_1 _18563_ (.A(_05782_),
    .B(_05922_),
    .X(_05923_));
 sky130_fd_sc_hd__o2111a_1 _18564_ (.A1(_05790_),
    .A2(_05917_),
    .B1(_05919_),
    .C1(_05921_),
    .D1(_05923_),
    .X(_05924_));
 sky130_fd_sc_hd__or2_2 _18565_ (.A(_05675_),
    .B(_05759_),
    .X(_05925_));
 sky130_fd_sc_hd__mux2_1 _18566_ (.A0(_05752_),
    .A1(_05762_),
    .S(_05674_),
    .X(_05926_));
 sky130_fd_sc_hd__nor2_1 _18567_ (.A(_05692_),
    .B(_05926_),
    .Y(_05927_));
 sky130_fd_sc_hd__a211o_1 _18568_ (.A1(_05692_),
    .A2(_05925_),
    .B1(_05927_),
    .C1(_05750_),
    .X(_05928_));
 sky130_fd_sc_hd__o211a_1 _18569_ (.A1(_05912_),
    .A2(_05913_),
    .B1(_05924_),
    .C1(_05928_),
    .X(_05929_));
 sky130_fd_sc_hd__a21bo_1 _18570_ (.A1(_05910_),
    .A2(_05911_),
    .B1_N(_05929_),
    .X(_05930_));
 sky130_fd_sc_hd__clkbuf_2 _18571_ (.A(_05930_),
    .X(\rvcpu.ALUResultE[4] ));
 sky130_fd_sc_hd__a21o_1 _18572_ (.A1(_05368_),
    .A2(_05401_),
    .B1(_05366_),
    .X(_05931_));
 sky130_fd_sc_hd__xnor2_1 _18573_ (.A(_05931_),
    .B(_05588_),
    .Y(_05932_));
 sky130_fd_sc_hd__a21oi_1 _18574_ (.A1(_05910_),
    .A2(_05591_),
    .B1(_05588_),
    .Y(_05933_));
 sky130_fd_sc_hd__a31o_1 _18575_ (.A1(_05588_),
    .A2(_05910_),
    .A3(_05591_),
    .B1(_05654_),
    .X(_05934_));
 sky130_fd_sc_hd__or2_1 _18576_ (.A(_05676_),
    .B(_05828_),
    .X(_05935_));
 sky130_fd_sc_hd__mux2_1 _18577_ (.A0(_05823_),
    .A1(_05825_),
    .S(_05675_),
    .X(_05936_));
 sky130_fd_sc_hd__mux2_1 _18578_ (.A0(_05935_),
    .A1(_05936_),
    .S(_05696_),
    .X(_05937_));
 sky130_fd_sc_hd__o211a_1 _18579_ (.A1(_05358_),
    .A2(_05664_),
    .B1(_05802_),
    .C1(_05689_),
    .X(_05938_));
 sky130_fd_sc_hd__a21o_1 _18580_ (.A1(_05669_),
    .A2(_05687_),
    .B1(_05938_),
    .X(_05939_));
 sky130_fd_sc_hd__nor2_1 _18581_ (.A(_05799_),
    .B(_05796_),
    .Y(_05940_));
 sky130_fd_sc_hd__a21oi_2 _18582_ (.A1(_05705_),
    .A2(_05939_),
    .B1(_05940_),
    .Y(_05941_));
 sky130_fd_sc_hd__o22a_1 _18583_ (.A1(_05360_),
    .A2(_05784_),
    .B1(_05732_),
    .B2(_05402_),
    .X(_05942_));
 sky130_fd_sc_hd__and2_1 _18584_ (.A(_05709_),
    .B(_05826_),
    .X(_05943_));
 sky130_fd_sc_hd__or2_2 _18585_ (.A(_05676_),
    .B(_05943_),
    .X(_05944_));
 sky130_fd_sc_hd__a22oi_1 _18586_ (.A1(_05588_),
    .A2(_05726_),
    .B1(_05879_),
    .B2(_05944_),
    .Y(_05945_));
 sky130_fd_sc_hd__o211a_1 _18587_ (.A1(_05790_),
    .A2(_05941_),
    .B1(_05942_),
    .C1(_05945_),
    .X(_05946_));
 sky130_fd_sc_hd__nor2_1 _18588_ (.A(_05705_),
    .B(_05831_),
    .Y(_05947_));
 sky130_fd_sc_hd__nor2_1 _18589_ (.A(_05676_),
    .B(_05800_),
    .Y(_05948_));
 sky130_fd_sc_hd__inv_2 _18590_ (.A(_05832_),
    .Y(_05949_));
 sky130_fd_sc_hd__mux2_1 _18591_ (.A0(_05822_),
    .A1(_05949_),
    .S(_05799_),
    .X(_05950_));
 sky130_fd_sc_hd__o32a_1 _18592_ (.A1(_05776_),
    .A2(_05947_),
    .A3(_05948_),
    .B1(_05782_),
    .B2(_05950_),
    .X(_05951_));
 sky130_fd_sc_hd__o211a_1 _18593_ (.A1(_05750_),
    .A2(_05937_),
    .B1(_05946_),
    .C1(_05951_),
    .X(_05952_));
 sky130_fd_sc_hd__o21a_1 _18594_ (.A1(_05933_),
    .A2(_05934_),
    .B1(_05952_),
    .X(_05953_));
 sky130_fd_sc_hd__o21ai_4 _18595_ (.A1(_05886_),
    .A2(_05932_),
    .B1(_05953_),
    .Y(\rvcpu.ALUResultE[5] ));
 sky130_fd_sc_hd__a21oi_1 _18596_ (.A1(_05361_),
    .A2(_05404_),
    .B1(_05356_),
    .Y(_05954_));
 sky130_fd_sc_hd__a311oi_1 _18597_ (.A1(_05356_),
    .A2(_05361_),
    .A3(_05404_),
    .B1(_05886_),
    .C1(_05954_),
    .Y(_05955_));
 sky130_fd_sc_hd__a21o_1 _18598_ (.A1(_05589_),
    .A2(_05593_),
    .B1(_05356_),
    .X(_05956_));
 sky130_fd_sc_hd__or2_1 _18599_ (.A(_05354_),
    .B(_05355_),
    .X(_05957_));
 sky130_fd_sc_hd__or3_1 _18600_ (.A(_05957_),
    .B(_05592_),
    .C(_05933_),
    .X(_05958_));
 sky130_fd_sc_hd__and3_1 _18601_ (.A(_05956_),
    .B(_05809_),
    .C(_05958_),
    .X(_05959_));
 sky130_fd_sc_hd__or3_2 _18602_ (.A(_05676_),
    .B(_05669_),
    .C(_05758_),
    .X(_05960_));
 sky130_fd_sc_hd__nand2_1 _18603_ (.A(_05799_),
    .B(_05840_),
    .Y(_05961_));
 sky130_fd_sc_hd__o21a_1 _18604_ (.A1(_05799_),
    .A2(_05843_),
    .B1(_05961_),
    .X(_05962_));
 sky130_fd_sc_hd__mux2_1 _18605_ (.A0(_05960_),
    .A1(_05962_),
    .S(_05696_),
    .X(_05963_));
 sky130_fd_sc_hd__nor2_1 _18606_ (.A(_05750_),
    .B(_05963_),
    .Y(_05964_));
 sky130_fd_sc_hd__o21ai_1 _18607_ (.A1(_05349_),
    .A2(_05664_),
    .B1(_05851_),
    .Y(_05965_));
 sky130_fd_sc_hd__mux2_1 _18608_ (.A0(_05914_),
    .A1(_05965_),
    .S(_05768_),
    .X(_05966_));
 sky130_fd_sc_hd__mux2_2 _18609_ (.A0(_05871_),
    .A1(_05966_),
    .S(_05799_),
    .X(_05967_));
 sky130_fd_sc_hd__nor2_1 _18610_ (.A(_05799_),
    .B(_05855_),
    .Y(_05968_));
 sky130_fd_sc_hd__a211o_1 _18611_ (.A1(_05705_),
    .A2(_05850_),
    .B1(_05968_),
    .C1(_05776_),
    .X(_05969_));
 sky130_fd_sc_hd__or2_1 _18612_ (.A(_05675_),
    .B(_05856_),
    .X(_05970_));
 sky130_fd_sc_hd__o21ai_2 _18613_ (.A1(_05799_),
    .A2(_05838_),
    .B1(_05970_),
    .Y(_05971_));
 sky130_fd_sc_hd__or2_1 _18614_ (.A(_05675_),
    .B(_05709_),
    .X(_05972_));
 sky130_fd_sc_hd__o2bb2a_1 _18615_ (.A1_N(_05879_),
    .A2_N(_05972_),
    .B1(_05957_),
    .B2(_05786_),
    .X(_05973_));
 sky130_fd_sc_hd__buf_2 _18616_ (.A(_05808_),
    .X(_05974_));
 sky130_fd_sc_hd__o2bb2a_1 _18617_ (.A1_N(_05354_),
    .A2_N(_05974_),
    .B1(_05784_),
    .B2(_05355_),
    .X(_05975_));
 sky130_fd_sc_hd__o211a_1 _18618_ (.A1(_05782_),
    .A2(_05971_),
    .B1(_05973_),
    .C1(_05975_),
    .X(_05976_));
 sky130_fd_sc_hd__o211a_1 _18619_ (.A1(_05790_),
    .A2(_05967_),
    .B1(_05969_),
    .C1(_05976_),
    .X(_05977_));
 sky130_fd_sc_hd__or4b_1 _18620_ (.A(_05955_),
    .B(_05959_),
    .C(_05964_),
    .D_N(_05977_),
    .X(_05978_));
 sky130_fd_sc_hd__clkbuf_2 _18621_ (.A(_05978_),
    .X(\rvcpu.ALUResultE[6] ));
 sky130_fd_sc_hd__a21oi_1 _18622_ (.A1(_05346_),
    .A2(_05405_),
    .B1(_05886_),
    .Y(_05979_));
 sky130_fd_sc_hd__o21a_1 _18623_ (.A1(_05346_),
    .A2(_05405_),
    .B1(_05979_),
    .X(_05980_));
 sky130_fd_sc_hd__nor2_1 _18624_ (.A(_05345_),
    .B(_05784_),
    .Y(_05981_));
 sky130_fd_sc_hd__a221o_1 _18625_ (.A1(_05346_),
    .A2(_05726_),
    .B1(_05974_),
    .B2(_05344_),
    .C1(_05981_),
    .X(_05982_));
 sky130_fd_sc_hd__a311o_1 _18626_ (.A1(_05696_),
    .A2(_05702_),
    .A3(_05691_),
    .B1(_05879_),
    .C1(_05982_),
    .X(_05983_));
 sky130_fd_sc_hd__nor2_1 _18627_ (.A(_05705_),
    .B(_05890_),
    .Y(_05984_));
 sky130_fd_sc_hd__a211o_1 _18628_ (.A1(_05706_),
    .A2(_05897_),
    .B1(_05984_),
    .C1(_05720_),
    .X(_05985_));
 sky130_fd_sc_hd__mux2_1 _18629_ (.A0(_05900_),
    .A1(_05904_),
    .S(_05675_),
    .X(_05986_));
 sky130_fd_sc_hd__or3_1 _18630_ (.A(_05741_),
    .B(_05375_),
    .C(_05719_),
    .X(_05987_));
 sky130_fd_sc_hd__o21a_1 _18631_ (.A1(_05692_),
    .A2(_05986_),
    .B1(_05987_),
    .X(_05988_));
 sky130_fd_sc_hd__mux2_1 _18632_ (.A0(_05901_),
    .A1(_05892_),
    .S(_05799_),
    .X(_05989_));
 sky130_fd_sc_hd__nand2_2 _18633_ (.A(_05363_),
    .B(_05692_),
    .Y(_05990_));
 sky130_fd_sc_hd__o22a_1 _18634_ (.A1(_05363_),
    .A2(_05988_),
    .B1(_05989_),
    .B2(_05990_),
    .X(_05991_));
 sky130_fd_sc_hd__a21oi_1 _18635_ (.A1(_05985_),
    .A2(_05991_),
    .B1(_05805_),
    .Y(_05992_));
 sky130_fd_sc_hd__a21oi_1 _18636_ (.A1(_05594_),
    .A2(_05956_),
    .B1(_05346_),
    .Y(_05993_));
 sky130_fd_sc_hd__and3_1 _18637_ (.A(_05346_),
    .B(_05594_),
    .C(_05956_),
    .X(_05994_));
 sky130_fd_sc_hd__or3_1 _18638_ (.A(_05993_),
    .B(_05654_),
    .C(_05994_),
    .X(_05995_));
 sky130_fd_sc_hd__or4b_1 _18639_ (.A(_05980_),
    .B(_05983_),
    .C(_05992_),
    .D_N(_05995_),
    .X(_05996_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _18640_ (.A(_05996_),
    .X(\rvcpu.ALUResultE[7] ));
 sky130_fd_sc_hd__or2_1 _18641_ (.A(_05425_),
    .B(_05426_),
    .X(_05997_));
 sky130_fd_sc_hd__nand2_1 _18642_ (.A(_05997_),
    .B(_05599_),
    .Y(_05998_));
 sky130_fd_sc_hd__o21a_1 _18643_ (.A1(_05997_),
    .A2(_05599_),
    .B1(_05809_),
    .X(_05999_));
 sky130_fd_sc_hd__xnor2_1 _18644_ (.A(_05997_),
    .B(_05406_),
    .Y(_06000_));
 sky130_fd_sc_hd__or2_1 _18645_ (.A(_05692_),
    .B(_05764_),
    .X(_06001_));
 sky130_fd_sc_hd__o211a_1 _18646_ (.A1(_05866_),
    .A2(_05754_),
    .B1(_06001_),
    .C1(_05720_),
    .X(_06002_));
 sky130_fd_sc_hd__a211oi_1 _18647_ (.A1(_05775_),
    .A2(_05780_),
    .B1(_06002_),
    .C1(_05805_),
    .Y(_06003_));
 sky130_fd_sc_hd__buf_2 _18648_ (.A(_05789_),
    .X(_06004_));
 sky130_fd_sc_hd__mux2_1 _18649_ (.A0(_05604_),
    .A1(_05596_),
    .S(_05664_),
    .X(_06005_));
 sky130_fd_sc_hd__mux2_1 _18650_ (.A0(_05965_),
    .A1(_06005_),
    .S(_05768_),
    .X(_06006_));
 sky130_fd_sc_hd__mux2_1 _18651_ (.A0(_05915_),
    .A1(_06006_),
    .S(_05705_),
    .X(_06007_));
 sky130_fd_sc_hd__nand2_1 _18652_ (.A(_05696_),
    .B(_06007_),
    .Y(_06008_));
 sky130_fd_sc_hd__a21o_1 _18653_ (.A1(_05771_),
    .A2(_05862_),
    .B1(_05696_),
    .X(_06009_));
 sky130_fd_sc_hd__and3_1 _18654_ (.A(_06004_),
    .B(_06008_),
    .C(_06009_),
    .X(_06010_));
 sky130_fd_sc_hd__o21a_1 _18655_ (.A1(_05421_),
    .A2(_05424_),
    .B1(_05729_),
    .X(_06011_));
 sky130_fd_sc_hd__a221o_1 _18656_ (.A1(_05427_),
    .A2(_05726_),
    .B1(_05974_),
    .B2(_05425_),
    .C1(_06011_),
    .X(_06012_));
 sky130_fd_sc_hd__a221o_1 _18657_ (.A1(_05693_),
    .A2(_05820_),
    .B1(_06010_),
    .B2(_05658_),
    .C1(_06012_),
    .X(_06013_));
 sky130_fd_sc_hd__a211o_1 _18658_ (.A1(_05238_),
    .A2(_06000_),
    .B1(_06003_),
    .C1(_06013_),
    .X(_06014_));
 sky130_fd_sc_hd__a21o_1 _18659_ (.A1(_05998_),
    .A2(_05999_),
    .B1(_06014_),
    .X(\rvcpu.ALUResultE[8] ));
 sky130_fd_sc_hd__a21oi_1 _18660_ (.A1(_05427_),
    .A2(_05406_),
    .B1(_05425_),
    .Y(_06015_));
 sky130_fd_sc_hd__xnor2_1 _18661_ (.A(_06015_),
    .B(_05431_),
    .Y(_06016_));
 sky130_fd_sc_hd__nor2_1 _18662_ (.A(_05604_),
    .B(_05424_),
    .Y(_06017_));
 sky130_fd_sc_hd__or2_1 _18663_ (.A(_05442_),
    .B(_05444_),
    .X(_06018_));
 sky130_fd_sc_hd__a211o_1 _18664_ (.A1(_05997_),
    .A2(_05599_),
    .B1(_06017_),
    .C1(_06018_),
    .X(_06019_));
 sky130_fd_sc_hd__a22oi_1 _18665_ (.A1(_05599_),
    .A2(_05601_),
    .B1(_06017_),
    .B2(_06018_),
    .Y(_06020_));
 sky130_fd_sc_hd__and3_1 _18666_ (.A(_05809_),
    .B(_06019_),
    .C(_06020_),
    .X(_06021_));
 sky130_fd_sc_hd__nand2_1 _18667_ (.A(_05866_),
    .B(_05696_),
    .Y(_06022_));
 sky130_fd_sc_hd__nand2_1 _18668_ (.A(_05775_),
    .B(_05833_),
    .Y(_06023_));
 sky130_fd_sc_hd__o221a_1 _18669_ (.A1(_05990_),
    .A2(_05824_),
    .B1(_05829_),
    .B2(_06022_),
    .C1(_06023_),
    .X(_06024_));
 sky130_fd_sc_hd__mux4_2 _18670_ (.A0(_05441_),
    .A1(_05421_),
    .A2(_05342_),
    .A3(_05349_),
    .S0(_05664_),
    .S1(_05669_),
    .X(_06025_));
 sky130_fd_sc_hd__mux2_1 _18671_ (.A0(_05939_),
    .A1(_06025_),
    .S(_05705_),
    .X(_06026_));
 sky130_fd_sc_hd__mux2_1 _18672_ (.A0(_05798_),
    .A1(_06026_),
    .S(_05696_),
    .X(_06027_));
 sky130_fd_sc_hd__a2bb2o_1 _18673_ (.A1_N(_05805_),
    .A2_N(_06024_),
    .B1(_06027_),
    .B2(_05702_),
    .X(_06028_));
 sky130_fd_sc_hd__nand2_1 _18674_ (.A(_05696_),
    .B(_05862_),
    .Y(_06029_));
 sky130_fd_sc_hd__nand2_1 _18675_ (.A(_05693_),
    .B(_05719_),
    .Y(_06030_));
 sky130_fd_sc_hd__nand2_1 _18676_ (.A(_06029_),
    .B(_06030_),
    .Y(_06031_));
 sky130_fd_sc_hd__o21a_1 _18677_ (.A1(_06031_),
    .A2(_05865_),
    .B1(_05820_),
    .X(_06032_));
 sky130_fd_sc_hd__nand2_1 _18678_ (.A(_05444_),
    .B(_05974_),
    .Y(_06033_));
 sky130_fd_sc_hd__o221a_1 _18679_ (.A1(_06018_),
    .A2(_05786_),
    .B1(_05784_),
    .B2(_05442_),
    .C1(_06033_),
    .X(_06034_));
 sky130_fd_sc_hd__or3b_1 _18680_ (.A(_06028_),
    .B(_06032_),
    .C_N(_06034_),
    .X(_06035_));
 sky130_fd_sc_hd__a211o_2 _18681_ (.A1(_05239_),
    .A2(_06016_),
    .B1(_06021_),
    .C1(_06035_),
    .X(\rvcpu.ALUResultE[9] ));
 sky130_fd_sc_hd__a31o_1 _18682_ (.A1(_05427_),
    .A2(_05406_),
    .A3(_05431_),
    .B1(_05445_),
    .X(_06036_));
 sky130_fd_sc_hd__nand2_1 _18683_ (.A(_05419_),
    .B(_06036_),
    .Y(_06037_));
 sky130_fd_sc_hd__o21a_1 _18684_ (.A1(_05419_),
    .A2(_06036_),
    .B1(_05239_),
    .X(_06038_));
 sky130_fd_sc_hd__a21boi_1 _18685_ (.A1(_05599_),
    .A2(_05601_),
    .B1_N(_05605_),
    .Y(_06039_));
 sky130_fd_sc_hd__nand2_1 _18686_ (.A(_05419_),
    .B(_06039_),
    .Y(_06040_));
 sky130_fd_sc_hd__or2_1 _18687_ (.A(_05419_),
    .B(_06039_),
    .X(_06041_));
 sky130_fd_sc_hd__and3_1 _18688_ (.A(_05809_),
    .B(_06040_),
    .C(_06041_),
    .X(_06042_));
 sky130_fd_sc_hd__a22o_1 _18689_ (.A1(_05781_),
    .A2(_05841_),
    .B1(_05857_),
    .B2(_05775_),
    .X(_06043_));
 sky130_fd_sc_hd__a31o_1 _18690_ (.A1(_05866_),
    .A2(_05697_),
    .A3(_05845_),
    .B1(_06043_),
    .X(_06044_));
 sky130_fd_sc_hd__mux4_1 _18691_ (.A0(_05606_),
    .A1(_05429_),
    .A2(_05604_),
    .A3(_05596_),
    .S0(_05664_),
    .S1(_05669_),
    .X(_06045_));
 sky130_fd_sc_hd__mux2_1 _18692_ (.A0(_05966_),
    .A1(_06045_),
    .S(_05705_),
    .X(_06046_));
 sky130_fd_sc_hd__inv_2 _18693_ (.A(_06046_),
    .Y(_06047_));
 sky130_fd_sc_hd__mux2_1 _18694_ (.A0(_05872_),
    .A1(_06047_),
    .S(_05697_),
    .X(_06048_));
 sky130_fd_sc_hd__nor2_1 _18695_ (.A(_05417_),
    .B(_05784_),
    .Y(_06049_));
 sky130_fd_sc_hd__a221o_1 _18696_ (.A1(_05419_),
    .A2(_05727_),
    .B1(_05974_),
    .B2(_05416_),
    .C1(_06049_),
    .X(_06050_));
 sky130_fd_sc_hd__a221o_1 _18697_ (.A1(_05749_),
    .A2(_06044_),
    .B1(_06048_),
    .B2(_05702_),
    .C1(_06050_),
    .X(_06051_));
 sky130_fd_sc_hd__or2_1 _18698_ (.A(_06032_),
    .B(_06051_),
    .X(_06052_));
 sky130_fd_sc_hd__a211o_2 _18699_ (.A1(_06037_),
    .A2(_06038_),
    .B1(_06042_),
    .C1(_06052_),
    .X(\rvcpu.ALUResultE[10] ));
 sky130_fd_sc_hd__a21oi_1 _18700_ (.A1(_05419_),
    .A2(_06036_),
    .B1(_05416_),
    .Y(_06053_));
 sky130_fd_sc_hd__xnor2_1 _18701_ (.A(_05410_),
    .B(_06053_),
    .Y(_06054_));
 sky130_fd_sc_hd__clkbuf_4 _18702_ (.A(_05809_),
    .X(_06055_));
 sky130_fd_sc_hd__nand3_1 _18703_ (.A(_05410_),
    .B(_05607_),
    .C(_06041_),
    .Y(_06056_));
 sky130_fd_sc_hd__a21o_1 _18704_ (.A1(_05607_),
    .A2(_06041_),
    .B1(_05410_),
    .X(_06057_));
 sky130_fd_sc_hd__mux2_1 _18705_ (.A0(_05673_),
    .A1(_05680_),
    .S(_05677_),
    .X(_06058_));
 sky130_fd_sc_hd__mux2_1 _18706_ (.A0(_05878_),
    .A1(_06058_),
    .S(_05697_),
    .X(_06059_));
 sky130_fd_sc_hd__a31o_1 _18707_ (.A1(_05697_),
    .A2(_05749_),
    .A3(_05906_),
    .B1(_05889_),
    .X(_06060_));
 sky130_fd_sc_hd__nand2_1 _18708_ (.A(_05775_),
    .B(_05893_),
    .Y(_06061_));
 sky130_fd_sc_hd__o211ai_1 _18709_ (.A1(_05990_),
    .A2(_05903_),
    .B1(_06060_),
    .C1(_06061_),
    .Y(_06062_));
 sky130_fd_sc_hd__o21ai_1 _18710_ (.A1(_05693_),
    .A2(_05864_),
    .B1(_05820_),
    .Y(_06063_));
 sky130_fd_sc_hd__o2bb2a_1 _18711_ (.A1_N(_05410_),
    .A2_N(_05726_),
    .B1(_05785_),
    .B2(_05447_),
    .X(_06064_));
 sky130_fd_sc_hd__o211a_1 _18712_ (.A1(_05449_),
    .A2(_05732_),
    .B1(_06063_),
    .C1(_06064_),
    .X(_06065_));
 sky130_fd_sc_hd__nand2_1 _18713_ (.A(_06062_),
    .B(_06065_),
    .Y(_06066_));
 sky130_fd_sc_hd__a21o_1 _18714_ (.A1(_05702_),
    .A2(_06059_),
    .B1(_06066_),
    .X(_06067_));
 sky130_fd_sc_hd__a31o_1 _18715_ (.A1(_06055_),
    .A2(_06056_),
    .A3(_06057_),
    .B1(_06067_),
    .X(_06068_));
 sky130_fd_sc_hd__a21o_1 _18716_ (.A1(_05239_),
    .A2(_06054_),
    .B1(_06068_),
    .X(\rvcpu.ALUResultE[11] ));
 sky130_fd_sc_hd__o31ai_2 _18717_ (.A1(_05410_),
    .A2(_05419_),
    .A3(_06039_),
    .B1(_05608_),
    .Y(_06069_));
 sky130_fd_sc_hd__xnor2_1 _18718_ (.A(_05436_),
    .B(_06069_),
    .Y(_06070_));
 sky130_fd_sc_hd__a2bb2o_1 _18719_ (.A1_N(_05776_),
    .A2_N(_05922_),
    .B1(_05926_),
    .B2(_05858_),
    .X(_06071_));
 sky130_fd_sc_hd__and3b_1 _18720_ (.A_N(_05925_),
    .B(_05697_),
    .C(_05837_),
    .X(_06072_));
 sky130_fd_sc_hd__a22o_1 _18721_ (.A1(_05436_),
    .A2(_05727_),
    .B1(_05730_),
    .B2(_05434_),
    .X(_06073_));
 sky130_fd_sc_hd__a211o_1 _18722_ (.A1(_05331_),
    .A2(_05974_),
    .B1(_06072_),
    .C1(_06073_),
    .X(_06074_));
 sky130_fd_sc_hd__o21ai_1 _18723_ (.A1(_05693_),
    .A2(_05944_),
    .B1(_05820_),
    .Y(_06075_));
 sky130_fd_sc_hd__or3b_1 _18724_ (.A(_06071_),
    .B(_06074_),
    .C_N(_06075_),
    .X(_06076_));
 sky130_fd_sc_hd__nand2_1 _18725_ (.A(_05658_),
    .B(_06004_),
    .Y(_06077_));
 sky130_fd_sc_hd__mux4_1 _18726_ (.A0(_05610_),
    .A1(_05408_),
    .A2(_05606_),
    .A3(_05429_),
    .S0(_05665_),
    .S1(_05670_),
    .X(_06078_));
 sky130_fd_sc_hd__mux2_1 _18727_ (.A0(_06006_),
    .A1(_06078_),
    .S(_05706_),
    .X(_06079_));
 sky130_fd_sc_hd__mux2_1 _18728_ (.A0(_05917_),
    .A1(_06079_),
    .S(_05697_),
    .X(_06080_));
 sky130_fd_sc_hd__inv_2 _18729_ (.A(_05436_),
    .Y(_06081_));
 sky130_fd_sc_hd__a21o_1 _18730_ (.A1(_05406_),
    .A2(_05433_),
    .B1(_05451_),
    .X(_06082_));
 sky130_fd_sc_hd__xnor2_1 _18731_ (.A(_06081_),
    .B(_06082_),
    .Y(_06083_));
 sky130_fd_sc_hd__a2bb2o_1 _18732_ (.A1_N(_06077_),
    .A2_N(_06080_),
    .B1(_06083_),
    .B2(_05239_),
    .X(_06084_));
 sky130_fd_sc_hd__a211o_1 _18733_ (.A1(_06055_),
    .A2(_06070_),
    .B1(_06076_),
    .C1(_06084_),
    .X(\rvcpu.ALUResultE[12] ));
 sky130_fd_sc_hd__or2_1 _18734_ (.A(_05324_),
    .B(_05332_),
    .X(_06085_));
 sky130_fd_sc_hd__a21oi_1 _18735_ (.A1(_05436_),
    .A2(_06082_),
    .B1(_05331_),
    .Y(_06086_));
 sky130_fd_sc_hd__or2_1 _18736_ (.A(_06085_),
    .B(_06086_),
    .X(_06087_));
 sky130_fd_sc_hd__a21oi_1 _18737_ (.A1(_06085_),
    .A2(_06086_),
    .B1(_05886_),
    .Y(_06088_));
 sky130_fd_sc_hd__nor2_1 _18738_ (.A(_05610_),
    .B(_05330_),
    .Y(_06089_));
 sky130_fd_sc_hd__a211o_1 _18739_ (.A1(_06081_),
    .A2(_06069_),
    .B1(_06089_),
    .C1(_06085_),
    .X(_06090_));
 sky130_fd_sc_hd__or3b_1 _18740_ (.A(_05436_),
    .B(_05438_),
    .C_N(_06069_),
    .X(_06091_));
 sky130_fd_sc_hd__a21oi_1 _18741_ (.A1(_06085_),
    .A2(_06089_),
    .B1(_05654_),
    .Y(_06092_));
 sky130_fd_sc_hd__inv_2 _18742_ (.A(_06025_),
    .Y(_06093_));
 sky130_fd_sc_hd__mux4_1 _18743_ (.A0(_05437_),
    .A1(_05610_),
    .A2(_05408_),
    .A3(_05606_),
    .S0(_05665_),
    .S1(_05670_),
    .X(_06094_));
 sky130_fd_sc_hd__mux2_1 _18744_ (.A0(_06093_),
    .A1(_06094_),
    .S(_05706_),
    .X(_06095_));
 sky130_fd_sc_hd__mux2_1 _18745_ (.A0(_05941_),
    .A1(_06095_),
    .S(_05697_),
    .X(_06096_));
 sky130_fd_sc_hd__or3_1 _18746_ (.A(_05693_),
    .B(_05805_),
    .C(_05935_),
    .X(_06097_));
 sky130_fd_sc_hd__nand2_1 _18747_ (.A(_05332_),
    .B(_05974_),
    .Y(_06098_));
 sky130_fd_sc_hd__o221a_1 _18748_ (.A1(_06085_),
    .A2(_05786_),
    .B1(_05784_),
    .B2(_05324_),
    .C1(_06098_),
    .X(_06099_));
 sky130_fd_sc_hd__o211a_1 _18749_ (.A1(_05658_),
    .A2(_06097_),
    .B1(_06099_),
    .C1(_06075_),
    .X(_06100_));
 sky130_fd_sc_hd__o221a_1 _18750_ (.A1(_05782_),
    .A2(_05936_),
    .B1(_05950_),
    .B2(_05776_),
    .C1(_06100_),
    .X(_06101_));
 sky130_fd_sc_hd__o21ai_1 _18751_ (.A1(_06077_),
    .A2(_06096_),
    .B1(_06101_),
    .Y(_06102_));
 sky130_fd_sc_hd__a31o_1 _18752_ (.A1(_06090_),
    .A2(_06091_),
    .A3(_06092_),
    .B1(_06102_),
    .X(_06103_));
 sky130_fd_sc_hd__a21o_1 _18753_ (.A1(_06087_),
    .A2(_06088_),
    .B1(_06103_),
    .X(\rvcpu.ALUResultE[13] ));
 sky130_fd_sc_hd__a21o_1 _18754_ (.A1(_05611_),
    .A2(_06091_),
    .B1(_05311_),
    .X(_06104_));
 sky130_fd_sc_hd__nand3_1 _18755_ (.A(_05311_),
    .B(_05611_),
    .C(_06091_),
    .Y(_06105_));
 sky130_fd_sc_hd__a31o_1 _18756_ (.A1(_05436_),
    .A2(_06082_),
    .A3(_05438_),
    .B1(_05333_),
    .X(_06106_));
 sky130_fd_sc_hd__xnor2_1 _18757_ (.A(_05311_),
    .B(_06106_),
    .Y(_06107_));
 sky130_fd_sc_hd__buf_2 _18758_ (.A(_05974_),
    .X(_06108_));
 sky130_fd_sc_hd__buf_2 _18759_ (.A(_05720_),
    .X(_06109_));
 sky130_fd_sc_hd__o22a_1 _18760_ (.A1(_06109_),
    .A2(_05971_),
    .B1(_05962_),
    .B2(_05990_),
    .X(_06110_));
 sky130_fd_sc_hd__o21ai_1 _18761_ (.A1(_05960_),
    .A2(_06022_),
    .B1(_06110_),
    .Y(_06111_));
 sky130_fd_sc_hd__mux4_1 _18762_ (.A0(_05307_),
    .A1(_05437_),
    .A2(_05610_),
    .A3(_05408_),
    .S0(_05665_),
    .S1(_05670_),
    .X(_06112_));
 sky130_fd_sc_hd__mux2_1 _18763_ (.A0(_06045_),
    .A1(_06112_),
    .S(_05706_),
    .X(_06113_));
 sky130_fd_sc_hd__or2_1 _18764_ (.A(_05693_),
    .B(_06113_),
    .X(_06114_));
 sky130_fd_sc_hd__o21ai_1 _18765_ (.A1(_05698_),
    .A2(_05967_),
    .B1(_06114_),
    .Y(_06115_));
 sky130_fd_sc_hd__or2_1 _18766_ (.A(_05334_),
    .B(_05310_),
    .X(_06116_));
 sky130_fd_sc_hd__a221o_1 _18767_ (.A1(_05311_),
    .A2(_05727_),
    .B1(_05730_),
    .B2(_06116_),
    .C1(_05820_),
    .X(_06117_));
 sky130_fd_sc_hd__a221o_1 _18768_ (.A1(_05749_),
    .A2(_06111_),
    .B1(_06115_),
    .B2(_05702_),
    .C1(_06117_),
    .X(_06118_));
 sky130_fd_sc_hd__a21oi_1 _18769_ (.A1(_05335_),
    .A2(_06108_),
    .B1(_06118_),
    .Y(_06119_));
 sky130_fd_sc_hd__o21ai_1 _18770_ (.A1(_05886_),
    .A2(_06107_),
    .B1(_06119_),
    .Y(_06120_));
 sky130_fd_sc_hd__a31o_1 _18771_ (.A1(_06055_),
    .A2(_06104_),
    .A3(_06105_),
    .B1(_06120_),
    .X(\rvcpu.ALUResultE[14] ));
 sky130_fd_sc_hd__a21oi_1 _18772_ (.A1(_05612_),
    .A2(_06104_),
    .B1(_05318_),
    .Y(_06121_));
 sky130_fd_sc_hd__a311oi_1 _18773_ (.A1(_05318_),
    .A2(_05612_),
    .A3(_06104_),
    .B1(_06121_),
    .C1(_05655_),
    .Y(_06122_));
 sky130_fd_sc_hd__a21oi_1 _18774_ (.A1(_05311_),
    .A2(_06106_),
    .B1(_05335_),
    .Y(_06123_));
 sky130_fd_sc_hd__xnor2_1 _18775_ (.A(_05318_),
    .B(_06123_),
    .Y(_06124_));
 sky130_fd_sc_hd__a2bb2o_1 _18776_ (.A1_N(_05315_),
    .A2_N(_05732_),
    .B1(_05730_),
    .B2(_05316_),
    .X(_06125_));
 sky130_fd_sc_hd__a211o_1 _18777_ (.A1(_05318_),
    .A2(_05728_),
    .B1(_05820_),
    .C1(_06125_),
    .X(_06126_));
 sky130_fd_sc_hd__o22a_1 _18778_ (.A1(_05990_),
    .A2(_05986_),
    .B1(_05989_),
    .B2(_06109_),
    .X(_06127_));
 sky130_fd_sc_hd__o31a_1 _18779_ (.A1(_05741_),
    .A2(_05658_),
    .A3(_06029_),
    .B1(_06127_),
    .X(_06128_));
 sky130_fd_sc_hd__a2bb2o_1 _18780_ (.A1_N(_05805_),
    .A2_N(_06128_),
    .B1(_05695_),
    .B2(_05703_),
    .X(_06129_));
 sky130_fd_sc_hd__a211o_1 _18781_ (.A1(_05239_),
    .A2(_06124_),
    .B1(_06126_),
    .C1(_06129_),
    .X(_06130_));
 sky130_fd_sc_hd__or2_1 _18782_ (.A(_06122_),
    .B(_06130_),
    .X(_06131_));
 sky130_fd_sc_hd__clkbuf_1 _18783_ (.A(_06131_),
    .X(\rvcpu.ALUResultE[15] ));
 sky130_fd_sc_hd__nor2_1 _18784_ (.A(_05454_),
    .B(_05513_),
    .Y(_06132_));
 sky130_fd_sc_hd__a21o_1 _18785_ (.A1(_05454_),
    .A2(_05513_),
    .B1(_05886_),
    .X(_06133_));
 sky130_fd_sc_hd__or2_1 _18786_ (.A(_05513_),
    .B(_05616_),
    .X(_06134_));
 sky130_fd_sc_hd__nand2_1 _18787_ (.A(_05513_),
    .B(_05616_),
    .Y(_06135_));
 sky130_fd_sc_hd__nand2_2 _18788_ (.A(_05658_),
    .B(_05749_),
    .Y(_06136_));
 sky130_fd_sc_hd__nor2_1 _18789_ (.A(_05721_),
    .B(_05734_),
    .Y(_06137_));
 sky130_fd_sc_hd__and3_1 _18790_ (.A(_05275_),
    .B(_05864_),
    .C(_05943_),
    .X(_06138_));
 sky130_fd_sc_hd__a21o_1 _18791_ (.A1(_06031_),
    .A2(_06138_),
    .B1(_05819_),
    .X(_06139_));
 sky130_fd_sc_hd__nand2_1 _18792_ (.A(_06137_),
    .B(_06139_),
    .Y(_06140_));
 sky130_fd_sc_hd__mux4_1 _18793_ (.A0(_05313_),
    .A1(_05320_),
    .A2(_05506_),
    .A3(_05334_),
    .S0(_05670_),
    .S1(_05769_),
    .X(_06141_));
 sky130_fd_sc_hd__nand2_1 _18794_ (.A(_05706_),
    .B(_06141_),
    .Y(_06142_));
 sky130_fd_sc_hd__o21ai_1 _18795_ (.A1(_05706_),
    .A2(_06078_),
    .B1(_06142_),
    .Y(_06143_));
 sky130_fd_sc_hd__o221a_1 _18796_ (.A1(_05658_),
    .A2(_05771_),
    .B1(_05720_),
    .B2(_06143_),
    .C1(_06004_),
    .X(_06144_));
 sky130_fd_sc_hd__a21oi_1 _18797_ (.A1(_05781_),
    .A2(_06007_),
    .B1(_05819_),
    .Y(_06145_));
 sky130_fd_sc_hd__a2bb2o_1 _18798_ (.A1_N(_05511_),
    .A2_N(_05784_),
    .B1(_05974_),
    .B2(_05510_),
    .X(_06146_));
 sky130_fd_sc_hd__a21o_1 _18799_ (.A1(_05513_),
    .A2(_05727_),
    .B1(_06146_),
    .X(_06147_));
 sky130_fd_sc_hd__a21oi_1 _18800_ (.A1(_06144_),
    .A2(_06145_),
    .B1(_06147_),
    .Y(_06148_));
 sky130_fd_sc_hd__o211ai_1 _18801_ (.A1(_06136_),
    .A2(_05765_),
    .B1(_06140_),
    .C1(_06148_),
    .Y(_06149_));
 sky130_fd_sc_hd__a31oi_1 _18802_ (.A1(_06134_),
    .A2(_05809_),
    .A3(_06135_),
    .B1(_06149_),
    .Y(_06150_));
 sky130_fd_sc_hd__o21ai_2 _18803_ (.A1(_06132_),
    .A2(_06133_),
    .B1(_06150_),
    .Y(\rvcpu.ALUResultE[16] ));
 sky130_fd_sc_hd__a21oi_1 _18804_ (.A1(_05454_),
    .A2(_05513_),
    .B1(_05510_),
    .Y(_06151_));
 sky130_fd_sc_hd__xnor2_1 _18805_ (.A(_05504_),
    .B(_06151_),
    .Y(_06152_));
 sky130_fd_sc_hd__a31oi_1 _18806_ (.A1(_05504_),
    .A2(_05567_),
    .A3(_06134_),
    .B1(_05655_),
    .Y(_06153_));
 sky130_fd_sc_hd__o211a_1 _18807_ (.A1(_05504_),
    .A2(_06134_),
    .B1(_06153_),
    .C1(_05568_),
    .X(_06154_));
 sky130_fd_sc_hd__a31o_1 _18808_ (.A1(_05698_),
    .A2(_06004_),
    .A3(_05798_),
    .B1(_05703_),
    .X(_06155_));
 sky130_fd_sc_hd__mux4_1 _18809_ (.A0(_05313_),
    .A1(_05334_),
    .A2(_05500_),
    .A3(_05506_),
    .S0(_05664_),
    .S1(_05768_),
    .X(_06156_));
 sky130_fd_sc_hd__inv_2 _18810_ (.A(_06156_),
    .Y(_06157_));
 sky130_fd_sc_hd__mux2_1 _18811_ (.A0(_06094_),
    .A1(_06157_),
    .S(_05706_),
    .X(_06158_));
 sky130_fd_sc_hd__inv_2 _18812_ (.A(_06158_),
    .Y(_06159_));
 sky130_fd_sc_hd__o22a_1 _18813_ (.A1(_05990_),
    .A2(_06026_),
    .B1(_06159_),
    .B2(_06109_),
    .X(_06160_));
 sky130_fd_sc_hd__a2bb2o_1 _18814_ (.A1_N(_05503_),
    .A2_N(_05785_),
    .B1(_05974_),
    .B2(_05502_),
    .X(_06161_));
 sky130_fd_sc_hd__a21oi_1 _18815_ (.A1(_05504_),
    .A2(_05727_),
    .B1(_06161_),
    .Y(_06162_));
 sky130_fd_sc_hd__o211a_1 _18816_ (.A1(_06136_),
    .A2(_05830_),
    .B1(_06140_),
    .C1(_06162_),
    .X(_06163_));
 sky130_fd_sc_hd__a21bo_1 _18817_ (.A1(_06155_),
    .A2(_06160_),
    .B1_N(_06163_),
    .X(_06164_));
 sky130_fd_sc_hd__a211o_1 _18818_ (.A1(_05239_),
    .A2(_06152_),
    .B1(_06154_),
    .C1(_06164_),
    .X(\rvcpu.ALUResultE[17] ));
 sky130_fd_sc_hd__o211a_1 _18819_ (.A1(_05338_),
    .A2(_05453_),
    .B1(_05504_),
    .C1(_05513_),
    .X(_06165_));
 sky130_fd_sc_hd__or3_1 _18820_ (.A(_05497_),
    .B(_05516_),
    .C(_06165_),
    .X(_06166_));
 sky130_fd_sc_hd__o21ai_1 _18821_ (.A1(_05516_),
    .A2(_06165_),
    .B1(_05497_),
    .Y(_06167_));
 sky130_fd_sc_hd__o31a_1 _18822_ (.A1(_05504_),
    .A2(_05513_),
    .A3(_05616_),
    .B1(_05569_),
    .X(_06168_));
 sky130_fd_sc_hd__nand2_1 _18823_ (.A(_05497_),
    .B(_06168_),
    .Y(_06169_));
 sky130_fd_sc_hd__o21a_1 _18824_ (.A1(_05497_),
    .A2(_06168_),
    .B1(_05809_),
    .X(_06170_));
 sky130_fd_sc_hd__mux4_1 _18825_ (.A0(_05313_),
    .A1(_05500_),
    .A2(_05506_),
    .A3(_05490_),
    .S0(_05768_),
    .S1(_05769_),
    .X(_06171_));
 sky130_fd_sc_hd__inv_2 _18826_ (.A(_06171_),
    .Y(_06172_));
 sky130_fd_sc_hd__mux2_1 _18827_ (.A0(_06112_),
    .A1(_06172_),
    .S(_05706_),
    .X(_06173_));
 sky130_fd_sc_hd__inv_2 _18828_ (.A(_06173_),
    .Y(_06174_));
 sky130_fd_sc_hd__a31o_1 _18829_ (.A1(_05697_),
    .A2(_06004_),
    .A3(_05872_),
    .B1(_05702_),
    .X(_06175_));
 sky130_fd_sc_hd__o221a_1 _18830_ (.A1(_05990_),
    .A2(_06047_),
    .B1(_06174_),
    .B2(_06109_),
    .C1(_06175_),
    .X(_06176_));
 sky130_fd_sc_hd__nor2_1 _18831_ (.A(_05494_),
    .B(_05732_),
    .Y(_06177_));
 sky130_fd_sc_hd__a221o_1 _18832_ (.A1(_05497_),
    .A2(_05727_),
    .B1(_05730_),
    .B2(_05495_),
    .C1(_06177_),
    .X(_06178_));
 sky130_fd_sc_hd__a21oi_1 _18833_ (.A1(_05658_),
    .A2(_06030_),
    .B1(_05734_),
    .Y(_06179_));
 sky130_fd_sc_hd__o21a_1 _18834_ (.A1(_05866_),
    .A2(_05864_),
    .B1(_06179_),
    .X(_06180_));
 sky130_fd_sc_hd__a211o_1 _18835_ (.A1(_05889_),
    .A2(_05846_),
    .B1(_06178_),
    .C1(_06180_),
    .X(_06181_));
 sky130_fd_sc_hd__a211o_1 _18836_ (.A1(_06169_),
    .A2(_06170_),
    .B1(_06176_),
    .C1(_06181_),
    .X(_06182_));
 sky130_fd_sc_hd__a31o_1 _18837_ (.A1(_05239_),
    .A2(_06166_),
    .A3(_06167_),
    .B1(_06182_),
    .X(\rvcpu.ALUResultE[18] ));
 sky130_fd_sc_hd__o21a_1 _18838_ (.A1(_05497_),
    .A2(_06168_),
    .B1(_05571_),
    .X(_06183_));
 sky130_fd_sc_hd__xnor2_1 _18839_ (.A(_05488_),
    .B(_06183_),
    .Y(_06184_));
 sky130_fd_sc_hd__mux2_1 _18840_ (.A0(_05700_),
    .A1(_05672_),
    .S(_05677_),
    .X(_06185_));
 sky130_fd_sc_hd__a31o_1 _18841_ (.A1(_05698_),
    .A2(_06004_),
    .A3(_05878_),
    .B1(_05703_),
    .X(_06186_));
 sky130_fd_sc_hd__o221a_1 _18842_ (.A1(_05990_),
    .A2(_06058_),
    .B1(_06185_),
    .B2(_06109_),
    .C1(_06186_),
    .X(_06187_));
 sky130_fd_sc_hd__o22ai_1 _18843_ (.A1(_05486_),
    .A2(_05785_),
    .B1(_05732_),
    .B2(_05487_),
    .Y(_06188_));
 sky130_fd_sc_hd__a2111o_1 _18844_ (.A1(_05488_),
    .A2(_05728_),
    .B1(_06180_),
    .C1(_06187_),
    .D1(_06188_),
    .X(_06189_));
 sky130_fd_sc_hd__a21oi_1 _18845_ (.A1(_05889_),
    .A2(_05907_),
    .B1(_06189_),
    .Y(_06190_));
 sky130_fd_sc_hd__and3_1 _18846_ (.A(_05563_),
    .B(_05494_),
    .C(_06167_),
    .X(_06191_));
 sky130_fd_sc_hd__a21oi_1 _18847_ (.A1(_05494_),
    .A2(_06167_),
    .B1(_05563_),
    .Y(_06192_));
 sky130_fd_sc_hd__or3_1 _18848_ (.A(_05886_),
    .B(_06191_),
    .C(_06192_),
    .X(_06193_));
 sky130_fd_sc_hd__o211ai_2 _18849_ (.A1(_05655_),
    .A2(_06184_),
    .B1(_06190_),
    .C1(_06193_),
    .Y(\rvcpu.ALUResultE[19] ));
 sky130_fd_sc_hd__a41o_1 _18850_ (.A1(_05454_),
    .A2(_05498_),
    .A3(_05504_),
    .A4(_05513_),
    .B1(_05519_),
    .X(_06194_));
 sky130_fd_sc_hd__xor2_1 _18851_ (.A(_05481_),
    .B(_06194_),
    .X(_06195_));
 sky130_fd_sc_hd__a31o_1 _18852_ (.A1(_05275_),
    .A2(_06031_),
    .A3(_05944_),
    .B1(_05819_),
    .X(_06196_));
 sky130_fd_sc_hd__and2_1 _18853_ (.A(_06137_),
    .B(_06196_),
    .X(_06197_));
 sky130_fd_sc_hd__a2bb2o_1 _18854_ (.A1_N(_05480_),
    .A2_N(_05785_),
    .B1(_06108_),
    .B2(_05479_),
    .X(_06198_));
 sky130_fd_sc_hd__a211o_1 _18855_ (.A1(_05481_),
    .A2(_05728_),
    .B1(_06197_),
    .C1(_06198_),
    .X(_06199_));
 sky130_fd_sc_hd__a211o_1 _18856_ (.A1(_05693_),
    .A2(_05925_),
    .B1(_05927_),
    .C1(_06136_),
    .X(_06200_));
 sky130_fd_sc_hd__mux4_1 _18857_ (.A0(_05475_),
    .A1(_05484_),
    .A2(_05490_),
    .A3(_05500_),
    .S0(_05665_),
    .S1(_05670_),
    .X(_06201_));
 sky130_fd_sc_hd__mux2_1 _18858_ (.A0(_06141_),
    .A1(_06201_),
    .S(_05706_),
    .X(_06202_));
 sky130_fd_sc_hd__nor2_1 _18859_ (.A(_06109_),
    .B(_06202_),
    .Y(_06203_));
 sky130_fd_sc_hd__a211o_1 _18860_ (.A1(_05781_),
    .A2(_06079_),
    .B1(_06203_),
    .C1(_05660_),
    .X(_06204_));
 sky130_fd_sc_hd__o21a_1 _18861_ (.A1(_05693_),
    .A2(_05917_),
    .B1(_05866_),
    .X(_06205_));
 sky130_fd_sc_hd__a21oi_1 _18862_ (.A1(_06200_),
    .A2(_06204_),
    .B1(_06205_),
    .Y(_06206_));
 sky130_fd_sc_hd__and3_1 _18863_ (.A(_05481_),
    .B(_05573_),
    .C(_05618_),
    .X(_06207_));
 sky130_fd_sc_hd__or3_1 _18864_ (.A(_05619_),
    .B(_05655_),
    .C(_06207_),
    .X(_06208_));
 sky130_fd_sc_hd__or3b_1 _18865_ (.A(_06199_),
    .B(_06206_),
    .C_N(_06208_),
    .X(_06209_));
 sky130_fd_sc_hd__a21o_1 _18866_ (.A1(_05240_),
    .A2(_06195_),
    .B1(_06209_),
    .X(\rvcpu.ALUResultE[20] ));
 sky130_fd_sc_hd__a21oi_1 _18867_ (.A1(_05481_),
    .A2(_06194_),
    .B1(_05479_),
    .Y(_06210_));
 sky130_fd_sc_hd__xnor2_1 _18868_ (.A(_05473_),
    .B(_06210_),
    .Y(_06211_));
 sky130_fd_sc_hd__or2b_1 _18869_ (.A(_05473_),
    .B_N(_05619_),
    .X(_06212_));
 sky130_fd_sc_hd__o21ai_1 _18870_ (.A1(_05622_),
    .A2(_05478_),
    .B1(_05473_),
    .Y(_06213_));
 sky130_fd_sc_hd__o21a_1 _18871_ (.A1(_05619_),
    .A2(_06213_),
    .B1(_06055_),
    .X(_06214_));
 sky130_fd_sc_hd__nand2_1 _18872_ (.A(_05694_),
    .B(_06095_),
    .Y(_06215_));
 sky130_fd_sc_hd__nor2_1 _18873_ (.A(_05694_),
    .B(_05941_),
    .Y(_06216_));
 sky130_fd_sc_hd__mux4_1 _18874_ (.A0(_05469_),
    .A1(_05475_),
    .A2(_05484_),
    .A3(_05490_),
    .S0(_05666_),
    .S1(_05670_),
    .X(_06217_));
 sky130_fd_sc_hd__mux2_1 _18875_ (.A0(_06156_),
    .A1(_06217_),
    .S(_05707_),
    .X(_06218_));
 sky130_fd_sc_hd__o221a_1 _18876_ (.A1(_05658_),
    .A2(_06216_),
    .B1(_06218_),
    .B2(_06109_),
    .C1(_06004_),
    .X(_06219_));
 sky130_fd_sc_hd__a22o_1 _18877_ (.A1(_05520_),
    .A2(_05730_),
    .B1(_06108_),
    .B2(_05472_),
    .X(_06220_));
 sky130_fd_sc_hd__a211o_1 _18878_ (.A1(_05473_),
    .A2(_05728_),
    .B1(_06197_),
    .C1(_06220_),
    .X(_06221_));
 sky130_fd_sc_hd__nor2_1 _18879_ (.A(_06136_),
    .B(_05937_),
    .Y(_06222_));
 sky130_fd_sc_hd__a211o_1 _18880_ (.A1(_06215_),
    .A2(_06219_),
    .B1(_06221_),
    .C1(_06222_),
    .X(_06223_));
 sky130_fd_sc_hd__a31o_1 _18881_ (.A1(_05623_),
    .A2(_06212_),
    .A3(_06214_),
    .B1(_06223_),
    .X(_06224_));
 sky130_fd_sc_hd__a21o_1 _18882_ (.A1(_05240_),
    .A2(_06211_),
    .B1(_06224_),
    .X(\rvcpu.ALUResultE[21] ));
 sky130_fd_sc_hd__a31o_1 _18883_ (.A1(_05473_),
    .A2(_05481_),
    .A3(_06194_),
    .B1(_05521_),
    .X(_06225_));
 sky130_fd_sc_hd__xor2_1 _18884_ (.A(_05467_),
    .B(_06225_),
    .X(_06226_));
 sky130_fd_sc_hd__nand3_1 _18885_ (.A(_05467_),
    .B(_05624_),
    .C(_06212_),
    .Y(_06227_));
 sky130_fd_sc_hd__a21o_1 _18886_ (.A1(_05624_),
    .A2(_06212_),
    .B1(_05467_),
    .X(_06228_));
 sky130_fd_sc_hd__and3_1 _18887_ (.A(_06055_),
    .B(_06227_),
    .C(_06228_),
    .X(_06229_));
 sky130_fd_sc_hd__mux4_1 _18888_ (.A0(_05463_),
    .A1(_05469_),
    .A2(_05475_),
    .A3(_05484_),
    .S0(_05666_),
    .S1(_05671_),
    .X(_06230_));
 sky130_fd_sc_hd__mux2_1 _18889_ (.A0(_06171_),
    .A1(_06230_),
    .S(_05707_),
    .X(_06231_));
 sky130_fd_sc_hd__o2bb2a_1 _18890_ (.A1_N(_05694_),
    .A2_N(_06113_),
    .B1(_06231_),
    .B2(_06109_),
    .X(_06232_));
 sky130_fd_sc_hd__o21ai_1 _18891_ (.A1(_05694_),
    .A2(_05967_),
    .B1(_05866_),
    .Y(_06233_));
 sky130_fd_sc_hd__nor2_1 _18892_ (.A(_06136_),
    .B(_05963_),
    .Y(_06234_));
 sky130_fd_sc_hd__a2bb2o_1 _18893_ (.A1_N(_05465_),
    .A2_N(_05785_),
    .B1(_06108_),
    .B2(_05466_),
    .X(_06235_));
 sky130_fd_sc_hd__a2111o_1 _18894_ (.A1(_05467_),
    .A2(_05728_),
    .B1(_06179_),
    .C1(_06234_),
    .D1(_06235_),
    .X(_06236_));
 sky130_fd_sc_hd__a31o_1 _18895_ (.A1(_06004_),
    .A2(_06232_),
    .A3(_06233_),
    .B1(_06236_),
    .X(_06237_));
 sky130_fd_sc_hd__a211o_1 _18896_ (.A1(_05240_),
    .A2(_06226_),
    .B1(_06229_),
    .C1(_06237_),
    .X(\rvcpu.ALUResultE[22] ));
 sky130_fd_sc_hd__a21oi_1 _18897_ (.A1(_05467_),
    .A2(_06225_),
    .B1(_05466_),
    .Y(_06238_));
 sky130_fd_sc_hd__xnor2_1 _18898_ (.A(_05461_),
    .B(_06238_),
    .Y(_06239_));
 sky130_fd_sc_hd__a21oi_1 _18899_ (.A1(_05627_),
    .A2(_06228_),
    .B1(_05461_),
    .Y(_06240_));
 sky130_fd_sc_hd__a31o_1 _18900_ (.A1(_05461_),
    .A2(_05627_),
    .A3(_06228_),
    .B1(_05655_),
    .X(_06241_));
 sky130_fd_sc_hd__nor2_1 _18901_ (.A(_06240_),
    .B(_06241_),
    .Y(_06242_));
 sky130_fd_sc_hd__mux2_1 _18902_ (.A0(_05701_),
    .A1(_05678_),
    .S(_05694_),
    .X(_06243_));
 sky130_fd_sc_hd__a2bb2o_1 _18903_ (.A1_N(_05459_),
    .A2_N(_05732_),
    .B1(_05730_),
    .B2(_05458_),
    .X(_06244_));
 sky130_fd_sc_hd__a211o_1 _18904_ (.A1(_05461_),
    .A2(_05728_),
    .B1(_06179_),
    .C1(_06244_),
    .X(_06245_));
 sky130_fd_sc_hd__a31o_1 _18905_ (.A1(_05698_),
    .A2(_05661_),
    .A3(_05691_),
    .B1(_06245_),
    .X(_06246_));
 sky130_fd_sc_hd__nor2_1 _18906_ (.A(_06136_),
    .B(_05988_),
    .Y(_06247_));
 sky130_fd_sc_hd__a211o_1 _18907_ (.A1(_05703_),
    .A2(_06243_),
    .B1(_06246_),
    .C1(_06247_),
    .X(_06248_));
 sky130_fd_sc_hd__a211o_1 _18908_ (.A1(_05240_),
    .A2(_06239_),
    .B1(_06242_),
    .C1(_06248_),
    .X(\rvcpu.ALUResultE[23] ));
 sky130_fd_sc_hd__or2_1 _18909_ (.A(_05525_),
    .B(_05537_),
    .X(_06249_));
 sky130_fd_sc_hd__nand2_1 _18910_ (.A(_05525_),
    .B(_05537_),
    .Y(_06250_));
 sky130_fd_sc_hd__a21oi_1 _18911_ (.A1(_05619_),
    .A2(_05620_),
    .B1(_05629_),
    .Y(_06251_));
 sky130_fd_sc_hd__or2_1 _18912_ (.A(_05535_),
    .B(_05536_),
    .X(_06252_));
 sky130_fd_sc_hd__a211o_1 _18913_ (.A1(_05619_),
    .A2(_05620_),
    .B1(_05629_),
    .C1(_06252_),
    .X(_06253_));
 sky130_fd_sc_hd__o211a_1 _18914_ (.A1(_05537_),
    .A2(_06251_),
    .B1(_06055_),
    .C1(_06253_),
    .X(_06254_));
 sky130_fd_sc_hd__mux4_1 _18915_ (.A0(_05456_),
    .A1(_05469_),
    .A2(_05533_),
    .A3(_05463_),
    .S0(_05670_),
    .S1(_05769_),
    .X(_06255_));
 sky130_fd_sc_hd__a21o_1 _18916_ (.A1(_05707_),
    .A2(_06255_),
    .B1(_06109_),
    .X(_06256_));
 sky130_fd_sc_hd__a21o_1 _18917_ (.A1(_05677_),
    .A2(_06201_),
    .B1(_06256_),
    .X(_06257_));
 sky130_fd_sc_hd__o221a_1 _18918_ (.A1(_05702_),
    .A2(_06010_),
    .B1(_06143_),
    .B2(_05990_),
    .C1(_06257_),
    .X(_06258_));
 sky130_fd_sc_hd__o31a_1 _18919_ (.A1(_05866_),
    .A2(_06031_),
    .A3(_06138_),
    .B1(_06137_),
    .X(_06259_));
 sky130_fd_sc_hd__a2bb2o_1 _18920_ (.A1_N(_05536_),
    .A2_N(_05785_),
    .B1(_05727_),
    .B2(_05537_),
    .X(_06260_));
 sky130_fd_sc_hd__o2bb2a_1 _18921_ (.A1_N(_05535_),
    .A2_N(_06108_),
    .B1(_06136_),
    .B2(_06001_),
    .X(_06261_));
 sky130_fd_sc_hd__or4b_1 _18922_ (.A(_06258_),
    .B(_06259_),
    .C(_06260_),
    .D_N(_06261_),
    .X(_06262_));
 sky130_fd_sc_hd__a311o_1 _18923_ (.A1(_05239_),
    .A2(_06249_),
    .A3(_06250_),
    .B1(_06254_),
    .C1(_06262_),
    .X(\rvcpu.ALUResultE[24] ));
 sky130_fd_sc_hd__a21o_1 _18924_ (.A1(_05525_),
    .A2(_05537_),
    .B1(_05535_),
    .X(_06263_));
 sky130_fd_sc_hd__nand2_1 _18925_ (.A(_05531_),
    .B(_06263_),
    .Y(_06264_));
 sky130_fd_sc_hd__or2_1 _18926_ (.A(_05531_),
    .B(_06263_),
    .X(_06265_));
 sky130_fd_sc_hd__o21ai_1 _18927_ (.A1(_05633_),
    .A2(_05534_),
    .B1(_05531_),
    .Y(_06266_));
 sky130_fd_sc_hd__a21o_1 _18928_ (.A1(_06252_),
    .A2(_05630_),
    .B1(_06266_),
    .X(_06267_));
 sky130_fd_sc_hd__or3_1 _18929_ (.A(_05531_),
    .B(_05537_),
    .C(_06251_),
    .X(_06268_));
 sky130_fd_sc_hd__a221o_1 _18930_ (.A1(_05551_),
    .A2(_05730_),
    .B1(_06108_),
    .B2(_05529_),
    .C1(_06259_),
    .X(_06269_));
 sky130_fd_sc_hd__mux2_1 _18931_ (.A0(_05456_),
    .A1(_05463_),
    .S(_05665_),
    .X(_06270_));
 sky130_fd_sc_hd__mux2_1 _18932_ (.A0(_05714_),
    .A1(_06270_),
    .S(_05670_),
    .X(_06271_));
 sky130_fd_sc_hd__mux2_1 _18933_ (.A0(_06217_),
    .A1(_06271_),
    .S(_05707_),
    .X(_06272_));
 sky130_fd_sc_hd__mux2_1 _18934_ (.A0(_06159_),
    .A1(_06272_),
    .S(_05697_),
    .X(_06273_));
 sky130_fd_sc_hd__a2bb2o_1 _18935_ (.A1_N(_05776_),
    .A2_N(_05829_),
    .B1(_05531_),
    .B2(_05727_),
    .X(_06274_));
 sky130_fd_sc_hd__a221o_1 _18936_ (.A1(_05661_),
    .A2(_06027_),
    .B1(_06273_),
    .B2(_05703_),
    .C1(_06274_),
    .X(_06275_));
 sky130_fd_sc_hd__or2_1 _18937_ (.A(_06269_),
    .B(_06275_),
    .X(_06276_));
 sky130_fd_sc_hd__a41o_1 _18938_ (.A1(_05634_),
    .A2(_06055_),
    .A3(_06267_),
    .A4(_06268_),
    .B1(_06276_),
    .X(_06277_));
 sky130_fd_sc_hd__a31o_1 _18939_ (.A1(_05240_),
    .A2(_06264_),
    .A3(_06265_),
    .B1(_06277_),
    .X(\rvcpu.ALUResultE[25] ));
 sky130_fd_sc_hd__a31o_1 _18940_ (.A1(_05525_),
    .A2(_05531_),
    .A3(_05537_),
    .B1(_05552_),
    .X(_06278_));
 sky130_fd_sc_hd__xor2_1 _18941_ (.A(_05549_),
    .B(_06278_),
    .X(_06279_));
 sky130_fd_sc_hd__o31a_1 _18942_ (.A1(_05531_),
    .A2(_05537_),
    .A3(_06251_),
    .B1(_05635_),
    .X(_06280_));
 sky130_fd_sc_hd__xor2_1 _18943_ (.A(_05549_),
    .B(_06280_),
    .X(_06281_));
 sky130_fd_sc_hd__mux4_1 _18944_ (.A0(_05456_),
    .A1(_05527_),
    .A2(_05533_),
    .A3(_05545_),
    .S0(_05768_),
    .S1(_05769_),
    .X(_06282_));
 sky130_fd_sc_hd__mux2_1 _18945_ (.A0(_06230_),
    .A1(_06282_),
    .S(_05707_),
    .X(_06283_));
 sky130_fd_sc_hd__mux2_1 _18946_ (.A0(_06174_),
    .A1(_06283_),
    .S(_05698_),
    .X(_06284_));
 sky130_fd_sc_hd__or2_1 _18947_ (.A(_06109_),
    .B(_05863_),
    .X(_06285_));
 sky130_fd_sc_hd__nor2_1 _18948_ (.A(_05548_),
    .B(_05785_),
    .Y(_06286_));
 sky130_fd_sc_hd__a221o_1 _18949_ (.A1(_05549_),
    .A2(_05727_),
    .B1(_06108_),
    .B2(_05547_),
    .C1(_06286_),
    .X(_06287_));
 sky130_fd_sc_hd__a31o_1 _18950_ (.A1(_05275_),
    .A2(_05733_),
    .A3(_06285_),
    .B1(_06287_),
    .X(_06288_));
 sky130_fd_sc_hd__a221o_1 _18951_ (.A1(_05806_),
    .A2(_05845_),
    .B1(_06048_),
    .B2(_05661_),
    .C1(_06288_),
    .X(_06289_));
 sky130_fd_sc_hd__a21o_1 _18952_ (.A1(_05703_),
    .A2(_06284_),
    .B1(_06289_),
    .X(_06290_));
 sky130_fd_sc_hd__a221o_1 _18953_ (.A1(_05240_),
    .A2(_06279_),
    .B1(_06281_),
    .B2(_06055_),
    .C1(_06290_),
    .X(\rvcpu.ALUResultE[26] ));
 sky130_fd_sc_hd__and2_1 _18954_ (.A(_05549_),
    .B(_06278_),
    .X(_06291_));
 sky130_fd_sc_hd__o21ai_1 _18955_ (.A1(_05547_),
    .A2(_06291_),
    .B1(_05543_),
    .Y(_06292_));
 sky130_fd_sc_hd__or3_1 _18956_ (.A(_05543_),
    .B(_05547_),
    .C(_06291_),
    .X(_06293_));
 sky130_fd_sc_hd__and3_1 _18957_ (.A(_05240_),
    .B(_06292_),
    .C(_06293_),
    .X(_06294_));
 sky130_fd_sc_hd__o21ai_1 _18958_ (.A1(_05549_),
    .A2(_06280_),
    .B1(_05638_),
    .Y(_06295_));
 sky130_fd_sc_hd__xnor2_1 _18959_ (.A(_05543_),
    .B(_06295_),
    .Y(_06296_));
 sky130_fd_sc_hd__mux2_1 _18960_ (.A0(_05715_),
    .A1(_05699_),
    .S(_05677_),
    .X(_06297_));
 sky130_fd_sc_hd__or2_1 _18961_ (.A(_05698_),
    .B(_06185_),
    .X(_06298_));
 sky130_fd_sc_hd__o211a_1 _18962_ (.A1(_05694_),
    .A2(_06297_),
    .B1(_06298_),
    .C1(_05703_),
    .X(_06299_));
 sky130_fd_sc_hd__a22o_1 _18963_ (.A1(_05543_),
    .A2(_05728_),
    .B1(_06108_),
    .B2(_05542_),
    .X(_06300_));
 sky130_fd_sc_hd__a311o_1 _18964_ (.A1(_05775_),
    .A2(_05724_),
    .A3(_05906_),
    .B1(_06299_),
    .C1(_06300_),
    .X(_06301_));
 sky130_fd_sc_hd__a22o_1 _18965_ (.A1(_05775_),
    .A2(_05906_),
    .B1(_06285_),
    .B2(_05275_),
    .X(_06302_));
 sky130_fd_sc_hd__a22o_1 _18966_ (.A1(_05661_),
    .A2(_06059_),
    .B1(_06302_),
    .B2(_05733_),
    .X(_06303_));
 sky130_fd_sc_hd__a211o_1 _18967_ (.A1(_05554_),
    .A2(_05730_),
    .B1(_06301_),
    .C1(_06303_),
    .X(_06304_));
 sky130_fd_sc_hd__a21o_1 _18968_ (.A1(_06055_),
    .A2(_06296_),
    .B1(_06304_),
    .X(_06305_));
 sky130_fd_sc_hd__or2_1 _18969_ (.A(_06294_),
    .B(_06305_),
    .X(_06306_));
 sky130_fd_sc_hd__buf_1 _18970_ (.A(_06306_),
    .X(\rvcpu.ALUResultE[27] ));
 sky130_fd_sc_hd__xnor2_1 _18971_ (.A(_05305_),
    .B(_05555_),
    .Y(_06307_));
 sky130_fd_sc_hd__a211oi_1 _18972_ (.A1(_05630_),
    .A2(_05631_),
    .B1(_05640_),
    .C1(_05305_),
    .Y(_06308_));
 sky130_fd_sc_hd__a211o_1 _18973_ (.A1(_05305_),
    .A2(_05641_),
    .B1(_05655_),
    .C1(_06308_),
    .X(_06309_));
 sky130_fd_sc_hd__mux4_1 _18974_ (.A0(_05300_),
    .A1(_05539_),
    .A2(_05545_),
    .A3(_05527_),
    .S0(_05666_),
    .S1(_05671_),
    .X(_06310_));
 sky130_fd_sc_hd__mux2_1 _18975_ (.A0(_06255_),
    .A1(_06310_),
    .S(_05707_),
    .X(_06311_));
 sky130_fd_sc_hd__mux2_1 _18976_ (.A0(_06202_),
    .A1(_06311_),
    .S(_05698_),
    .X(_06312_));
 sky130_fd_sc_hd__nand2_1 _18977_ (.A(_05866_),
    .B(_06004_),
    .Y(_06313_));
 sky130_fd_sc_hd__nor2_1 _18978_ (.A(_06313_),
    .B(_06080_),
    .Y(_06314_));
 sky130_fd_sc_hd__o31a_1 _18979_ (.A1(_05694_),
    .A2(_05819_),
    .A3(_05944_),
    .B1(_06137_),
    .X(_06315_));
 sky130_fd_sc_hd__a2bb2o_1 _18980_ (.A1_N(_05303_),
    .A2_N(_05785_),
    .B1(_06108_),
    .B2(_05302_),
    .X(_06316_));
 sky130_fd_sc_hd__o22a_1 _18981_ (.A1(_05305_),
    .A2(_05786_),
    .B1(_05776_),
    .B2(_05925_),
    .X(_06317_));
 sky130_fd_sc_hd__or4b_1 _18982_ (.A(_06314_),
    .B(_06315_),
    .C(_06316_),
    .D_N(_06317_),
    .X(_06318_));
 sky130_fd_sc_hd__a21oi_1 _18983_ (.A1(_05703_),
    .A2(_06312_),
    .B1(_06318_),
    .Y(_06319_));
 sky130_fd_sc_hd__o211ai_4 _18984_ (.A1(_05886_),
    .A2(_06307_),
    .B1(_06309_),
    .C1(_06319_),
    .Y(\rvcpu.ALUResultE[28] ));
 sky130_fd_sc_hd__nor2_1 _18985_ (.A(_05305_),
    .B(_05555_),
    .Y(_06320_));
 sky130_fd_sc_hd__or3_1 _18986_ (.A(_05302_),
    .B(_06320_),
    .C(_05561_),
    .X(_06321_));
 sky130_fd_sc_hd__o21ai_1 _18987_ (.A1(_05302_),
    .A2(_06320_),
    .B1(_05561_),
    .Y(_06322_));
 sky130_fd_sc_hd__nand2_1 _18988_ (.A(_05561_),
    .B(_05644_),
    .Y(_06323_));
 sky130_fd_sc_hd__a21o_1 _18989_ (.A1(_05305_),
    .A2(_05641_),
    .B1(_06323_),
    .X(_06324_));
 sky130_fd_sc_hd__a31oi_1 _18990_ (.A1(_05305_),
    .A2(_05562_),
    .A3(_05641_),
    .B1(_05655_),
    .Y(_06325_));
 sky130_fd_sc_hd__nor2_1 _18991_ (.A(_05298_),
    .B(_05785_),
    .Y(_06326_));
 sky130_fd_sc_hd__a221o_1 _18992_ (.A1(_05561_),
    .A2(_05728_),
    .B1(_06108_),
    .B2(_05556_),
    .C1(_06326_),
    .X(_06327_));
 sky130_fd_sc_hd__mux2_1 _18993_ (.A0(_05713_),
    .A1(_05708_),
    .S(_05768_),
    .X(_06328_));
 sky130_fd_sc_hd__mux2_1 _18994_ (.A0(_06271_),
    .A1(_06328_),
    .S(_05707_),
    .X(_06329_));
 sky130_fd_sc_hd__mux2_1 _18995_ (.A0(_06218_),
    .A1(_06329_),
    .S(_05698_),
    .X(_06330_));
 sky130_fd_sc_hd__a21bo_1 _18996_ (.A1(_06004_),
    .A2(_06330_),
    .B1_N(_06097_),
    .X(_06331_));
 sky130_fd_sc_hd__a2bb2o_1 _18997_ (.A1_N(_06313_),
    .A2_N(_06096_),
    .B1(_06331_),
    .B2(_05658_),
    .X(_06332_));
 sky130_fd_sc_hd__or3_1 _18998_ (.A(_06315_),
    .B(_06327_),
    .C(_06332_),
    .X(_06333_));
 sky130_fd_sc_hd__a31o_1 _18999_ (.A1(_05645_),
    .A2(_06324_),
    .A3(_06325_),
    .B1(_06333_),
    .X(_06334_));
 sky130_fd_sc_hd__a31o_1 _19000_ (.A1(_05240_),
    .A2(_06321_),
    .A3(_06322_),
    .B1(_06334_),
    .X(\rvcpu.ALUResultE[29] ));
 sky130_fd_sc_hd__and2_1 _19001_ (.A(_05288_),
    .B(_05289_),
    .X(_06335_));
 sky130_fd_sc_hd__nor2_1 _19002_ (.A(_05298_),
    .B(_05558_),
    .Y(_06336_));
 sky130_fd_sc_hd__and2_1 _19003_ (.A(_06335_),
    .B(_06336_),
    .X(_06337_));
 sky130_fd_sc_hd__o21ai_1 _19004_ (.A1(_06335_),
    .A2(_06336_),
    .B1(_05240_),
    .Y(_06338_));
 sky130_fd_sc_hd__nand2_1 _19005_ (.A(_05290_),
    .B(_05647_),
    .Y(_06339_));
 sky130_fd_sc_hd__o21a_1 _19006_ (.A1(_05290_),
    .A2(_05647_),
    .B1(_06055_),
    .X(_06340_));
 sky130_fd_sc_hd__nor2_1 _19007_ (.A(_05776_),
    .B(_05960_),
    .Y(_06341_));
 sky130_fd_sc_hd__a2bb2o_1 _19008_ (.A1_N(_05288_),
    .A2_N(_05732_),
    .B1(_05730_),
    .B2(_05289_),
    .X(_06342_));
 sky130_fd_sc_hd__a211o_1 _19009_ (.A1(_06335_),
    .A2(_05728_),
    .B1(_06137_),
    .C1(_06342_),
    .X(_06343_));
 sky130_fd_sc_hd__a211o_1 _19010_ (.A1(_05661_),
    .A2(_06115_),
    .B1(_06341_),
    .C1(_06343_),
    .X(_06344_));
 sky130_fd_sc_hd__nor2_1 _19011_ (.A(_05671_),
    .B(_05757_),
    .Y(_06345_));
 sky130_fd_sc_hd__mux2_1 _19012_ (.A0(_05300_),
    .A1(_05539_),
    .S(_05666_),
    .X(_06346_));
 sky130_fd_sc_hd__a221o_1 _19013_ (.A1(_05755_),
    .A2(_06345_),
    .B1(_06346_),
    .B2(_05671_),
    .C1(_05677_),
    .X(_06347_));
 sky130_fd_sc_hd__o21a_1 _19014_ (.A1(_05707_),
    .A2(_06282_),
    .B1(_06347_),
    .X(_06348_));
 sky130_fd_sc_hd__or2_1 _19015_ (.A(_05698_),
    .B(_06231_),
    .X(_06349_));
 sky130_fd_sc_hd__o211a_1 _19016_ (.A1(_05694_),
    .A2(_06348_),
    .B1(_06349_),
    .C1(_05703_),
    .X(_06350_));
 sky130_fd_sc_hd__a211o_1 _19017_ (.A1(_06339_),
    .A2(_06340_),
    .B1(_06344_),
    .C1(_06350_),
    .X(_06351_));
 sky130_fd_sc_hd__o21bai_2 _19018_ (.A1(_06337_),
    .A2(_06338_),
    .B1_N(_06351_),
    .Y(\rvcpu.ALUResultE[30] ));
 sky130_fd_sc_hd__nand2_1 _19019_ (.A(\rvcpu.dp.plde.ImmExtE[0] ),
    .B(\rvcpu.dp.plde.PCE[0] ),
    .Y(_06352_));
 sky130_fd_sc_hd__or2_1 _19020_ (.A(\rvcpu.dp.plde.ImmExtE[0] ),
    .B(\rvcpu.dp.plde.PCE[0] ),
    .X(_06353_));
 sky130_fd_sc_hd__and2_1 _19021_ (.A(_06352_),
    .B(_06353_),
    .X(_06354_));
 sky130_fd_sc_hd__clkbuf_4 _19022_ (.A(\rvcpu.dp.plde.luiE ),
    .X(_06355_));
 sky130_fd_sc_hd__mux2_1 _19023_ (.A0(_06354_),
    .A1(\rvcpu.dp.plde.ImmExtE[0] ),
    .S(_06355_),
    .X(_06356_));
 sky130_fd_sc_hd__clkbuf_1 _19024_ (.A(_06356_),
    .X(\rvcpu.dp.lAuiPCE[0] ));
 sky130_fd_sc_hd__xor2_2 _19025_ (.A(\rvcpu.dp.plde.ImmExtE[1] ),
    .B(\rvcpu.dp.plde.PCE[1] ),
    .X(_06357_));
 sky130_fd_sc_hd__xnor2_1 _19026_ (.A(_06352_),
    .B(_06357_),
    .Y(_06358_));
 sky130_fd_sc_hd__mux2_1 _19027_ (.A0(_06358_),
    .A1(\rvcpu.dp.plde.ImmExtE[1] ),
    .S(_06355_),
    .X(_06359_));
 sky130_fd_sc_hd__clkbuf_1 _19028_ (.A(_06359_),
    .X(\rvcpu.dp.lAuiPCE[1] ));
 sky130_fd_sc_hd__nand2_1 _19029_ (.A(\rvcpu.dp.plde.ImmExtE[2] ),
    .B(\rvcpu.dp.plde.PCE[2] ),
    .Y(_06360_));
 sky130_fd_sc_hd__or2_1 _19030_ (.A(\rvcpu.dp.plde.ImmExtE[2] ),
    .B(\rvcpu.dp.plde.PCE[2] ),
    .X(_06361_));
 sky130_fd_sc_hd__nand2_1 _19031_ (.A(_06360_),
    .B(_06361_),
    .Y(_06362_));
 sky130_fd_sc_hd__and2_1 _19032_ (.A(\rvcpu.dp.plde.ImmExtE[1] ),
    .B(\rvcpu.dp.plde.PCE[1] ),
    .X(_06363_));
 sky130_fd_sc_hd__a31oi_4 _19033_ (.A1(\rvcpu.dp.plde.ImmExtE[0] ),
    .A2(\rvcpu.dp.plde.PCE[0] ),
    .A3(_06357_),
    .B1(_06363_),
    .Y(_06364_));
 sky130_fd_sc_hd__xor2_2 _19034_ (.A(_06362_),
    .B(_06364_),
    .X(_06365_));
 sky130_fd_sc_hd__mux2_1 _19035_ (.A0(_06365_),
    .A1(\rvcpu.dp.plde.ImmExtE[2] ),
    .S(_06355_),
    .X(_06366_));
 sky130_fd_sc_hd__clkbuf_1 _19036_ (.A(_06366_),
    .X(\rvcpu.dp.lAuiPCE[2] ));
 sky130_fd_sc_hd__nand2_1 _19037_ (.A(\rvcpu.dp.plde.ImmExtE[3] ),
    .B(\rvcpu.dp.plde.PCE[3] ),
    .Y(_06367_));
 sky130_fd_sc_hd__or2_1 _19038_ (.A(\rvcpu.dp.plde.ImmExtE[3] ),
    .B(\rvcpu.dp.plde.PCE[3] ),
    .X(_06368_));
 sky130_fd_sc_hd__nand2_1 _19039_ (.A(_06367_),
    .B(_06368_),
    .Y(_06369_));
 sky130_fd_sc_hd__o21ai_2 _19040_ (.A1(_06362_),
    .A2(_06364_),
    .B1(_06360_),
    .Y(_06370_));
 sky130_fd_sc_hd__xnor2_2 _19041_ (.A(_06369_),
    .B(_06370_),
    .Y(_06371_));
 sky130_fd_sc_hd__mux2_1 _19042_ (.A0(_06371_),
    .A1(\rvcpu.dp.plde.ImmExtE[3] ),
    .S(_06355_),
    .X(_06372_));
 sky130_fd_sc_hd__clkbuf_1 _19043_ (.A(_06372_),
    .X(\rvcpu.dp.lAuiPCE[3] ));
 sky130_fd_sc_hd__and2_1 _19044_ (.A(\rvcpu.dp.plde.ImmExtE[4] ),
    .B(\rvcpu.dp.plde.PCE[4] ),
    .X(_06373_));
 sky130_fd_sc_hd__nor2_1 _19045_ (.A(\rvcpu.dp.plde.ImmExtE[4] ),
    .B(\rvcpu.dp.plde.PCE[4] ),
    .Y(_06374_));
 sky130_fd_sc_hd__nor2_1 _19046_ (.A(_06373_),
    .B(_06374_),
    .Y(_06375_));
 sky130_fd_sc_hd__a21boi_2 _19047_ (.A1(_06368_),
    .A2(_06370_),
    .B1_N(_06367_),
    .Y(_06376_));
 sky130_fd_sc_hd__xnor2_2 _19048_ (.A(_06375_),
    .B(_06376_),
    .Y(_06377_));
 sky130_fd_sc_hd__mux2_1 _19049_ (.A0(_06377_),
    .A1(\rvcpu.dp.plde.ImmExtE[4] ),
    .S(_06355_),
    .X(_06378_));
 sky130_fd_sc_hd__clkbuf_1 _19050_ (.A(_06378_),
    .X(\rvcpu.dp.lAuiPCE[4] ));
 sky130_fd_sc_hd__nand2_1 _19051_ (.A(\rvcpu.dp.plde.ImmExtE[4] ),
    .B(\rvcpu.dp.plde.PCE[4] ),
    .Y(_06379_));
 sky130_fd_sc_hd__o21a_1 _19052_ (.A1(_06374_),
    .A2(_06376_),
    .B1(_06379_),
    .X(_06380_));
 sky130_fd_sc_hd__nor2_1 _19053_ (.A(\rvcpu.dp.plde.ImmExtE[5] ),
    .B(\rvcpu.dp.plde.PCE[5] ),
    .Y(_06381_));
 sky130_fd_sc_hd__and2_1 _19054_ (.A(\rvcpu.dp.plde.ImmExtE[5] ),
    .B(\rvcpu.dp.plde.PCE[5] ),
    .X(_06382_));
 sky130_fd_sc_hd__nor2_1 _19055_ (.A(_06381_),
    .B(_06382_),
    .Y(_06383_));
 sky130_fd_sc_hd__xnor2_2 _19056_ (.A(_06380_),
    .B(_06383_),
    .Y(_06384_));
 sky130_fd_sc_hd__mux2_1 _19057_ (.A0(_06384_),
    .A1(\rvcpu.dp.plde.ImmExtE[5] ),
    .S(_06355_),
    .X(_06385_));
 sky130_fd_sc_hd__clkbuf_1 _19058_ (.A(_06385_),
    .X(\rvcpu.dp.lAuiPCE[5] ));
 sky130_fd_sc_hd__nand2_1 _19059_ (.A(\rvcpu.dp.plde.ImmExtE[6] ),
    .B(\rvcpu.dp.plde.PCE[6] ),
    .Y(_06386_));
 sky130_fd_sc_hd__or2_1 _19060_ (.A(\rvcpu.dp.plde.ImmExtE[6] ),
    .B(\rvcpu.dp.plde.PCE[6] ),
    .X(_06387_));
 sky130_fd_sc_hd__nand2_1 _19061_ (.A(_06386_),
    .B(_06387_),
    .Y(_06388_));
 sky130_fd_sc_hd__inv_2 _19062_ (.A(_06382_),
    .Y(_06389_));
 sky130_fd_sc_hd__o211a_1 _19063_ (.A1(_06374_),
    .A2(_06376_),
    .B1(_06389_),
    .C1(_06379_),
    .X(_06390_));
 sky130_fd_sc_hd__nor2_1 _19064_ (.A(_06381_),
    .B(_06390_),
    .Y(_06391_));
 sky130_fd_sc_hd__xnor2_2 _19065_ (.A(_06388_),
    .B(_06391_),
    .Y(_06392_));
 sky130_fd_sc_hd__mux2_1 _19066_ (.A0(_06392_),
    .A1(\rvcpu.dp.plde.ImmExtE[6] ),
    .S(_06355_),
    .X(_06393_));
 sky130_fd_sc_hd__clkbuf_1 _19067_ (.A(_06393_),
    .X(\rvcpu.dp.lAuiPCE[6] ));
 sky130_fd_sc_hd__nand2_1 _19068_ (.A(\rvcpu.dp.plde.ImmExtE[7] ),
    .B(\rvcpu.dp.plde.PCE[7] ),
    .Y(_06394_));
 sky130_fd_sc_hd__or2_1 _19069_ (.A(\rvcpu.dp.plde.ImmExtE[7] ),
    .B(\rvcpu.dp.plde.PCE[7] ),
    .X(_06395_));
 sky130_fd_sc_hd__nand2_1 _19070_ (.A(_06394_),
    .B(_06395_),
    .Y(_06396_));
 sky130_fd_sc_hd__o31a_1 _19071_ (.A1(_06381_),
    .A2(_06388_),
    .A3(_06390_),
    .B1(_06386_),
    .X(_06397_));
 sky130_fd_sc_hd__xor2_2 _19072_ (.A(_06396_),
    .B(_06397_),
    .X(_06398_));
 sky130_fd_sc_hd__mux2_1 _19073_ (.A0(_06398_),
    .A1(\rvcpu.dp.plde.ImmExtE[7] ),
    .S(_06355_),
    .X(_06399_));
 sky130_fd_sc_hd__clkbuf_1 _19074_ (.A(_06399_),
    .X(\rvcpu.dp.lAuiPCE[7] ));
 sky130_fd_sc_hd__or2_1 _19075_ (.A(\rvcpu.dp.plde.ImmExtE[8] ),
    .B(\rvcpu.dp.plde.PCE[8] ),
    .X(_06400_));
 sky130_fd_sc_hd__nand2_1 _19076_ (.A(\rvcpu.dp.plde.ImmExtE[8] ),
    .B(\rvcpu.dp.plde.PCE[8] ),
    .Y(_06401_));
 sky130_fd_sc_hd__nand2_1 _19077_ (.A(_06400_),
    .B(_06401_),
    .Y(_06402_));
 sky130_fd_sc_hd__o21ai_2 _19078_ (.A1(_06396_),
    .A2(_06397_),
    .B1(_06394_),
    .Y(_06403_));
 sky130_fd_sc_hd__xnor2_1 _19079_ (.A(_06402_),
    .B(_06403_),
    .Y(_06404_));
 sky130_fd_sc_hd__mux2_1 _19080_ (.A0(_06404_),
    .A1(\rvcpu.dp.plde.ImmExtE[8] ),
    .S(_06355_),
    .X(_06405_));
 sky130_fd_sc_hd__clkbuf_1 _19081_ (.A(_06405_),
    .X(\rvcpu.dp.lAuiPCE[8] ));
 sky130_fd_sc_hd__and2_1 _19082_ (.A(\rvcpu.dp.plde.ImmExtE[9] ),
    .B(\rvcpu.dp.plde.PCE[9] ),
    .X(_06406_));
 sky130_fd_sc_hd__nor2_1 _19083_ (.A(\rvcpu.dp.plde.ImmExtE[9] ),
    .B(\rvcpu.dp.plde.PCE[9] ),
    .Y(_06407_));
 sky130_fd_sc_hd__nor2_1 _19084_ (.A(_06406_),
    .B(_06407_),
    .Y(_06408_));
 sky130_fd_sc_hd__and2_1 _19085_ (.A(\rvcpu.dp.plde.ImmExtE[8] ),
    .B(\rvcpu.dp.plde.PCE[8] ),
    .X(_06409_));
 sky130_fd_sc_hd__a21oi_1 _19086_ (.A1(_06400_),
    .A2(_06403_),
    .B1(_06409_),
    .Y(_06410_));
 sky130_fd_sc_hd__xnor2_2 _19087_ (.A(_06408_),
    .B(_06410_),
    .Y(_06411_));
 sky130_fd_sc_hd__mux2_1 _19088_ (.A0(_06411_),
    .A1(\rvcpu.dp.plde.ImmExtE[9] ),
    .S(_06355_),
    .X(_06412_));
 sky130_fd_sc_hd__clkbuf_1 _19089_ (.A(_06412_),
    .X(\rvcpu.dp.lAuiPCE[9] ));
 sky130_fd_sc_hd__nor2_1 _19090_ (.A(\rvcpu.dp.plde.ImmExtE[10] ),
    .B(\rvcpu.dp.plde.PCE[10] ),
    .Y(_06413_));
 sky130_fd_sc_hd__nand2_1 _19091_ (.A(\rvcpu.dp.plde.ImmExtE[10] ),
    .B(\rvcpu.dp.plde.PCE[10] ),
    .Y(_06414_));
 sky130_fd_sc_hd__and2b_1 _19092_ (.A_N(_06413_),
    .B(_06414_),
    .X(_06415_));
 sky130_fd_sc_hd__a211oi_2 _19093_ (.A1(_06400_),
    .A2(_06403_),
    .B1(_06406_),
    .C1(_06409_),
    .Y(_06416_));
 sky130_fd_sc_hd__or2_1 _19094_ (.A(_06407_),
    .B(_06416_),
    .X(_06417_));
 sky130_fd_sc_hd__xnor2_1 _19095_ (.A(_06415_),
    .B(_06417_),
    .Y(_06418_));
 sky130_fd_sc_hd__clkbuf_4 _19096_ (.A(\rvcpu.dp.plde.luiE ),
    .X(_06419_));
 sky130_fd_sc_hd__mux2_1 _19097_ (.A0(_06418_),
    .A1(\rvcpu.dp.plde.ImmExtE[10] ),
    .S(_06419_),
    .X(_06420_));
 sky130_fd_sc_hd__clkbuf_1 _19098_ (.A(_06420_),
    .X(\rvcpu.dp.lAuiPCE[10] ));
 sky130_fd_sc_hd__or2_1 _19099_ (.A(\rvcpu.dp.plde.ImmExtE[11] ),
    .B(\rvcpu.dp.plde.PCE[11] ),
    .X(_06421_));
 sky130_fd_sc_hd__nand2_1 _19100_ (.A(\rvcpu.dp.plde.ImmExtE[11] ),
    .B(\rvcpu.dp.plde.PCE[11] ),
    .Y(_06422_));
 sky130_fd_sc_hd__nand2_1 _19101_ (.A(_06421_),
    .B(_06422_),
    .Y(_06423_));
 sky130_fd_sc_hd__o21ai_1 _19102_ (.A1(_06413_),
    .A2(_06417_),
    .B1(_06414_),
    .Y(_06424_));
 sky130_fd_sc_hd__xnor2_1 _19103_ (.A(_06423_),
    .B(_06424_),
    .Y(_06425_));
 sky130_fd_sc_hd__mux2_1 _19104_ (.A0(_06425_),
    .A1(\rvcpu.dp.plde.ImmExtE[11] ),
    .S(_06419_),
    .X(_06426_));
 sky130_fd_sc_hd__clkbuf_1 _19105_ (.A(_06426_),
    .X(\rvcpu.dp.lAuiPCE[11] ));
 sky130_fd_sc_hd__and2_1 _19106_ (.A(\rvcpu.dp.plde.ImmExtE[12] ),
    .B(\rvcpu.dp.plde.PCE[12] ),
    .X(_06427_));
 sky130_fd_sc_hd__nor2_1 _19107_ (.A(\rvcpu.dp.plde.ImmExtE[12] ),
    .B(\rvcpu.dp.plde.PCE[12] ),
    .Y(_06428_));
 sky130_fd_sc_hd__nor2_1 _19108_ (.A(_06427_),
    .B(_06428_),
    .Y(_06429_));
 sky130_fd_sc_hd__o311ai_4 _19109_ (.A1(_06407_),
    .A2(_06413_),
    .A3(_06416_),
    .B1(_06422_),
    .C1(_06414_),
    .Y(_06430_));
 sky130_fd_sc_hd__nand2_1 _19110_ (.A(_06421_),
    .B(_06430_),
    .Y(_06431_));
 sky130_fd_sc_hd__xnor2_1 _19111_ (.A(_06429_),
    .B(_06431_),
    .Y(_06432_));
 sky130_fd_sc_hd__mux2_1 _19112_ (.A0(_06432_),
    .A1(\rvcpu.dp.plde.ImmExtE[12] ),
    .S(_06419_),
    .X(_06433_));
 sky130_fd_sc_hd__clkbuf_1 _19113_ (.A(_06433_),
    .X(\rvcpu.dp.lAuiPCE[12] ));
 sky130_fd_sc_hd__nor2_1 _19114_ (.A(\rvcpu.dp.plde.ImmExtE[13] ),
    .B(\rvcpu.dp.plde.PCE[13] ),
    .Y(_06434_));
 sky130_fd_sc_hd__and2_1 _19115_ (.A(\rvcpu.dp.plde.ImmExtE[13] ),
    .B(\rvcpu.dp.plde.PCE[13] ),
    .X(_06435_));
 sky130_fd_sc_hd__or2_1 _19116_ (.A(_06434_),
    .B(_06435_),
    .X(_06436_));
 sky130_fd_sc_hd__a31o_1 _19117_ (.A1(_06421_),
    .A2(_06429_),
    .A3(_06430_),
    .B1(_06427_),
    .X(_06437_));
 sky130_fd_sc_hd__xnor2_1 _19118_ (.A(_06436_),
    .B(_06437_),
    .Y(_06438_));
 sky130_fd_sc_hd__mux2_1 _19119_ (.A0(_06438_),
    .A1(\rvcpu.dp.plde.ImmExtE[13] ),
    .S(_06419_),
    .X(_06439_));
 sky130_fd_sc_hd__clkbuf_1 _19120_ (.A(_06439_),
    .X(\rvcpu.dp.lAuiPCE[13] ));
 sky130_fd_sc_hd__inv_2 _19121_ (.A(_06434_),
    .Y(_06440_));
 sky130_fd_sc_hd__nand2_1 _19122_ (.A(\rvcpu.dp.plde.ImmExtE[14] ),
    .B(\rvcpu.dp.plde.PCE[14] ),
    .Y(_06441_));
 sky130_fd_sc_hd__or2_1 _19123_ (.A(\rvcpu.dp.plde.ImmExtE[14] ),
    .B(\rvcpu.dp.plde.PCE[14] ),
    .X(_06442_));
 sky130_fd_sc_hd__and2_1 _19124_ (.A(_06441_),
    .B(_06442_),
    .X(_06443_));
 sky130_fd_sc_hd__a311o_1 _19125_ (.A1(_06421_),
    .A2(_06429_),
    .A3(_06430_),
    .B1(_06435_),
    .C1(_06427_),
    .X(_06444_));
 sky130_fd_sc_hd__nand3_1 _19126_ (.A(_06440_),
    .B(_06443_),
    .C(_06444_),
    .Y(_06445_));
 sky130_fd_sc_hd__a21o_1 _19127_ (.A1(_06440_),
    .A2(_06444_),
    .B1(_06443_),
    .X(_06446_));
 sky130_fd_sc_hd__and2_1 _19128_ (.A(_06445_),
    .B(_06446_),
    .X(_06447_));
 sky130_fd_sc_hd__mux2_1 _19129_ (.A0(_06447_),
    .A1(\rvcpu.dp.plde.ImmExtE[14] ),
    .S(_06419_),
    .X(_06448_));
 sky130_fd_sc_hd__clkbuf_1 _19130_ (.A(_06448_),
    .X(\rvcpu.dp.lAuiPCE[14] ));
 sky130_fd_sc_hd__nor2_1 _19131_ (.A(\rvcpu.dp.plde.ImmExtE[15] ),
    .B(\rvcpu.dp.plde.PCE[15] ),
    .Y(_06449_));
 sky130_fd_sc_hd__nand2_1 _19132_ (.A(\rvcpu.dp.plde.ImmExtE[15] ),
    .B(\rvcpu.dp.plde.PCE[15] ),
    .Y(_06450_));
 sky130_fd_sc_hd__or2b_1 _19133_ (.A(_06449_),
    .B_N(_06450_),
    .X(_06451_));
 sky130_fd_sc_hd__nand2_1 _19134_ (.A(_06441_),
    .B(_06445_),
    .Y(_06452_));
 sky130_fd_sc_hd__xnor2_1 _19135_ (.A(_06451_),
    .B(_06452_),
    .Y(_06453_));
 sky130_fd_sc_hd__mux2_1 _19136_ (.A0(_06453_),
    .A1(\rvcpu.dp.plde.ImmExtE[15] ),
    .S(_06419_),
    .X(_06454_));
 sky130_fd_sc_hd__clkbuf_1 _19137_ (.A(_06454_),
    .X(\rvcpu.dp.lAuiPCE[15] ));
 sky130_fd_sc_hd__or2_1 _19138_ (.A(\rvcpu.dp.plde.ImmExtE[16] ),
    .B(\rvcpu.dp.plde.PCE[16] ),
    .X(_06455_));
 sky130_fd_sc_hd__nand2_1 _19139_ (.A(\rvcpu.dp.plde.ImmExtE[16] ),
    .B(\rvcpu.dp.plde.PCE[16] ),
    .Y(_06456_));
 sky130_fd_sc_hd__and2_1 _19140_ (.A(_06455_),
    .B(_06456_),
    .X(_06457_));
 sky130_fd_sc_hd__nand2_1 _19141_ (.A(_06441_),
    .B(_06450_),
    .Y(_06458_));
 sky130_fd_sc_hd__inv_2 _19142_ (.A(_06458_),
    .Y(_06459_));
 sky130_fd_sc_hd__a21o_1 _19143_ (.A1(_06445_),
    .A2(_06459_),
    .B1(_06449_),
    .X(_06460_));
 sky130_fd_sc_hd__xnor2_1 _19144_ (.A(_06457_),
    .B(_06460_),
    .Y(_06461_));
 sky130_fd_sc_hd__mux2_1 _19145_ (.A0(_06461_),
    .A1(\rvcpu.dp.plde.ImmExtE[16] ),
    .S(_06419_),
    .X(_06462_));
 sky130_fd_sc_hd__clkbuf_1 _19146_ (.A(_06462_),
    .X(\rvcpu.dp.lAuiPCE[16] ));
 sky130_fd_sc_hd__nor2_1 _19147_ (.A(\rvcpu.dp.plde.ImmExtE[17] ),
    .B(\rvcpu.dp.plde.PCE[17] ),
    .Y(_06463_));
 sky130_fd_sc_hd__nand2_1 _19148_ (.A(\rvcpu.dp.plde.ImmExtE[17] ),
    .B(\rvcpu.dp.plde.PCE[17] ),
    .Y(_06464_));
 sky130_fd_sc_hd__or2b_1 _19149_ (.A(_06463_),
    .B_N(_06464_),
    .X(_06465_));
 sky130_fd_sc_hd__inv_2 _19150_ (.A(_06457_),
    .Y(_06466_));
 sky130_fd_sc_hd__o21ai_1 _19151_ (.A1(_06466_),
    .A2(_06460_),
    .B1(_06456_),
    .Y(_06467_));
 sky130_fd_sc_hd__xnor2_1 _19152_ (.A(_06465_),
    .B(_06467_),
    .Y(_06468_));
 sky130_fd_sc_hd__mux2_1 _19153_ (.A0(_06468_),
    .A1(\rvcpu.dp.plde.ImmExtE[17] ),
    .S(_06419_),
    .X(_06469_));
 sky130_fd_sc_hd__clkbuf_1 _19154_ (.A(_06469_),
    .X(\rvcpu.dp.lAuiPCE[17] ));
 sky130_fd_sc_hd__nand3b_1 _19155_ (.A_N(_06463_),
    .B(\rvcpu.dp.plde.PCE[16] ),
    .C(\rvcpu.dp.plde.ImmExtE[16] ),
    .Y(_06470_));
 sky130_fd_sc_hd__nand2_1 _19156_ (.A(_06464_),
    .B(_06470_),
    .Y(_06471_));
 sky130_fd_sc_hd__a2111oi_1 _19157_ (.A1(_06445_),
    .A2(_06459_),
    .B1(_06465_),
    .C1(_06449_),
    .D1(_06466_),
    .Y(_06472_));
 sky130_fd_sc_hd__nand2_1 _19158_ (.A(\rvcpu.dp.plde.ImmExtE[18] ),
    .B(\rvcpu.dp.plde.PCE[18] ),
    .Y(_06473_));
 sky130_fd_sc_hd__or2_1 _19159_ (.A(\rvcpu.dp.plde.ImmExtE[18] ),
    .B(\rvcpu.dp.plde.PCE[18] ),
    .X(_06474_));
 sky130_fd_sc_hd__and2_1 _19160_ (.A(_06473_),
    .B(_06474_),
    .X(_06475_));
 sky130_fd_sc_hd__o21ai_2 _19161_ (.A1(_06471_),
    .A2(net38),
    .B1(_06475_),
    .Y(_06476_));
 sky130_fd_sc_hd__or3_1 _19162_ (.A(_06475_),
    .B(_06471_),
    .C(net38),
    .X(_06477_));
 sky130_fd_sc_hd__and2_1 _19163_ (.A(_06476_),
    .B(_06477_),
    .X(_06478_));
 sky130_fd_sc_hd__mux2_1 _19164_ (.A0(_06478_),
    .A1(\rvcpu.dp.plde.ImmExtE[18] ),
    .S(_06419_),
    .X(_06479_));
 sky130_fd_sc_hd__clkbuf_1 _19165_ (.A(_06479_),
    .X(\rvcpu.dp.lAuiPCE[18] ));
 sky130_fd_sc_hd__nor2_1 _19166_ (.A(\rvcpu.dp.plde.ImmExtE[19] ),
    .B(\rvcpu.dp.plde.PCE[19] ),
    .Y(_06480_));
 sky130_fd_sc_hd__nand2_1 _19167_ (.A(\rvcpu.dp.plde.ImmExtE[19] ),
    .B(\rvcpu.dp.plde.PCE[19] ),
    .Y(_06481_));
 sky130_fd_sc_hd__or2b_1 _19168_ (.A(_06480_),
    .B_N(_06481_),
    .X(_06482_));
 sky130_fd_sc_hd__nand2_1 _19169_ (.A(_06473_),
    .B(_06476_),
    .Y(_06483_));
 sky130_fd_sc_hd__xnor2_1 _19170_ (.A(_06482_),
    .B(_06483_),
    .Y(_06484_));
 sky130_fd_sc_hd__mux2_1 _19171_ (.A0(_06484_),
    .A1(\rvcpu.dp.plde.ImmExtE[19] ),
    .S(_06419_),
    .X(_06485_));
 sky130_fd_sc_hd__clkbuf_1 _19172_ (.A(_06485_),
    .X(\rvcpu.dp.lAuiPCE[19] ));
 sky130_fd_sc_hd__or2_1 _19173_ (.A(\rvcpu.dp.plde.ImmExtE[20] ),
    .B(\rvcpu.dp.plde.PCE[20] ),
    .X(_06486_));
 sky130_fd_sc_hd__nand2_1 _19174_ (.A(\rvcpu.dp.plde.ImmExtE[20] ),
    .B(\rvcpu.dp.plde.PCE[20] ),
    .Y(_06487_));
 sky130_fd_sc_hd__nand2_1 _19175_ (.A(_06486_),
    .B(_06487_),
    .Y(_06488_));
 sky130_fd_sc_hd__a31o_1 _19176_ (.A1(_06473_),
    .A2(_06476_),
    .A3(_06481_),
    .B1(_06480_),
    .X(_06489_));
 sky130_fd_sc_hd__nand2_1 _19177_ (.A(_06488_),
    .B(_06489_),
    .Y(_06490_));
 sky130_fd_sc_hd__a311o_1 _19178_ (.A1(_06473_),
    .A2(_06476_),
    .A3(_06481_),
    .B1(_06488_),
    .C1(_06480_),
    .X(_06491_));
 sky130_fd_sc_hd__and2_1 _19179_ (.A(_06490_),
    .B(_06491_),
    .X(_06492_));
 sky130_fd_sc_hd__clkbuf_4 _19180_ (.A(\rvcpu.dp.plde.luiE ),
    .X(_06493_));
 sky130_fd_sc_hd__mux2_1 _19181_ (.A0(_06492_),
    .A1(\rvcpu.dp.plde.ImmExtE[20] ),
    .S(_06493_),
    .X(_06494_));
 sky130_fd_sc_hd__clkbuf_1 _19182_ (.A(_06494_),
    .X(\rvcpu.dp.lAuiPCE[20] ));
 sky130_fd_sc_hd__nor2_1 _19183_ (.A(\rvcpu.dp.plde.ImmExtE[21] ),
    .B(\rvcpu.dp.plde.PCE[21] ),
    .Y(_06495_));
 sky130_fd_sc_hd__nand2_1 _19184_ (.A(\rvcpu.dp.plde.ImmExtE[21] ),
    .B(\rvcpu.dp.plde.PCE[21] ),
    .Y(_06496_));
 sky130_fd_sc_hd__or2b_1 _19185_ (.A(_06495_),
    .B_N(_06496_),
    .X(_06497_));
 sky130_fd_sc_hd__nand2_1 _19186_ (.A(_06487_),
    .B(_06491_),
    .Y(_06498_));
 sky130_fd_sc_hd__xnor2_1 _19187_ (.A(_06497_),
    .B(_06498_),
    .Y(_06499_));
 sky130_fd_sc_hd__mux2_1 _19188_ (.A0(_06499_),
    .A1(\rvcpu.dp.plde.ImmExtE[21] ),
    .S(_06493_),
    .X(_06500_));
 sky130_fd_sc_hd__clkbuf_1 _19189_ (.A(_06500_),
    .X(\rvcpu.dp.lAuiPCE[21] ));
 sky130_fd_sc_hd__nand2_1 _19190_ (.A(\rvcpu.dp.plde.ImmExtE[22] ),
    .B(\rvcpu.dp.plde.PCE[22] ),
    .Y(_06501_));
 sky130_fd_sc_hd__or2_1 _19191_ (.A(\rvcpu.dp.plde.ImmExtE[22] ),
    .B(\rvcpu.dp.plde.PCE[22] ),
    .X(_06502_));
 sky130_fd_sc_hd__nand2_1 _19192_ (.A(_06501_),
    .B(_06502_),
    .Y(_06503_));
 sky130_fd_sc_hd__a31o_1 _19193_ (.A1(_06487_),
    .A2(_06491_),
    .A3(_06496_),
    .B1(_06495_),
    .X(_06504_));
 sky130_fd_sc_hd__xor2_1 _19194_ (.A(_06503_),
    .B(_06504_),
    .X(_06505_));
 sky130_fd_sc_hd__mux2_1 _19195_ (.A0(_06505_),
    .A1(\rvcpu.dp.plde.ImmExtE[22] ),
    .S(_06493_),
    .X(_06506_));
 sky130_fd_sc_hd__clkbuf_1 _19196_ (.A(_06506_),
    .X(\rvcpu.dp.lAuiPCE[22] ));
 sky130_fd_sc_hd__nor2_1 _19197_ (.A(\rvcpu.dp.plde.ImmExtE[23] ),
    .B(\rvcpu.dp.plde.PCE[23] ),
    .Y(_06507_));
 sky130_fd_sc_hd__nand2_1 _19198_ (.A(\rvcpu.dp.plde.ImmExtE[23] ),
    .B(\rvcpu.dp.plde.PCE[23] ),
    .Y(_06508_));
 sky130_fd_sc_hd__or2b_1 _19199_ (.A(_06507_),
    .B_N(_06508_),
    .X(_06509_));
 sky130_fd_sc_hd__a311o_1 _19200_ (.A1(_06487_),
    .A2(_06491_),
    .A3(_06496_),
    .B1(_06503_),
    .C1(_06495_),
    .X(_06510_));
 sky130_fd_sc_hd__nand2_1 _19201_ (.A(_06501_),
    .B(_06510_),
    .Y(_06511_));
 sky130_fd_sc_hd__xnor2_1 _19202_ (.A(_06509_),
    .B(_06511_),
    .Y(_06512_));
 sky130_fd_sc_hd__mux2_1 _19203_ (.A0(_06512_),
    .A1(\rvcpu.dp.plde.ImmExtE[23] ),
    .S(_06493_),
    .X(_06513_));
 sky130_fd_sc_hd__clkbuf_1 _19204_ (.A(_06513_),
    .X(\rvcpu.dp.lAuiPCE[23] ));
 sky130_fd_sc_hd__nand2_1 _19205_ (.A(\rvcpu.dp.plde.ImmExtE[24] ),
    .B(\rvcpu.dp.plde.PCE[24] ),
    .Y(_06514_));
 sky130_fd_sc_hd__or2_1 _19206_ (.A(\rvcpu.dp.plde.ImmExtE[24] ),
    .B(\rvcpu.dp.plde.PCE[24] ),
    .X(_06515_));
 sky130_fd_sc_hd__and2_1 _19207_ (.A(_06514_),
    .B(_06515_),
    .X(_06516_));
 sky130_fd_sc_hd__a31o_1 _19208_ (.A1(_06501_),
    .A2(_06510_),
    .A3(_06508_),
    .B1(_06507_),
    .X(_06517_));
 sky130_fd_sc_hd__xnor2_1 _19209_ (.A(_06516_),
    .B(_06517_),
    .Y(_06518_));
 sky130_fd_sc_hd__mux2_1 _19210_ (.A0(_06518_),
    .A1(\rvcpu.dp.plde.ImmExtE[24] ),
    .S(_06493_),
    .X(_06519_));
 sky130_fd_sc_hd__clkbuf_1 _19211_ (.A(_06519_),
    .X(\rvcpu.dp.lAuiPCE[24] ));
 sky130_fd_sc_hd__inv_2 _19212_ (.A(_06516_),
    .Y(_06520_));
 sky130_fd_sc_hd__o21ai_1 _19213_ (.A1(_06520_),
    .A2(_06517_),
    .B1(_06514_),
    .Y(_06521_));
 sky130_fd_sc_hd__or2_1 _19214_ (.A(\rvcpu.dp.plde.ImmExtE[25] ),
    .B(\rvcpu.dp.plde.PCE[25] ),
    .X(_06522_));
 sky130_fd_sc_hd__nand2_1 _19215_ (.A(\rvcpu.dp.plde.ImmExtE[25] ),
    .B(\rvcpu.dp.plde.PCE[25] ),
    .Y(_06523_));
 sky130_fd_sc_hd__nand2_1 _19216_ (.A(_06522_),
    .B(_06523_),
    .Y(_06524_));
 sky130_fd_sc_hd__xnor2_1 _19217_ (.A(_06521_),
    .B(_06524_),
    .Y(_06525_));
 sky130_fd_sc_hd__mux2_1 _19218_ (.A0(_06525_),
    .A1(\rvcpu.dp.plde.ImmExtE[25] ),
    .S(_06493_),
    .X(_06526_));
 sky130_fd_sc_hd__clkbuf_1 _19219_ (.A(_06526_),
    .X(\rvcpu.dp.lAuiPCE[25] ));
 sky130_fd_sc_hd__nand2_1 _19220_ (.A(\rvcpu.dp.plde.ImmExtE[26] ),
    .B(\rvcpu.dp.plde.PCE[26] ),
    .Y(_06527_));
 sky130_fd_sc_hd__or2_1 _19221_ (.A(\rvcpu.dp.plde.ImmExtE[26] ),
    .B(\rvcpu.dp.plde.PCE[26] ),
    .X(_06528_));
 sky130_fd_sc_hd__nand2_1 _19222_ (.A(_06527_),
    .B(_06528_),
    .Y(_06529_));
 sky130_fd_sc_hd__a21boi_2 _19223_ (.A1(_06521_),
    .A2(_06522_),
    .B1_N(_06523_),
    .Y(_06530_));
 sky130_fd_sc_hd__xor2_1 _19224_ (.A(_06529_),
    .B(_06530_),
    .X(_06531_));
 sky130_fd_sc_hd__mux2_1 _19225_ (.A0(_06531_),
    .A1(\rvcpu.dp.plde.ImmExtE[26] ),
    .S(_06493_),
    .X(_06532_));
 sky130_fd_sc_hd__clkbuf_1 _19226_ (.A(_06532_),
    .X(\rvcpu.dp.lAuiPCE[26] ));
 sky130_fd_sc_hd__nor2_1 _19227_ (.A(\rvcpu.dp.plde.ImmExtE[26] ),
    .B(\rvcpu.dp.plde.PCE[26] ),
    .Y(_06533_));
 sky130_fd_sc_hd__o21ai_1 _19228_ (.A1(_06533_),
    .A2(_06530_),
    .B1(_06527_),
    .Y(_06534_));
 sky130_fd_sc_hd__or2_1 _19229_ (.A(\rvcpu.dp.plde.ImmExtE[27] ),
    .B(\rvcpu.dp.plde.PCE[27] ),
    .X(_06535_));
 sky130_fd_sc_hd__nand2_1 _19230_ (.A(\rvcpu.dp.plde.ImmExtE[27] ),
    .B(\rvcpu.dp.plde.PCE[27] ),
    .Y(_06536_));
 sky130_fd_sc_hd__nand2_1 _19231_ (.A(_06535_),
    .B(_06536_),
    .Y(_06537_));
 sky130_fd_sc_hd__xnor2_1 _19232_ (.A(_06534_),
    .B(_06537_),
    .Y(_06538_));
 sky130_fd_sc_hd__mux2_1 _19233_ (.A0(_06538_),
    .A1(\rvcpu.dp.plde.ImmExtE[27] ),
    .S(_06493_),
    .X(_06539_));
 sky130_fd_sc_hd__clkbuf_1 _19234_ (.A(_06539_),
    .X(\rvcpu.dp.lAuiPCE[27] ));
 sky130_fd_sc_hd__and2_1 _19235_ (.A(\rvcpu.dp.plde.ImmExtE[28] ),
    .B(\rvcpu.dp.plde.PCE[28] ),
    .X(_06540_));
 sky130_fd_sc_hd__nor2_1 _19236_ (.A(\rvcpu.dp.plde.ImmExtE[28] ),
    .B(\rvcpu.dp.plde.PCE[28] ),
    .Y(_06541_));
 sky130_fd_sc_hd__nor2_1 _19237_ (.A(_06540_),
    .B(_06541_),
    .Y(_06542_));
 sky130_fd_sc_hd__o211ai_1 _19238_ (.A1(_06533_),
    .A2(_06530_),
    .B1(_06536_),
    .C1(_06527_),
    .Y(_06543_));
 sky130_fd_sc_hd__nand2_1 _19239_ (.A(_06535_),
    .B(_06543_),
    .Y(_06544_));
 sky130_fd_sc_hd__xnor2_1 _19240_ (.A(_06542_),
    .B(_06544_),
    .Y(_06545_));
 sky130_fd_sc_hd__mux2_1 _19241_ (.A0(_06545_),
    .A1(\rvcpu.dp.plde.ImmExtE[28] ),
    .S(_06493_),
    .X(_06546_));
 sky130_fd_sc_hd__clkbuf_1 _19242_ (.A(_06546_),
    .X(\rvcpu.dp.lAuiPCE[28] ));
 sky130_fd_sc_hd__a31o_1 _19243_ (.A1(_06535_),
    .A2(_06542_),
    .A3(_06543_),
    .B1(_06540_),
    .X(_06547_));
 sky130_fd_sc_hd__or2_1 _19244_ (.A(\rvcpu.dp.plde.ImmExtE[29] ),
    .B(\rvcpu.dp.plde.PCE[29] ),
    .X(_06548_));
 sky130_fd_sc_hd__nand2_1 _19245_ (.A(\rvcpu.dp.plde.ImmExtE[29] ),
    .B(\rvcpu.dp.plde.PCE[29] ),
    .Y(_06549_));
 sky130_fd_sc_hd__nand2_1 _19246_ (.A(_06548_),
    .B(_06549_),
    .Y(_06550_));
 sky130_fd_sc_hd__xnor2_1 _19247_ (.A(_06547_),
    .B(_06550_),
    .Y(_06551_));
 sky130_fd_sc_hd__mux2_1 _19248_ (.A0(_06551_),
    .A1(\rvcpu.dp.plde.ImmExtE[29] ),
    .S(_06493_),
    .X(_06552_));
 sky130_fd_sc_hd__clkbuf_1 _19249_ (.A(_06552_),
    .X(\rvcpu.dp.lAuiPCE[29] ));
 sky130_fd_sc_hd__and2_1 _19250_ (.A(\rvcpu.dp.plde.ImmExtE[30] ),
    .B(\rvcpu.dp.plde.PCE[30] ),
    .X(_06553_));
 sky130_fd_sc_hd__nor2_1 _19251_ (.A(\rvcpu.dp.plde.ImmExtE[30] ),
    .B(\rvcpu.dp.plde.PCE[30] ),
    .Y(_06554_));
 sky130_fd_sc_hd__nor2_1 _19252_ (.A(_06553_),
    .B(_06554_),
    .Y(_06555_));
 sky130_fd_sc_hd__or2b_1 _19253_ (.A(_06547_),
    .B_N(_06549_),
    .X(_06556_));
 sky130_fd_sc_hd__nand2_1 _19254_ (.A(_06548_),
    .B(_06556_),
    .Y(_06557_));
 sky130_fd_sc_hd__xnor2_1 _19255_ (.A(_06555_),
    .B(_06557_),
    .Y(_06558_));
 sky130_fd_sc_hd__mux2_1 _19256_ (.A0(_06558_),
    .A1(\rvcpu.dp.plde.ImmExtE[30] ),
    .S(\rvcpu.dp.plde.luiE ),
    .X(_06559_));
 sky130_fd_sc_hd__clkbuf_1 _19257_ (.A(_06559_),
    .X(\rvcpu.dp.lAuiPCE[30] ));
 sky130_fd_sc_hd__a31o_1 _19258_ (.A1(_06548_),
    .A2(_06555_),
    .A3(_06556_),
    .B1(_06553_),
    .X(_06560_));
 sky130_fd_sc_hd__xnor2_1 _19259_ (.A(\rvcpu.dp.plde.ImmExtE[31] ),
    .B(\rvcpu.dp.plde.PCE[31] ),
    .Y(_06561_));
 sky130_fd_sc_hd__xnor2_1 _19260_ (.A(_06560_),
    .B(_06561_),
    .Y(_06562_));
 sky130_fd_sc_hd__mux2_1 _19261_ (.A0(_06562_),
    .A1(\rvcpu.dp.plde.ImmExtE[31] ),
    .S(\rvcpu.dp.plde.luiE ),
    .X(_06563_));
 sky130_fd_sc_hd__clkbuf_1 _19262_ (.A(_06563_),
    .X(\rvcpu.dp.lAuiPCE[31] ));
 sky130_fd_sc_hd__and2_1 _19263_ (.A(_05275_),
    .B(_05280_),
    .X(_06564_));
 sky130_fd_sc_hd__o21a_1 _19264_ (.A1(_06564_),
    .A2(_05559_),
    .B1(_05655_),
    .X(_06565_));
 sky130_fd_sc_hd__a2bb2o_1 _19265_ (.A1_N(_05655_),
    .A2_N(_05743_),
    .B1(_06565_),
    .B2(_05281_),
    .X(_00002_));
 sky130_fd_sc_hd__or3b_1 _19266_ (.A(\rvcpu.dp.plfd.InstrD[3] ),
    .B(\rvcpu.dp.plfd.InstrD[2] ),
    .C_N(\rvcpu.dp.plfd.InstrD[0] ),
    .X(_06566_));
 sky130_fd_sc_hd__nor3b_2 _19267_ (.A(_06566_),
    .B(\rvcpu.dp.plfd.InstrD[6] ),
    .C_N(\rvcpu.dp.plfd.InstrD[4] ),
    .Y(_06567_));
 sky130_fd_sc_hd__inv_2 _19268_ (.A(\rvcpu.dp.plfd.InstrD[14] ),
    .Y(_06568_));
 sky130_fd_sc_hd__a311o_1 _19269_ (.A1(\rvcpu.c.ad.funct7b5 ),
    .A2(_06568_),
    .A3(\rvcpu.c.ad.opb5 ),
    .B1(\rvcpu.dp.plfd.InstrD[12] ),
    .C1(\rvcpu.dp.plfd.InstrD[13] ),
    .X(_06569_));
 sky130_fd_sc_hd__inv_2 _19270_ (.A(\rvcpu.c.ad.funct7b5 ),
    .Y(_06570_));
 sky130_fd_sc_hd__o211ai_1 _19271_ (.A1(_06570_),
    .A2(\rvcpu.dp.plfd.InstrD[13] ),
    .B1(\rvcpu.dp.plfd.InstrD[12] ),
    .C1(\rvcpu.dp.plfd.InstrD[14] ),
    .Y(_06571_));
 sky130_fd_sc_hd__nor2_1 _19272_ (.A(\rvcpu.dp.plfd.InstrD[4] ),
    .B(_06566_),
    .Y(_06572_));
 sky130_fd_sc_hd__and3_1 _19273_ (.A(\rvcpu.dp.plfd.InstrD[6] ),
    .B(\rvcpu.c.ad.opb5 ),
    .C(_06572_),
    .X(_06573_));
 sky130_fd_sc_hd__a31o_1 _19274_ (.A1(_06567_),
    .A2(_06569_),
    .A3(_06571_),
    .B1(_06573_),
    .X(_04447_));
 sky130_fd_sc_hd__and2b_1 _19275_ (.A_N(\rvcpu.dp.plfd.InstrD[13] ),
    .B(\rvcpu.dp.plfd.InstrD[12] ),
    .X(_06574_));
 sky130_fd_sc_hd__nand2_1 _19276_ (.A(\rvcpu.dp.plfd.InstrD[14] ),
    .B(\rvcpu.c.ad.opb5 ),
    .Y(_06575_));
 sky130_fd_sc_hd__or3b_1 _19277_ (.A(_06575_),
    .B(\rvcpu.c.ad.funct7b5 ),
    .C_N(_06574_),
    .X(_06576_));
 sky130_fd_sc_hd__o211a_1 _19278_ (.A1(\rvcpu.dp.plfd.InstrD[14] ),
    .A2(_06574_),
    .B1(_06576_),
    .C1(_06567_),
    .X(_04448_));
 sky130_fd_sc_hd__a21oi_1 _19279_ (.A1(_06570_),
    .A2(\rvcpu.dp.plfd.InstrD[12] ),
    .B1(\rvcpu.dp.plfd.InstrD[13] ),
    .Y(_06577_));
 sky130_fd_sc_hd__mux2_1 _19280_ (.A0(\rvcpu.dp.plfd.InstrD[13] ),
    .A1(_06577_),
    .S(\rvcpu.dp.plfd.InstrD[14] ),
    .X(_06578_));
 sky130_fd_sc_hd__and2_1 _19281_ (.A(_06567_),
    .B(_06578_),
    .X(_06579_));
 sky130_fd_sc_hd__clkbuf_1 _19282_ (.A(_06579_),
    .X(_04449_));
 sky130_fd_sc_hd__o211a_1 _19283_ (.A1(_06570_),
    .A2(_06575_),
    .B1(_06574_),
    .C1(_06567_),
    .X(_04450_));
 sky130_fd_sc_hd__nand2b_2 _19284_ (.A_N(\rvcpu.dp.plem.funct3M[1] ),
    .B(\rvcpu.dp.plem.funct3M[0] ),
    .Y(_06580_));
 sky130_fd_sc_hd__or3b_1 _19285_ (.A(\rvcpu.dp.plem.funct3M[0] ),
    .B(\rvcpu.dp.plem.funct3M[2] ),
    .C_N(\rvcpu.dp.plem.funct3M[1] ),
    .X(_06581_));
 sky130_fd_sc_hd__clkbuf_4 _19286_ (.A(_06581_),
    .X(_06582_));
 sky130_fd_sc_hd__nand2_2 _19287_ (.A(_06580_),
    .B(_06582_),
    .Y(_06583_));
 sky130_fd_sc_hd__clkinv_4 _19288_ (.A(net1),
    .Y(_06584_));
 sky130_fd_sc_hd__buf_8 _19289_ (.A(_06584_),
    .X(_06585_));
 sky130_fd_sc_hd__nand2_2 _19290_ (.A(_06585_),
    .B(\rvcpu.dp.plem.ALUResultM[1] ),
    .Y(_06586_));
 sky130_fd_sc_hd__buf_4 _19291_ (.A(_06585_),
    .X(_06587_));
 sky130_fd_sc_hd__nand2_2 _19292_ (.A(_06587_),
    .B(\rvcpu.dp.plem.ALUResultM[0] ),
    .Y(_06588_));
 sky130_fd_sc_hd__and2_1 _19293_ (.A(_06586_),
    .B(_06588_),
    .X(_06589_));
 sky130_fd_sc_hd__or2_1 _19294_ (.A(_06583_),
    .B(_06589_),
    .X(_06590_));
 sky130_fd_sc_hd__buf_8 _19295_ (.A(net1),
    .X(_06591_));
 sky130_fd_sc_hd__nor2_8 _19296_ (.A(_06591_),
    .B(_05347_),
    .Y(_06592_));
 sky130_fd_sc_hd__and2_1 _19297_ (.A(_06585_),
    .B(\rvcpu.dp.plem.ALUResultM[7] ),
    .X(_06593_));
 sky130_fd_sc_hd__buf_8 _19298_ (.A(_06593_),
    .X(_06594_));
 sky130_fd_sc_hd__nor2_4 _19299_ (.A(_06592_),
    .B(_06594_),
    .Y(_06595_));
 sky130_fd_sc_hd__clkbuf_16 _19300_ (.A(_06595_),
    .X(_06596_));
 sky130_fd_sc_hd__and2_1 _19301_ (.A(_06585_),
    .B(\rvcpu.dp.plem.ALUResultM[5] ),
    .X(_06597_));
 sky130_fd_sc_hd__buf_6 _19302_ (.A(_06597_),
    .X(_06598_));
 sky130_fd_sc_hd__buf_6 _19303_ (.A(_06598_),
    .X(_06599_));
 sky130_fd_sc_hd__clkbuf_16 _19304_ (.A(_06599_),
    .X(_06600_));
 sky130_fd_sc_hd__buf_8 _19305_ (.A(_06600_),
    .X(_06601_));
 sky130_fd_sc_hd__clkbuf_8 _19306_ (.A(_06601_),
    .X(_06602_));
 sky130_fd_sc_hd__buf_8 _19307_ (.A(_06602_),
    .X(_06603_));
 sky130_fd_sc_hd__buf_4 _19308_ (.A(_06603_),
    .X(_06604_));
 sky130_fd_sc_hd__clkbuf_16 _19309_ (.A(_05185_),
    .X(_06605_));
 sky130_fd_sc_hd__nand2_8 _19310_ (.A(_06584_),
    .B(\rvcpu.dp.plem.ALUResultM[3] ),
    .Y(_06606_));
 sky130_fd_sc_hd__nor2_4 _19311_ (.A(\rvcpu.dp.plem.ALUResultM[4] ),
    .B(_06606_),
    .Y(_06607_));
 sky130_fd_sc_hd__nand2_8 _19312_ (.A(_06605_),
    .B(_06607_),
    .Y(_06608_));
 sky130_fd_sc_hd__buf_6 _19313_ (.A(_06608_),
    .X(_06609_));
 sky130_fd_sc_hd__buf_8 _19314_ (.A(_06609_),
    .X(_06610_));
 sky130_fd_sc_hd__buf_8 _19315_ (.A(_06610_),
    .X(_06611_));
 sky130_fd_sc_hd__buf_8 _19316_ (.A(_06611_),
    .X(_06612_));
 sky130_fd_sc_hd__buf_6 _19317_ (.A(_06612_),
    .X(_06613_));
 sky130_fd_sc_hd__nand2_4 _19318_ (.A(_06585_),
    .B(\rvcpu.dp.plem.ALUResultM[4] ),
    .Y(_06614_));
 sky130_fd_sc_hd__nor2_8 _19319_ (.A(\rvcpu.dp.plem.ALUResultM[3] ),
    .B(_06614_),
    .Y(_06615_));
 sky130_fd_sc_hd__nand2_4 _19320_ (.A(_06605_),
    .B(_06615_),
    .Y(_06616_));
 sky130_fd_sc_hd__buf_6 _19321_ (.A(_06616_),
    .X(_06617_));
 sky130_fd_sc_hd__clkbuf_8 _19322_ (.A(_06617_),
    .X(_06618_));
 sky130_fd_sc_hd__buf_6 _19323_ (.A(_06618_),
    .X(_06619_));
 sky130_fd_sc_hd__buf_8 _19324_ (.A(_06619_),
    .X(_06620_));
 sky130_fd_sc_hd__buf_4 _19325_ (.A(_06620_),
    .X(_06621_));
 sky130_fd_sc_hd__inv_4 _19326_ (.A(\rvcpu.dp.plem.ALUResultM[4] ),
    .Y(_06622_));
 sky130_fd_sc_hd__nor2_8 _19327_ (.A(_06622_),
    .B(_06606_),
    .Y(_06623_));
 sky130_fd_sc_hd__nand2_4 _19328_ (.A(_06605_),
    .B(_06623_),
    .Y(_06624_));
 sky130_fd_sc_hd__buf_6 _19329_ (.A(_06624_),
    .X(_06625_));
 sky130_fd_sc_hd__clkbuf_8 _19330_ (.A(_06625_),
    .X(_06626_));
 sky130_fd_sc_hd__clkbuf_8 _19331_ (.A(_06626_),
    .X(_06627_));
 sky130_fd_sc_hd__buf_6 _19332_ (.A(_06627_),
    .X(_06628_));
 sky130_fd_sc_hd__buf_8 _19333_ (.A(_06628_),
    .X(_06629_));
 sky130_fd_sc_hd__buf_6 _19334_ (.A(_06629_),
    .X(_06630_));
 sky130_fd_sc_hd__nand2_8 _19335_ (.A(net122),
    .B(_06607_),
    .Y(_06631_));
 sky130_fd_sc_hd__buf_8 _19336_ (.A(_06631_),
    .X(_06632_));
 sky130_fd_sc_hd__buf_6 _19337_ (.A(_06632_),
    .X(_06633_));
 sky130_fd_sc_hd__buf_8 _19338_ (.A(_06633_),
    .X(_06634_));
 sky130_fd_sc_hd__buf_6 _19339_ (.A(_06634_),
    .X(_06635_));
 sky130_fd_sc_hd__buf_6 _19340_ (.A(_06635_),
    .X(_06636_));
 sky130_fd_sc_hd__o22a_1 _19341_ (.A1(\datamem.data_ram[14][16] ),
    .A2(_06630_),
    .B1(_06636_),
    .B2(\datamem.data_ram[11][16] ),
    .X(_06637_));
 sky130_fd_sc_hd__o221a_1 _19342_ (.A1(\datamem.data_ram[10][16] ),
    .A2(_06613_),
    .B1(_06621_),
    .B2(\datamem.data_ram[12][16] ),
    .C1(_06637_),
    .X(_06638_));
 sky130_fd_sc_hd__nand2_8 _19343_ (.A(net122),
    .B(_06584_),
    .Y(_06639_));
 sky130_fd_sc_hd__nor2_8 _19344_ (.A(net1),
    .B(_05371_),
    .Y(_06640_));
 sky130_fd_sc_hd__nor2_8 _19345_ (.A(_06591_),
    .B(_06622_),
    .Y(_06641_));
 sky130_fd_sc_hd__nor2_4 _19346_ (.A(_06640_),
    .B(_06641_),
    .Y(_06642_));
 sky130_fd_sc_hd__nand2_4 _19347_ (.A(_06639_),
    .B(_06642_),
    .Y(_06643_));
 sky130_fd_sc_hd__clkbuf_8 _19348_ (.A(_06643_),
    .X(_06644_));
 sky130_fd_sc_hd__buf_8 _19349_ (.A(_06644_),
    .X(_06645_));
 sky130_fd_sc_hd__buf_8 _19350_ (.A(_06645_),
    .X(_06646_));
 sky130_fd_sc_hd__buf_6 _19351_ (.A(_06646_),
    .X(_06647_));
 sky130_fd_sc_hd__clkbuf_8 _19352_ (.A(_06647_),
    .X(_06648_));
 sky130_fd_sc_hd__buf_6 _19353_ (.A(_06648_),
    .X(_06649_));
 sky130_fd_sc_hd__nor2_2 _19354_ (.A(_05185_),
    .B(net1),
    .Y(_06650_));
 sky130_fd_sc_hd__buf_6 _19355_ (.A(_06650_),
    .X(_06651_));
 sky130_fd_sc_hd__clkbuf_16 _19356_ (.A(_06651_),
    .X(_06652_));
 sky130_fd_sc_hd__nand2_8 _19357_ (.A(_06652_),
    .B(_06642_),
    .Y(_06653_));
 sky130_fd_sc_hd__clkbuf_8 _19358_ (.A(_06653_),
    .X(_06654_));
 sky130_fd_sc_hd__clkbuf_8 _19359_ (.A(_06654_),
    .X(_06655_));
 sky130_fd_sc_hd__buf_4 _19360_ (.A(_06655_),
    .X(_06656_));
 sky130_fd_sc_hd__buf_6 _19361_ (.A(_06656_),
    .X(_06657_));
 sky130_fd_sc_hd__buf_8 _19362_ (.A(_06657_),
    .X(_06658_));
 sky130_fd_sc_hd__clkbuf_8 _19363_ (.A(_06658_),
    .X(_06659_));
 sky130_fd_sc_hd__nand2_8 _19364_ (.A(net122),
    .B(_06615_),
    .Y(_06660_));
 sky130_fd_sc_hd__buf_8 _19365_ (.A(_06660_),
    .X(_06661_));
 sky130_fd_sc_hd__buf_6 _19366_ (.A(_06661_),
    .X(_06662_));
 sky130_fd_sc_hd__buf_8 _19367_ (.A(_06662_),
    .X(_06663_));
 sky130_fd_sc_hd__buf_8 _19368_ (.A(_06663_),
    .X(_06664_));
 sky130_fd_sc_hd__buf_4 _19369_ (.A(_06664_),
    .X(_06665_));
 sky130_fd_sc_hd__clkbuf_16 _19370_ (.A(\rvcpu.dp.plem.ALUResultM[2] ),
    .X(_06666_));
 sky130_fd_sc_hd__nand2_8 _19371_ (.A(_06666_),
    .B(_06623_),
    .Y(_06667_));
 sky130_fd_sc_hd__buf_4 _19372_ (.A(_06667_),
    .X(_06668_));
 sky130_fd_sc_hd__buf_4 _19373_ (.A(_06668_),
    .X(_06669_));
 sky130_fd_sc_hd__clkbuf_8 _19374_ (.A(_06669_),
    .X(_06670_));
 sky130_fd_sc_hd__buf_8 _19375_ (.A(_06670_),
    .X(_06671_));
 sky130_fd_sc_hd__clkbuf_8 _19376_ (.A(_06671_),
    .X(_06672_));
 sky130_fd_sc_hd__o22a_1 _19377_ (.A1(\datamem.data_ram[13][16] ),
    .A2(_06665_),
    .B1(_06672_),
    .B2(\datamem.data_ram[15][16] ),
    .X(_06673_));
 sky130_fd_sc_hd__o221a_1 _19378_ (.A1(\datamem.data_ram[8][16] ),
    .A2(_06649_),
    .B1(_06659_),
    .B2(\datamem.data_ram[9][16] ),
    .C1(_06673_),
    .X(_06674_));
 sky130_fd_sc_hd__nand2_1 _19379_ (.A(_06585_),
    .B(\rvcpu.dp.plem.ALUResultM[5] ),
    .Y(_06675_));
 sky130_fd_sc_hd__buf_8 _19380_ (.A(_06675_),
    .X(_06676_));
 sky130_fd_sc_hd__clkbuf_16 _19381_ (.A(_06676_),
    .X(_06677_));
 sky130_fd_sc_hd__buf_6 _19382_ (.A(_06677_),
    .X(_06678_));
 sky130_fd_sc_hd__buf_8 _19383_ (.A(_06678_),
    .X(_06679_));
 sky130_fd_sc_hd__clkbuf_16 _19384_ (.A(_06679_),
    .X(_06680_));
 sky130_fd_sc_hd__buf_6 _19385_ (.A(_06680_),
    .X(_06681_));
 sky130_fd_sc_hd__buf_8 _19386_ (.A(_06627_),
    .X(_06682_));
 sky130_fd_sc_hd__buf_6 _19387_ (.A(_06682_),
    .X(_06683_));
 sky130_fd_sc_hd__buf_6 _19388_ (.A(_06616_),
    .X(_06684_));
 sky130_fd_sc_hd__clkbuf_8 _19389_ (.A(_06684_),
    .X(_06685_));
 sky130_fd_sc_hd__buf_8 _19390_ (.A(_06685_),
    .X(_06686_));
 sky130_fd_sc_hd__buf_6 _19391_ (.A(_06686_),
    .X(_06687_));
 sky130_fd_sc_hd__buf_6 _19392_ (.A(_06687_),
    .X(_06688_));
 sky130_fd_sc_hd__clkbuf_8 _19393_ (.A(_06608_),
    .X(_06689_));
 sky130_fd_sc_hd__buf_6 _19394_ (.A(_06689_),
    .X(_06690_));
 sky130_fd_sc_hd__buf_6 _19395_ (.A(_06690_),
    .X(_06691_));
 sky130_fd_sc_hd__buf_8 _19396_ (.A(_06691_),
    .X(_06692_));
 sky130_fd_sc_hd__o22a_1 _19397_ (.A1(\datamem.data_ram[2][16] ),
    .A2(_06692_),
    .B1(_06635_),
    .B2(\datamem.data_ram[3][16] ),
    .X(_06693_));
 sky130_fd_sc_hd__o221a_1 _19398_ (.A1(\datamem.data_ram[6][16] ),
    .A2(_06683_),
    .B1(_06688_),
    .B2(\datamem.data_ram[4][16] ),
    .C1(_06693_),
    .X(_06694_));
 sky130_fd_sc_hd__buf_6 _19399_ (.A(_06645_),
    .X(_06695_));
 sky130_fd_sc_hd__clkbuf_8 _19400_ (.A(_06695_),
    .X(_06696_));
 sky130_fd_sc_hd__buf_6 _19401_ (.A(_06696_),
    .X(_06697_));
 sky130_fd_sc_hd__clkbuf_8 _19402_ (.A(_06697_),
    .X(_06698_));
 sky130_fd_sc_hd__clkbuf_8 _19403_ (.A(_06655_),
    .X(_06699_));
 sky130_fd_sc_hd__buf_6 _19404_ (.A(_06699_),
    .X(_06700_));
 sky130_fd_sc_hd__clkbuf_8 _19405_ (.A(_06700_),
    .X(_06701_));
 sky130_fd_sc_hd__buf_6 _19406_ (.A(_06662_),
    .X(_06702_));
 sky130_fd_sc_hd__buf_6 _19407_ (.A(_06702_),
    .X(_06703_));
 sky130_fd_sc_hd__buf_8 _19408_ (.A(_06667_),
    .X(_06704_));
 sky130_fd_sc_hd__clkbuf_8 _19409_ (.A(_06704_),
    .X(_06705_));
 sky130_fd_sc_hd__clkbuf_8 _19410_ (.A(_06705_),
    .X(_06706_));
 sky130_fd_sc_hd__buf_6 _19411_ (.A(_06706_),
    .X(_06707_));
 sky130_fd_sc_hd__o22a_1 _19412_ (.A1(\datamem.data_ram[5][16] ),
    .A2(_06703_),
    .B1(_06707_),
    .B2(\datamem.data_ram[7][16] ),
    .X(_06708_));
 sky130_fd_sc_hd__o221a_1 _19413_ (.A1(\datamem.data_ram[0][16] ),
    .A2(_06698_),
    .B1(_06701_),
    .B2(\datamem.data_ram[1][16] ),
    .C1(_06708_),
    .X(_06709_));
 sky130_fd_sc_hd__and3_1 _19414_ (.A(_06681_),
    .B(_06694_),
    .C(_06709_),
    .X(_06710_));
 sky130_fd_sc_hd__a31o_1 _19415_ (.A1(_06604_),
    .A2(_06638_),
    .A3(_06674_),
    .B1(_06710_),
    .X(_06711_));
 sky130_fd_sc_hd__buf_4 _19416_ (.A(_06594_),
    .X(_06712_));
 sky130_fd_sc_hd__buf_6 _19417_ (.A(_06712_),
    .X(_06713_));
 sky130_fd_sc_hd__buf_8 _19418_ (.A(_06592_),
    .X(_06714_));
 sky130_fd_sc_hd__buf_8 _19419_ (.A(_06714_),
    .X(_06715_));
 sky130_fd_sc_hd__clkbuf_8 _19420_ (.A(_06715_),
    .X(_06716_));
 sky130_fd_sc_hd__buf_6 _19421_ (.A(_06625_),
    .X(_06717_));
 sky130_fd_sc_hd__buf_4 _19422_ (.A(_06717_),
    .X(_06718_));
 sky130_fd_sc_hd__buf_8 _19423_ (.A(_06718_),
    .X(_06719_));
 sky130_fd_sc_hd__o22a_1 _19424_ (.A1(\datamem.data_ram[38][16] ),
    .A2(_06719_),
    .B1(_06687_),
    .B2(\datamem.data_ram[36][16] ),
    .X(_06720_));
 sky130_fd_sc_hd__buf_6 _19425_ (.A(_06660_),
    .X(_06721_));
 sky130_fd_sc_hd__buf_6 _19426_ (.A(_06721_),
    .X(_06722_));
 sky130_fd_sc_hd__clkbuf_8 _19427_ (.A(_06722_),
    .X(_06723_));
 sky130_fd_sc_hd__clkbuf_8 _19428_ (.A(_06723_),
    .X(_06724_));
 sky130_fd_sc_hd__clkbuf_8 _19429_ (.A(_06668_),
    .X(_06725_));
 sky130_fd_sc_hd__buf_6 _19430_ (.A(_06725_),
    .X(_06726_));
 sky130_fd_sc_hd__o22a_1 _19431_ (.A1(\datamem.data_ram[39][16] ),
    .A2(_06726_),
    .B1(_06699_),
    .B2(\datamem.data_ram[33][16] ),
    .X(_06727_));
 sky130_fd_sc_hd__buf_6 _19432_ (.A(_06690_),
    .X(_06728_));
 sky130_fd_sc_hd__clkbuf_8 _19433_ (.A(_06631_),
    .X(_06729_));
 sky130_fd_sc_hd__clkbuf_8 _19434_ (.A(_06729_),
    .X(_06730_));
 sky130_fd_sc_hd__buf_6 _19435_ (.A(_06730_),
    .X(_06731_));
 sky130_fd_sc_hd__buf_8 _19436_ (.A(_06676_),
    .X(_06732_));
 sky130_fd_sc_hd__buf_8 _19437_ (.A(_06732_),
    .X(_06733_));
 sky130_fd_sc_hd__o221a_1 _19438_ (.A1(\datamem.data_ram[34][16] ),
    .A2(_06728_),
    .B1(_06731_),
    .B2(\datamem.data_ram[35][16] ),
    .C1(_06733_),
    .X(_06734_));
 sky130_fd_sc_hd__o211a_1 _19439_ (.A1(\datamem.data_ram[37][16] ),
    .A2(_06724_),
    .B1(_06727_),
    .C1(_06734_),
    .X(_06735_));
 sky130_fd_sc_hd__o211a_1 _19440_ (.A1(\datamem.data_ram[32][16] ),
    .A2(_06698_),
    .B1(_06720_),
    .C1(_06735_),
    .X(_06736_));
 sky130_fd_sc_hd__clkbuf_8 _19441_ (.A(_06730_),
    .X(_06737_));
 sky130_fd_sc_hd__buf_6 _19442_ (.A(_06737_),
    .X(_06738_));
 sky130_fd_sc_hd__buf_6 _19443_ (.A(_06738_),
    .X(_06739_));
 sky130_fd_sc_hd__o22a_1 _19444_ (.A1(\datamem.data_ram[44][16] ),
    .A2(_06687_),
    .B1(_06700_),
    .B2(\datamem.data_ram[41][16] ),
    .X(_06740_));
 sky130_fd_sc_hd__buf_8 _19445_ (.A(_06599_),
    .X(_06741_));
 sky130_fd_sc_hd__buf_8 _19446_ (.A(_06741_),
    .X(_06742_));
 sky130_fd_sc_hd__clkbuf_8 _19447_ (.A(_06624_),
    .X(_06743_));
 sky130_fd_sc_hd__buf_6 _19448_ (.A(_06743_),
    .X(_06744_));
 sky130_fd_sc_hd__o22a_1 _19449_ (.A1(\datamem.data_ram[46][16] ),
    .A2(_06744_),
    .B1(_06695_),
    .B2(\datamem.data_ram[40][16] ),
    .X(_06745_));
 sky130_fd_sc_hd__o221a_1 _19450_ (.A1(\datamem.data_ram[42][16] ),
    .A2(_06728_),
    .B1(_06726_),
    .B2(\datamem.data_ram[47][16] ),
    .C1(_06745_),
    .X(_06746_));
 sky130_fd_sc_hd__o211a_1 _19451_ (.A1(\datamem.data_ram[45][16] ),
    .A2(_06724_),
    .B1(_06742_),
    .C1(_06746_),
    .X(_06747_));
 sky130_fd_sc_hd__o211a_1 _19452_ (.A1(\datamem.data_ram[43][16] ),
    .A2(_06739_),
    .B1(_06740_),
    .C1(_06747_),
    .X(_06748_));
 sky130_fd_sc_hd__or3_1 _19453_ (.A(_06716_),
    .B(_06736_),
    .C(_06748_),
    .X(_06749_));
 sky130_fd_sc_hd__nand2_8 _19454_ (.A(_06585_),
    .B(\rvcpu.dp.plem.ALUResultM[6] ),
    .Y(_06750_));
 sky130_fd_sc_hd__buf_8 _19455_ (.A(_06750_),
    .X(_06751_));
 sky130_fd_sc_hd__buf_8 _19456_ (.A(_06751_),
    .X(_06752_));
 sky130_fd_sc_hd__buf_6 _19457_ (.A(_06752_),
    .X(_06753_));
 sky130_fd_sc_hd__buf_8 _19458_ (.A(_06728_),
    .X(_06754_));
 sky130_fd_sc_hd__o22a_1 _19459_ (.A1(\datamem.data_ram[58][16] ),
    .A2(_06754_),
    .B1(_06671_),
    .B2(\datamem.data_ram[63][16] ),
    .X(_06755_));
 sky130_fd_sc_hd__o22a_1 _19460_ (.A1(\datamem.data_ram[61][16] ),
    .A2(_06722_),
    .B1(_06655_),
    .B2(\datamem.data_ram[57][16] ),
    .X(_06756_));
 sky130_fd_sc_hd__o221a_1 _19461_ (.A1(\datamem.data_ram[56][16] ),
    .A2(_06696_),
    .B1(_06686_),
    .B2(\datamem.data_ram[60][16] ),
    .C1(_06756_),
    .X(_06757_));
 sky130_fd_sc_hd__o211a_1 _19462_ (.A1(\datamem.data_ram[62][16] ),
    .A2(_06719_),
    .B1(_06742_),
    .C1(_06757_),
    .X(_06758_));
 sky130_fd_sc_hd__o211a_1 _19463_ (.A1(\datamem.data_ram[59][16] ),
    .A2(_06739_),
    .B1(_06755_),
    .C1(_06758_),
    .X(_06759_));
 sky130_fd_sc_hd__buf_6 _19464_ (.A(_06725_),
    .X(_06760_));
 sky130_fd_sc_hd__clkbuf_8 _19465_ (.A(_06760_),
    .X(_06761_));
 sky130_fd_sc_hd__o22a_1 _19466_ (.A1(\datamem.data_ram[48][16] ),
    .A2(_06697_),
    .B1(_06761_),
    .B2(\datamem.data_ram[55][16] ),
    .X(_06762_));
 sky130_fd_sc_hd__buf_6 _19467_ (.A(_06744_),
    .X(_06763_));
 sky130_fd_sc_hd__clkbuf_8 _19468_ (.A(_06763_),
    .X(_06764_));
 sky130_fd_sc_hd__buf_6 _19469_ (.A(_06684_),
    .X(_06765_));
 sky130_fd_sc_hd__buf_6 _19470_ (.A(_06765_),
    .X(_06766_));
 sky130_fd_sc_hd__o22a_1 _19471_ (.A1(\datamem.data_ram[52][16] ),
    .A2(_06766_),
    .B1(_06699_),
    .B2(\datamem.data_ram[49][16] ),
    .X(_06767_));
 sky130_fd_sc_hd__clkbuf_8 _19472_ (.A(_06722_),
    .X(_06768_));
 sky130_fd_sc_hd__buf_8 _19473_ (.A(_06732_),
    .X(_06769_));
 sky130_fd_sc_hd__o221a_1 _19474_ (.A1(\datamem.data_ram[50][16] ),
    .A2(_06728_),
    .B1(_06768_),
    .B2(\datamem.data_ram[53][16] ),
    .C1(_06769_),
    .X(_06770_));
 sky130_fd_sc_hd__o211a_1 _19475_ (.A1(\datamem.data_ram[54][16] ),
    .A2(_06764_),
    .B1(_06767_),
    .C1(_06770_),
    .X(_06771_));
 sky130_fd_sc_hd__o211a_1 _19476_ (.A1(\datamem.data_ram[51][16] ),
    .A2(_06739_),
    .B1(_06762_),
    .C1(_06771_),
    .X(_06772_));
 sky130_fd_sc_hd__or3_2 _19477_ (.A(_06753_),
    .B(_06759_),
    .C(_06772_),
    .X(_06773_));
 sky130_fd_sc_hd__or2_1 _19478_ (.A(\datamem.data_ram[19][16] ),
    .B(_06636_),
    .X(_06774_));
 sky130_fd_sc_hd__o22a_1 _19479_ (.A1(\datamem.data_ram[21][16] ),
    .A2(_06665_),
    .B1(_06621_),
    .B2(\datamem.data_ram[20][16] ),
    .X(_06775_));
 sky130_fd_sc_hd__buf_8 _19480_ (.A(_06679_),
    .X(_06776_));
 sky130_fd_sc_hd__buf_8 _19481_ (.A(_06776_),
    .X(_06777_));
 sky130_fd_sc_hd__clkbuf_8 _19482_ (.A(_06646_),
    .X(_06778_));
 sky130_fd_sc_hd__buf_6 _19483_ (.A(_06778_),
    .X(_06779_));
 sky130_fd_sc_hd__buf_8 _19484_ (.A(_06654_),
    .X(_06780_));
 sky130_fd_sc_hd__buf_6 _19485_ (.A(_06780_),
    .X(_06781_));
 sky130_fd_sc_hd__buf_8 _19486_ (.A(_06781_),
    .X(_06782_));
 sky130_fd_sc_hd__buf_8 _19487_ (.A(_06782_),
    .X(_06783_));
 sky130_fd_sc_hd__buf_8 _19488_ (.A(_06670_),
    .X(_06784_));
 sky130_fd_sc_hd__o22a_1 _19489_ (.A1(\datamem.data_ram[18][16] ),
    .A2(_06611_),
    .B1(_06784_),
    .B2(\datamem.data_ram[23][16] ),
    .X(_06785_));
 sky130_fd_sc_hd__o221a_1 _19490_ (.A1(\datamem.data_ram[16][16] ),
    .A2(_06779_),
    .B1(_06783_),
    .B2(\datamem.data_ram[17][16] ),
    .C1(_06785_),
    .X(_06786_));
 sky130_fd_sc_hd__o211a_1 _19491_ (.A1(\datamem.data_ram[22][16] ),
    .A2(_06630_),
    .B1(_06777_),
    .C1(_06786_),
    .X(_06787_));
 sky130_fd_sc_hd__o22a_1 _19492_ (.A1(\datamem.data_ram[30][16] ),
    .A2(_06629_),
    .B1(_06620_),
    .B2(\datamem.data_ram[28][16] ),
    .X(_06788_));
 sky130_fd_sc_hd__clkbuf_8 _19493_ (.A(_06655_),
    .X(_06789_));
 sky130_fd_sc_hd__buf_8 _19494_ (.A(_06789_),
    .X(_06790_));
 sky130_fd_sc_hd__o22a_1 _19495_ (.A1(\datamem.data_ram[24][16] ),
    .A2(_06647_),
    .B1(_06790_),
    .B2(\datamem.data_ram[25][16] ),
    .X(_06791_));
 sky130_fd_sc_hd__o221a_1 _19496_ (.A1(\datamem.data_ram[26][16] ),
    .A2(_06611_),
    .B1(_06784_),
    .B2(\datamem.data_ram[31][16] ),
    .C1(_06601_),
    .X(_06792_));
 sky130_fd_sc_hd__o211a_1 _19497_ (.A1(\datamem.data_ram[29][16] ),
    .A2(_06664_),
    .B1(_06791_),
    .C1(_06792_),
    .X(_06793_));
 sky130_fd_sc_hd__o211a_1 _19498_ (.A1(\datamem.data_ram[27][16] ),
    .A2(_06636_),
    .B1(_06788_),
    .C1(_06793_),
    .X(_06794_));
 sky130_fd_sc_hd__a31o_1 _19499_ (.A1(_06774_),
    .A2(_06775_),
    .A3(_06787_),
    .B1(_06794_),
    .X(_06795_));
 sky130_fd_sc_hd__nor2_8 _19500_ (.A(\rvcpu.dp.plem.ALUResultM[7] ),
    .B(_06750_),
    .Y(_06796_));
 sky130_fd_sc_hd__buf_8 _19501_ (.A(_06796_),
    .X(_06797_));
 sky130_fd_sc_hd__a32o_1 _19502_ (.A1(_06713_),
    .A2(_06749_),
    .A3(_06773_),
    .B1(_06795_),
    .B2(_06797_),
    .X(_06798_));
 sky130_fd_sc_hd__a21oi_4 _19503_ (.A1(_06596_),
    .A2(_06711_),
    .B1(_06798_),
    .Y(_06799_));
 sky130_fd_sc_hd__o22a_1 _19504_ (.A1(\datamem.data_ram[53][24] ),
    .A2(_06723_),
    .B1(_06731_),
    .B2(\datamem.data_ram[51][24] ),
    .X(_06800_));
 sky130_fd_sc_hd__o221a_1 _19505_ (.A1(\datamem.data_ram[54][24] ),
    .A2(_06682_),
    .B1(_06790_),
    .B2(\datamem.data_ram[49][24] ),
    .C1(_06800_),
    .X(_06801_));
 sky130_fd_sc_hd__clkbuf_8 _19506_ (.A(_06689_),
    .X(_06802_));
 sky130_fd_sc_hd__clkbuf_8 _19507_ (.A(_06802_),
    .X(_06803_));
 sky130_fd_sc_hd__clkbuf_8 _19508_ (.A(_06803_),
    .X(_06804_));
 sky130_fd_sc_hd__clkbuf_8 _19509_ (.A(_06685_),
    .X(_06805_));
 sky130_fd_sc_hd__buf_6 _19510_ (.A(_06805_),
    .X(_06806_));
 sky130_fd_sc_hd__buf_6 _19511_ (.A(_06695_),
    .X(_06807_));
 sky130_fd_sc_hd__o22a_1 _19512_ (.A1(\datamem.data_ram[48][24] ),
    .A2(_06807_),
    .B1(_06726_),
    .B2(\datamem.data_ram[55][24] ),
    .X(_06808_));
 sky130_fd_sc_hd__o221a_1 _19513_ (.A1(\datamem.data_ram[50][24] ),
    .A2(_06804_),
    .B1(_06806_),
    .B2(\datamem.data_ram[52][24] ),
    .C1(_06808_),
    .X(_06809_));
 sky130_fd_sc_hd__buf_8 _19514_ (.A(_06741_),
    .X(_06810_));
 sky130_fd_sc_hd__buf_4 _19515_ (.A(_06644_),
    .X(_06811_));
 sky130_fd_sc_hd__clkbuf_8 _19516_ (.A(_06729_),
    .X(_06812_));
 sky130_fd_sc_hd__o22a_1 _19517_ (.A1(\datamem.data_ram[56][24] ),
    .A2(_06811_),
    .B1(_06812_),
    .B2(\datamem.data_ram[59][24] ),
    .X(_06813_));
 sky130_fd_sc_hd__o221a_1 _19518_ (.A1(\datamem.data_ram[63][24] ),
    .A2(_06670_),
    .B1(_06781_),
    .B2(\datamem.data_ram[57][24] ),
    .C1(_06813_),
    .X(_06814_));
 sky130_fd_sc_hd__buf_6 _19519_ (.A(_06661_),
    .X(_06815_));
 sky130_fd_sc_hd__o22a_1 _19520_ (.A1(\datamem.data_ram[62][24] ),
    .A2(_06626_),
    .B1(_06685_),
    .B2(\datamem.data_ram[60][24] ),
    .X(_06816_));
 sky130_fd_sc_hd__o221a_1 _19521_ (.A1(\datamem.data_ram[58][24] ),
    .A2(_06803_),
    .B1(_06815_),
    .B2(\datamem.data_ram[61][24] ),
    .C1(_06816_),
    .X(_06817_));
 sky130_fd_sc_hd__and3_1 _19522_ (.A(_06810_),
    .B(_06814_),
    .C(_06817_),
    .X(_06818_));
 sky130_fd_sc_hd__a31o_1 _19523_ (.A1(_06776_),
    .A2(_06801_),
    .A3(_06809_),
    .B1(_06818_),
    .X(_06819_));
 sky130_fd_sc_hd__buf_6 _19524_ (.A(_06644_),
    .X(_06820_));
 sky130_fd_sc_hd__buf_8 _19525_ (.A(_06820_),
    .X(_06821_));
 sky130_fd_sc_hd__o22a_1 _19526_ (.A1(\datamem.data_ram[40][24] ),
    .A2(_06821_),
    .B1(_06805_),
    .B2(\datamem.data_ram[44][24] ),
    .X(_06822_));
 sky130_fd_sc_hd__clkbuf_8 _19527_ (.A(_06722_),
    .X(_06823_));
 sky130_fd_sc_hd__o22a_1 _19528_ (.A1(\datamem.data_ram[42][24] ),
    .A2(_06802_),
    .B1(_06669_),
    .B2(\datamem.data_ram[47][24] ),
    .X(_06824_));
 sky130_fd_sc_hd__o221a_1 _19529_ (.A1(\datamem.data_ram[46][24] ),
    .A2(_06626_),
    .B1(_06812_),
    .B2(\datamem.data_ram[43][24] ),
    .C1(_06599_),
    .X(_06825_));
 sky130_fd_sc_hd__o211a_1 _19530_ (.A1(\datamem.data_ram[45][24] ),
    .A2(_06823_),
    .B1(_06824_),
    .C1(_06825_),
    .X(_06826_));
 sky130_fd_sc_hd__o211a_1 _19531_ (.A1(\datamem.data_ram[41][24] ),
    .A2(_06790_),
    .B1(_06822_),
    .C1(_06826_),
    .X(_06827_));
 sky130_fd_sc_hd__clkbuf_8 _19532_ (.A(_06812_),
    .X(_06828_));
 sky130_fd_sc_hd__buf_6 _19533_ (.A(_06828_),
    .X(_06829_));
 sky130_fd_sc_hd__o22a_1 _19534_ (.A1(\datamem.data_ram[38][24] ),
    .A2(_06718_),
    .B1(_06686_),
    .B2(\datamem.data_ram[36][24] ),
    .X(_06830_));
 sky130_fd_sc_hd__o22a_1 _19535_ (.A1(\datamem.data_ram[34][24] ),
    .A2(_06689_),
    .B1(_06668_),
    .B2(\datamem.data_ram[39][24] ),
    .X(_06831_));
 sky130_fd_sc_hd__o221a_1 _19536_ (.A1(\datamem.data_ram[32][24] ),
    .A2(_06811_),
    .B1(_06655_),
    .B2(\datamem.data_ram[33][24] ),
    .C1(_06831_),
    .X(_06832_));
 sky130_fd_sc_hd__o211a_1 _19537_ (.A1(\datamem.data_ram[37][24] ),
    .A2(_06823_),
    .B1(_06733_),
    .C1(_06832_),
    .X(_06833_));
 sky130_fd_sc_hd__o211a_1 _19538_ (.A1(\datamem.data_ram[35][24] ),
    .A2(_06829_),
    .B1(_06830_),
    .C1(_06833_),
    .X(_06834_));
 sky130_fd_sc_hd__or3_1 _19539_ (.A(_06827_),
    .B(_06714_),
    .C(_06834_),
    .X(_06835_));
 sky130_fd_sc_hd__o211a_1 _19540_ (.A1(_06753_),
    .A2(_06819_),
    .B1(_06712_),
    .C1(_06835_),
    .X(_06836_));
 sky130_fd_sc_hd__buf_6 _19541_ (.A(_06807_),
    .X(_06837_));
 sky130_fd_sc_hd__o22a_1 _19542_ (.A1(\datamem.data_ram[24][24] ),
    .A2(_06837_),
    .B1(_06806_),
    .B2(\datamem.data_ram[28][24] ),
    .X(_06838_));
 sky130_fd_sc_hd__o22a_1 _19543_ (.A1(\datamem.data_ram[30][24] ),
    .A2(_06717_),
    .B1(_06812_),
    .B2(\datamem.data_ram[27][24] ),
    .X(_06839_));
 sky130_fd_sc_hd__o221a_1 _19544_ (.A1(\datamem.data_ram[29][24] ),
    .A2(_06815_),
    .B1(_06670_),
    .B2(\datamem.data_ram[31][24] ),
    .C1(_06839_),
    .X(_06840_));
 sky130_fd_sc_hd__o211a_1 _19545_ (.A1(\datamem.data_ram[25][24] ),
    .A2(_06790_),
    .B1(_06840_),
    .C1(_06810_),
    .X(_06841_));
 sky130_fd_sc_hd__o211a_1 _19546_ (.A1(\datamem.data_ram[26][24] ),
    .A2(_06612_),
    .B1(_06838_),
    .C1(_06841_),
    .X(_06842_));
 sky130_fd_sc_hd__o22a_1 _19547_ (.A1(\datamem.data_ram[21][24] ),
    .A2(_06724_),
    .B1(_06671_),
    .B2(\datamem.data_ram[23][24] ),
    .X(_06843_));
 sky130_fd_sc_hd__o22a_1 _19548_ (.A1(\datamem.data_ram[22][24] ),
    .A2(_06718_),
    .B1(_06696_),
    .B2(\datamem.data_ram[16][24] ),
    .X(_06844_));
 sky130_fd_sc_hd__o221a_1 _19549_ (.A1(\datamem.data_ram[18][24] ),
    .A2(_06803_),
    .B1(_06731_),
    .B2(\datamem.data_ram[19][24] ),
    .C1(_06733_),
    .X(_06845_));
 sky130_fd_sc_hd__o211a_1 _19550_ (.A1(\datamem.data_ram[20][24] ),
    .A2(_06687_),
    .B1(_06844_),
    .C1(_06845_),
    .X(_06846_));
 sky130_fd_sc_hd__o211a_1 _19551_ (.A1(\datamem.data_ram[17][24] ),
    .A2(_06658_),
    .B1(_06843_),
    .C1(_06846_),
    .X(_06847_));
 sky130_fd_sc_hd__o22a_1 _19552_ (.A1(\datamem.data_ram[13][24] ),
    .A2(_06823_),
    .B1(_06789_),
    .B2(\datamem.data_ram[9][24] ),
    .X(_06848_));
 sky130_fd_sc_hd__o22a_1 _19553_ (.A1(\datamem.data_ram[14][24] ),
    .A2(_06625_),
    .B1(_06689_),
    .B2(\datamem.data_ram[10][24] ),
    .X(_06849_));
 sky130_fd_sc_hd__o221a_1 _19554_ (.A1(\datamem.data_ram[8][24] ),
    .A2(_06820_),
    .B1(_06669_),
    .B2(\datamem.data_ram[15][24] ),
    .C1(_06849_),
    .X(_06850_));
 sky130_fd_sc_hd__buf_8 _19555_ (.A(_06599_),
    .X(_06851_));
 sky130_fd_sc_hd__o211a_1 _19556_ (.A1(\datamem.data_ram[12][24] ),
    .A2(_06805_),
    .B1(_06850_),
    .C1(_06851_),
    .X(_06852_));
 sky130_fd_sc_hd__o211a_1 _19557_ (.A1(\datamem.data_ram[11][24] ),
    .A2(_06829_),
    .B1(_06848_),
    .C1(_06852_),
    .X(_06853_));
 sky130_fd_sc_hd__o22a_1 _19558_ (.A1(\datamem.data_ram[6][24] ),
    .A2(_06718_),
    .B1(_06686_),
    .B2(\datamem.data_ram[4][24] ),
    .X(_06854_));
 sky130_fd_sc_hd__o22a_1 _19559_ (.A1(\datamem.data_ram[0][24] ),
    .A2(_06811_),
    .B1(_06669_),
    .B2(\datamem.data_ram[7][24] ),
    .X(_06855_));
 sky130_fd_sc_hd__o221a_1 _19560_ (.A1(\datamem.data_ram[2][24] ),
    .A2(_06802_),
    .B1(_06655_),
    .B2(\datamem.data_ram[1][24] ),
    .C1(_06732_),
    .X(_06856_));
 sky130_fd_sc_hd__o211a_1 _19561_ (.A1(\datamem.data_ram[5][24] ),
    .A2(_06823_),
    .B1(_06855_),
    .C1(_06856_),
    .X(_06857_));
 sky130_fd_sc_hd__o211a_1 _19562_ (.A1(\datamem.data_ram[3][24] ),
    .A2(_06829_),
    .B1(_06854_),
    .C1(_06857_),
    .X(_06858_));
 sky130_fd_sc_hd__or3_1 _19563_ (.A(_06714_),
    .B(_06853_),
    .C(_06858_),
    .X(_06859_));
 sky130_fd_sc_hd__nand2_8 _19564_ (.A(_06585_),
    .B(\rvcpu.dp.plem.ALUResultM[7] ),
    .Y(_06860_));
 sky130_fd_sc_hd__o311a_1 _19565_ (.A1(_06752_),
    .A2(_06842_),
    .A3(_06847_),
    .B1(_06859_),
    .C1(_06860_),
    .X(_06861_));
 sky130_fd_sc_hd__nor2_4 _19566_ (.A(_06836_),
    .B(_06861_),
    .Y(_06862_));
 sky130_fd_sc_hd__buf_8 _19567_ (.A(_06829_),
    .X(_06863_));
 sky130_fd_sc_hd__or2_1 _19568_ (.A(\datamem.data_ram[3][8] ),
    .B(_06863_),
    .X(_06864_));
 sky130_fd_sc_hd__clkbuf_8 _19569_ (.A(_06724_),
    .X(_06865_));
 sky130_fd_sc_hd__o22a_1 _19570_ (.A1(\datamem.data_ram[5][8] ),
    .A2(_06865_),
    .B1(_06672_),
    .B2(\datamem.data_ram[7][8] ),
    .X(_06866_));
 sky130_fd_sc_hd__o22a_1 _19571_ (.A1(\datamem.data_ram[6][8] ),
    .A2(_06718_),
    .B1(_06789_),
    .B2(\datamem.data_ram[1][8] ),
    .X(_06867_));
 sky130_fd_sc_hd__o221a_1 _19572_ (.A1(\datamem.data_ram[2][8] ),
    .A2(_06804_),
    .B1(_06837_),
    .B2(\datamem.data_ram[0][8] ),
    .C1(_06867_),
    .X(_06868_));
 sky130_fd_sc_hd__o211a_1 _19573_ (.A1(\datamem.data_ram[4][8] ),
    .A2(_06620_),
    .B1(_06868_),
    .C1(_06776_),
    .X(_06869_));
 sky130_fd_sc_hd__o22a_1 _19574_ (.A1(\datamem.data_ram[13][8] ),
    .A2(_06724_),
    .B1(_06837_),
    .B2(\datamem.data_ram[8][8] ),
    .X(_06870_));
 sky130_fd_sc_hd__o22a_1 _19575_ (.A1(\datamem.data_ram[12][8] ),
    .A2(_06686_),
    .B1(_06656_),
    .B2(\datamem.data_ram[9][8] ),
    .X(_06871_));
 sky130_fd_sc_hd__o221a_1 _19576_ (.A1(\datamem.data_ram[11][8] ),
    .A2(_06731_),
    .B1(_06726_),
    .B2(\datamem.data_ram[15][8] ),
    .C1(_06741_),
    .X(_06872_));
 sky130_fd_sc_hd__o211a_1 _19577_ (.A1(\datamem.data_ram[10][8] ),
    .A2(_06754_),
    .B1(_06871_),
    .C1(_06872_),
    .X(_06873_));
 sky130_fd_sc_hd__o211a_1 _19578_ (.A1(\datamem.data_ram[14][8] ),
    .A2(_06683_),
    .B1(_06870_),
    .C1(_06873_),
    .X(_06874_));
 sky130_fd_sc_hd__a31o_1 _19579_ (.A1(_06864_),
    .A2(_06866_),
    .A3(_06869_),
    .B1(_06874_),
    .X(_06875_));
 sky130_fd_sc_hd__o22a_1 _19580_ (.A1(\datamem.data_ram[32][8] ),
    .A2(_06821_),
    .B1(_06618_),
    .B2(\datamem.data_ram[36][8] ),
    .X(_06876_));
 sky130_fd_sc_hd__o22a_1 _19581_ (.A1(\datamem.data_ram[35][8] ),
    .A2(_06632_),
    .B1(_06669_),
    .B2(\datamem.data_ram[39][8] ),
    .X(_06877_));
 sky130_fd_sc_hd__o221a_1 _19582_ (.A1(\datamem.data_ram[34][8] ),
    .A2(_06609_),
    .B1(_06780_),
    .B2(\datamem.data_ram[33][8] ),
    .C1(_06677_),
    .X(_06878_));
 sky130_fd_sc_hd__o211a_1 _19583_ (.A1(\datamem.data_ram[37][8] ),
    .A2(_06815_),
    .B1(_06877_),
    .C1(_06878_),
    .X(_06879_));
 sky130_fd_sc_hd__o211a_1 _19584_ (.A1(\datamem.data_ram[38][8] ),
    .A2(_06628_),
    .B1(_06876_),
    .C1(_06879_),
    .X(_06880_));
 sky130_fd_sc_hd__o22a_1 _19585_ (.A1(\datamem.data_ram[44][8] ),
    .A2(_06618_),
    .B1(_06781_),
    .B2(\datamem.data_ram[41][8] ),
    .X(_06881_));
 sky130_fd_sc_hd__o22a_1 _19586_ (.A1(\datamem.data_ram[42][8] ),
    .A2(_06689_),
    .B1(_06644_),
    .B2(\datamem.data_ram[40][8] ),
    .X(_06882_));
 sky130_fd_sc_hd__o221a_1 _19587_ (.A1(\datamem.data_ram[46][8] ),
    .A2(_06743_),
    .B1(_06661_),
    .B2(\datamem.data_ram[45][8] ),
    .C1(_06882_),
    .X(_06883_));
 sky130_fd_sc_hd__o211a_1 _19588_ (.A1(\datamem.data_ram[47][8] ),
    .A2(_06670_),
    .B1(_06883_),
    .C1(_06851_),
    .X(_06884_));
 sky130_fd_sc_hd__o211a_1 _19589_ (.A1(\datamem.data_ram[43][8] ),
    .A2(_06634_),
    .B1(_06881_),
    .C1(_06884_),
    .X(_06885_));
 sky130_fd_sc_hd__or3_1 _19590_ (.A(_06714_),
    .B(_06880_),
    .C(_06885_),
    .X(_06886_));
 sky130_fd_sc_hd__o22a_1 _19591_ (.A1(\datamem.data_ram[58][8] ),
    .A2(_06610_),
    .B1(_06821_),
    .B2(\datamem.data_ram[56][8] ),
    .X(_06887_));
 sky130_fd_sc_hd__o22a_1 _19592_ (.A1(\datamem.data_ram[61][8] ),
    .A2(_06721_),
    .B1(_06654_),
    .B2(\datamem.data_ram[57][8] ),
    .X(_06888_));
 sky130_fd_sc_hd__o221a_1 _19593_ (.A1(\datamem.data_ram[62][8] ),
    .A2(_06743_),
    .B1(_06617_),
    .B2(\datamem.data_ram[60][8] ),
    .C1(_06888_),
    .X(_06889_));
 sky130_fd_sc_hd__o211a_1 _19594_ (.A1(\datamem.data_ram[63][8] ),
    .A2(_06670_),
    .B1(_06889_),
    .C1(_06851_),
    .X(_06890_));
 sky130_fd_sc_hd__o211a_1 _19595_ (.A1(\datamem.data_ram[59][8] ),
    .A2(_06634_),
    .B1(_06887_),
    .C1(_06890_),
    .X(_06891_));
 sky130_fd_sc_hd__o22a_1 _19596_ (.A1(\datamem.data_ram[53][8] ),
    .A2(_06815_),
    .B1(_06670_),
    .B2(\datamem.data_ram[55][8] ),
    .X(_06892_));
 sky130_fd_sc_hd__o22a_1 _19597_ (.A1(\datamem.data_ram[54][8] ),
    .A2(_06626_),
    .B1(_06811_),
    .B2(\datamem.data_ram[48][8] ),
    .X(_06893_));
 sky130_fd_sc_hd__o221a_1 _19598_ (.A1(\datamem.data_ram[50][8] ),
    .A2(_06609_),
    .B1(_06780_),
    .B2(\datamem.data_ram[49][8] ),
    .C1(_06677_),
    .X(_06894_));
 sky130_fd_sc_hd__o211a_1 _19599_ (.A1(\datamem.data_ram[52][8] ),
    .A2(_06805_),
    .B1(_06893_),
    .C1(_06894_),
    .X(_06895_));
 sky130_fd_sc_hd__o211a_1 _19600_ (.A1(\datamem.data_ram[51][8] ),
    .A2(_06634_),
    .B1(_06892_),
    .C1(_06895_),
    .X(_06896_));
 sky130_fd_sc_hd__or3_1 _19601_ (.A(_06751_),
    .B(_06891_),
    .C(_06896_),
    .X(_06897_));
 sky130_fd_sc_hd__o22a_1 _19602_ (.A1(\datamem.data_ram[16][8] ),
    .A2(_06696_),
    .B1(_06731_),
    .B2(\datamem.data_ram[19][8] ),
    .X(_06898_));
 sky130_fd_sc_hd__o221a_1 _19603_ (.A1(\datamem.data_ram[18][8] ),
    .A2(_06804_),
    .B1(_06806_),
    .B2(\datamem.data_ram[20][8] ),
    .C1(_06898_),
    .X(_06899_));
 sky130_fd_sc_hd__o22a_1 _19604_ (.A1(\datamem.data_ram[21][8] ),
    .A2(_06723_),
    .B1(_06726_),
    .B2(\datamem.data_ram[23][8] ),
    .X(_06900_));
 sky130_fd_sc_hd__o221a_1 _19605_ (.A1(\datamem.data_ram[22][8] ),
    .A2(_06682_),
    .B1(_06790_),
    .B2(\datamem.data_ram[17][8] ),
    .C1(_06900_),
    .X(_06901_));
 sky130_fd_sc_hd__o22a_1 _19606_ (.A1(\datamem.data_ram[26][8] ),
    .A2(_06802_),
    .B1(_06669_),
    .B2(\datamem.data_ram[31][8] ),
    .X(_06902_));
 sky130_fd_sc_hd__o221a_1 _19607_ (.A1(\datamem.data_ram[29][8] ),
    .A2(_06823_),
    .B1(_06807_),
    .B2(\datamem.data_ram[24][8] ),
    .C1(_06902_),
    .X(_06903_));
 sky130_fd_sc_hd__o22a_1 _19608_ (.A1(\datamem.data_ram[30][8] ),
    .A2(_06717_),
    .B1(_06685_),
    .B2(\datamem.data_ram[28][8] ),
    .X(_06904_));
 sky130_fd_sc_hd__o221a_1 _19609_ (.A1(\datamem.data_ram[27][8] ),
    .A2(_06828_),
    .B1(_06789_),
    .B2(\datamem.data_ram[25][8] ),
    .C1(_06904_),
    .X(_06905_));
 sky130_fd_sc_hd__and3_1 _19610_ (.A(_06810_),
    .B(_06903_),
    .C(_06905_),
    .X(_06906_));
 sky130_fd_sc_hd__a31o_1 _19611_ (.A1(_06680_),
    .A2(_06899_),
    .A3(_06901_),
    .B1(_06906_),
    .X(_06907_));
 sky130_fd_sc_hd__a32o_1 _19612_ (.A1(_06712_),
    .A2(_06886_),
    .A3(_06897_),
    .B1(_06797_),
    .B2(_06907_),
    .X(_06908_));
 sky130_fd_sc_hd__a21oi_4 _19613_ (.A1(_06596_),
    .A2(_06875_),
    .B1(_06908_),
    .Y(_06909_));
 sky130_fd_sc_hd__mux2_1 _19614_ (.A0(_06862_),
    .A1(_06909_),
    .S(_06586_),
    .X(_06910_));
 sky130_fd_sc_hd__nor2_2 _19615_ (.A(_06591_),
    .B(_05386_),
    .Y(_06911_));
 sky130_fd_sc_hd__nand2_1 _19616_ (.A(_05391_),
    .B(_06911_),
    .Y(_06912_));
 sky130_fd_sc_hd__mux2_1 _19617_ (.A0(_06799_),
    .A1(_06910_),
    .S(_06912_),
    .X(_06913_));
 sky130_fd_sc_hd__or2_1 _19618_ (.A(_06586_),
    .B(_06580_),
    .X(_06914_));
 sky130_fd_sc_hd__buf_2 _19619_ (.A(_06914_),
    .X(_06915_));
 sky130_fd_sc_hd__buf_4 _19620_ (.A(_06753_),
    .X(_06916_));
 sky130_fd_sc_hd__nand2_8 _19621_ (.A(_05371_),
    .B(_06641_),
    .Y(_06917_));
 sky130_fd_sc_hd__nor2_1 _19622_ (.A(_06605_),
    .B(_06917_),
    .Y(_06918_));
 sky130_fd_sc_hd__clkbuf_8 _19623_ (.A(_06918_),
    .X(_06919_));
 sky130_fd_sc_hd__buf_4 _19624_ (.A(_06919_),
    .X(_06920_));
 sky130_fd_sc_hd__buf_4 _19625_ (.A(_06920_),
    .X(_06921_));
 sky130_fd_sc_hd__nand2_8 _19626_ (.A(\rvcpu.dp.plem.ALUResultM[4] ),
    .B(_06640_),
    .Y(_06922_));
 sky130_fd_sc_hd__nor2_1 _19627_ (.A(_06605_),
    .B(_06922_),
    .Y(_06923_));
 sky130_fd_sc_hd__buf_4 _19628_ (.A(_06923_),
    .X(_06924_));
 sky130_fd_sc_hd__buf_4 _19629_ (.A(_06924_),
    .X(_06925_));
 sky130_fd_sc_hd__buf_4 _19630_ (.A(_06925_),
    .X(_06926_));
 sky130_fd_sc_hd__clkbuf_4 _19631_ (.A(_06926_),
    .X(_06927_));
 sky130_fd_sc_hd__nand2_4 _19632_ (.A(_06622_),
    .B(_06640_),
    .Y(_06928_));
 sky130_fd_sc_hd__nor2_1 _19633_ (.A(_06666_),
    .B(_06928_),
    .Y(_06929_));
 sky130_fd_sc_hd__clkbuf_8 _19634_ (.A(_06929_),
    .X(_06930_));
 sky130_fd_sc_hd__clkbuf_8 _19635_ (.A(_06930_),
    .X(_06931_));
 sky130_fd_sc_hd__buf_4 _19636_ (.A(_06931_),
    .X(_06932_));
 sky130_fd_sc_hd__buf_6 _19637_ (.A(_06651_),
    .X(_06933_));
 sky130_fd_sc_hd__nand2_8 _19638_ (.A(_06606_),
    .B(_06614_),
    .Y(_06934_));
 sky130_fd_sc_hd__nor2_8 _19639_ (.A(_06933_),
    .B(_06934_),
    .Y(_06935_));
 sky130_fd_sc_hd__buf_4 _19640_ (.A(_06935_),
    .X(_06936_));
 sky130_fd_sc_hd__buf_4 _19641_ (.A(_06936_),
    .X(_06937_));
 sky130_fd_sc_hd__a22o_1 _19642_ (.A1(\datamem.data_ram[34][0] ),
    .A2(_06932_),
    .B1(_06937_),
    .B2(\datamem.data_ram[32][0] ),
    .X(_06938_));
 sky130_fd_sc_hd__a221o_1 _19643_ (.A1(\datamem.data_ram[37][0] ),
    .A2(_06921_),
    .B1(_06927_),
    .B2(\datamem.data_ram[39][0] ),
    .C1(_06938_),
    .X(_06939_));
 sky130_fd_sc_hd__buf_6 _19644_ (.A(_06928_),
    .X(_06940_));
 sky130_fd_sc_hd__nor2_8 _19645_ (.A(_06605_),
    .B(_06940_),
    .Y(_06941_));
 sky130_fd_sc_hd__buf_4 _19646_ (.A(_06941_),
    .X(_06942_));
 sky130_fd_sc_hd__buf_4 _19647_ (.A(_06942_),
    .X(_06943_));
 sky130_fd_sc_hd__buf_6 _19648_ (.A(_06639_),
    .X(_06944_));
 sky130_fd_sc_hd__nor2_2 _19649_ (.A(_06944_),
    .B(_06934_),
    .Y(_06945_));
 sky130_fd_sc_hd__buf_4 _19650_ (.A(_06945_),
    .X(_06946_));
 sky130_fd_sc_hd__clkbuf_8 _19651_ (.A(_06946_),
    .X(_06947_));
 sky130_fd_sc_hd__buf_4 _19652_ (.A(_06947_),
    .X(_06948_));
 sky130_fd_sc_hd__clkbuf_8 _19653_ (.A(_06948_),
    .X(_06949_));
 sky130_fd_sc_hd__nor2_8 _19654_ (.A(\rvcpu.dp.plem.ALUResultM[2] ),
    .B(_06922_),
    .Y(_06950_));
 sky130_fd_sc_hd__buf_4 _19655_ (.A(_06950_),
    .X(_06951_));
 sky130_fd_sc_hd__buf_4 _19656_ (.A(_06951_),
    .X(_06952_));
 sky130_fd_sc_hd__nor2_8 _19657_ (.A(_06666_),
    .B(_06917_),
    .Y(_06953_));
 sky130_fd_sc_hd__buf_4 _19658_ (.A(_06953_),
    .X(_06954_));
 sky130_fd_sc_hd__buf_4 _19659_ (.A(_06954_),
    .X(_06955_));
 sky130_fd_sc_hd__a22o_1 _19660_ (.A1(\datamem.data_ram[38][0] ),
    .A2(_06952_),
    .B1(_06955_),
    .B2(\datamem.data_ram[36][0] ),
    .X(_06956_));
 sky130_fd_sc_hd__a221o_1 _19661_ (.A1(\datamem.data_ram[35][0] ),
    .A2(_06943_),
    .B1(_06949_),
    .B2(\datamem.data_ram[33][0] ),
    .C1(_06956_),
    .X(_06957_));
 sky130_fd_sc_hd__buf_4 _19662_ (.A(_06947_),
    .X(_06958_));
 sky130_fd_sc_hd__a22o_1 _19663_ (.A1(\datamem.data_ram[42][0] ),
    .A2(_06931_),
    .B1(_06925_),
    .B2(\datamem.data_ram[47][0] ),
    .X(_06959_));
 sky130_fd_sc_hd__a221o_1 _19664_ (.A1(\datamem.data_ram[46][0] ),
    .A2(_06952_),
    .B1(_06958_),
    .B2(\datamem.data_ram[41][0] ),
    .C1(_06959_),
    .X(_06960_));
 sky130_fd_sc_hd__buf_4 _19665_ (.A(_06941_),
    .X(_06961_));
 sky130_fd_sc_hd__a22o_1 _19666_ (.A1(\datamem.data_ram[40][0] ),
    .A2(_06936_),
    .B1(_06954_),
    .B2(\datamem.data_ram[44][0] ),
    .X(_06962_));
 sky130_fd_sc_hd__a221o_1 _19667_ (.A1(\datamem.data_ram[45][0] ),
    .A2(_06920_),
    .B1(_06961_),
    .B2(\datamem.data_ram[43][0] ),
    .C1(_06962_),
    .X(_06963_));
 sky130_fd_sc_hd__or3_1 _19668_ (.A(_06680_),
    .B(_06960_),
    .C(_06963_),
    .X(_06964_));
 sky130_fd_sc_hd__o31a_1 _19669_ (.A1(_06603_),
    .A2(_06939_),
    .A3(_06957_),
    .B1(_06964_),
    .X(_06965_));
 sky130_fd_sc_hd__buf_4 _19670_ (.A(_06943_),
    .X(_06966_));
 sky130_fd_sc_hd__buf_6 _19671_ (.A(_06810_),
    .X(_06967_));
 sky130_fd_sc_hd__a221o_1 _19672_ (.A1(\datamem.data_ram[51][0] ),
    .A2(_06966_),
    .B1(_06927_),
    .B2(\datamem.data_ram[55][0] ),
    .C1(_06967_),
    .X(_06968_));
 sky130_fd_sc_hd__buf_4 _19673_ (.A(_06920_),
    .X(_06969_));
 sky130_fd_sc_hd__clkbuf_4 _19674_ (.A(_06969_),
    .X(_06970_));
 sky130_fd_sc_hd__a22o_1 _19675_ (.A1(\datamem.data_ram[54][0] ),
    .A2(_06951_),
    .B1(_06958_),
    .B2(\datamem.data_ram[49][0] ),
    .X(_06971_));
 sky130_fd_sc_hd__a21o_1 _19676_ (.A1(\datamem.data_ram[50][0] ),
    .A2(_06932_),
    .B1(_06971_),
    .X(_06972_));
 sky130_fd_sc_hd__buf_6 _19677_ (.A(_06936_),
    .X(_06973_));
 sky130_fd_sc_hd__a22o_1 _19678_ (.A1(\datamem.data_ram[48][0] ),
    .A2(_06973_),
    .B1(_06955_),
    .B2(\datamem.data_ram[52][0] ),
    .X(_06974_));
 sky130_fd_sc_hd__a211o_1 _19679_ (.A1(\datamem.data_ram[53][0] ),
    .A2(_06970_),
    .B1(_06972_),
    .C1(_06974_),
    .X(_06975_));
 sky130_fd_sc_hd__buf_4 _19680_ (.A(_06954_),
    .X(_06976_));
 sky130_fd_sc_hd__buf_4 _19681_ (.A(_06976_),
    .X(_06977_));
 sky130_fd_sc_hd__buf_4 _19682_ (.A(_06951_),
    .X(_06978_));
 sky130_fd_sc_hd__a22o_1 _19683_ (.A1(\datamem.data_ram[62][0] ),
    .A2(_06978_),
    .B1(_06926_),
    .B2(\datamem.data_ram[63][0] ),
    .X(_06979_));
 sky130_fd_sc_hd__a22o_1 _19684_ (.A1(\datamem.data_ram[56][0] ),
    .A2(_06936_),
    .B1(_06947_),
    .B2(\datamem.data_ram[57][0] ),
    .X(_06980_));
 sky130_fd_sc_hd__a221o_1 _19685_ (.A1(\datamem.data_ram[58][0] ),
    .A2(_06931_),
    .B1(_06942_),
    .B2(\datamem.data_ram[59][0] ),
    .C1(_06769_),
    .X(_06981_));
 sky130_fd_sc_hd__a211o_1 _19686_ (.A1(\datamem.data_ram[61][0] ),
    .A2(_06969_),
    .B1(_06980_),
    .C1(_06981_),
    .X(_06982_));
 sky130_fd_sc_hd__a211o_1 _19687_ (.A1(\datamem.data_ram[60][0] ),
    .A2(_06977_),
    .B1(_06979_),
    .C1(_06982_),
    .X(_06983_));
 sky130_fd_sc_hd__o211a_1 _19688_ (.A1(_06968_),
    .A2(_06975_),
    .B1(_06983_),
    .C1(_06716_),
    .X(_06984_));
 sky130_fd_sc_hd__clkbuf_8 _19689_ (.A(_06860_),
    .X(_06985_));
 sky130_fd_sc_hd__a211o_1 _19690_ (.A1(_06916_),
    .A2(_06965_),
    .B1(_06984_),
    .C1(_06985_),
    .X(_06986_));
 sky130_fd_sc_hd__inv_2 _19691_ (.A(_06582_),
    .Y(_06987_));
 sky130_fd_sc_hd__o22a_2 _19692_ (.A1(_06586_),
    .A2(_06987_),
    .B1(_06583_),
    .B2(_06588_),
    .X(_06988_));
 sky130_fd_sc_hd__buf_4 _19693_ (.A(_06931_),
    .X(_06989_));
 sky130_fd_sc_hd__clkbuf_8 _19694_ (.A(_06937_),
    .X(_06990_));
 sky130_fd_sc_hd__a22o_1 _19695_ (.A1(\datamem.data_ram[12][0] ),
    .A2(_06955_),
    .B1(_06958_),
    .B2(\datamem.data_ram[9][0] ),
    .X(_06991_));
 sky130_fd_sc_hd__a221o_1 _19696_ (.A1(\datamem.data_ram[10][0] ),
    .A2(_06989_),
    .B1(_06990_),
    .B2(\datamem.data_ram[8][0] ),
    .C1(_06991_),
    .X(_06992_));
 sky130_fd_sc_hd__buf_4 _19697_ (.A(_06925_),
    .X(_06993_));
 sky130_fd_sc_hd__a22o_1 _19698_ (.A1(\datamem.data_ram[14][0] ),
    .A2(_06952_),
    .B1(_06961_),
    .B2(\datamem.data_ram[11][0] ),
    .X(_06994_));
 sky130_fd_sc_hd__a221o_1 _19699_ (.A1(\datamem.data_ram[13][0] ),
    .A2(_06921_),
    .B1(_06993_),
    .B2(\datamem.data_ram[15][0] ),
    .C1(_06994_),
    .X(_06995_));
 sky130_fd_sc_hd__or3_1 _19700_ (.A(_06777_),
    .B(_06992_),
    .C(_06995_),
    .X(_06996_));
 sky130_fd_sc_hd__clkbuf_8 _19701_ (.A(_06949_),
    .X(_06997_));
 sky130_fd_sc_hd__a22o_1 _19702_ (.A1(\datamem.data_ram[7][0] ),
    .A2(_06926_),
    .B1(_06955_),
    .B2(\datamem.data_ram[4][0] ),
    .X(_06998_));
 sky130_fd_sc_hd__a211o_1 _19703_ (.A1(\datamem.data_ram[5][0] ),
    .A2(_06970_),
    .B1(_06967_),
    .C1(_06998_),
    .X(_06999_));
 sky130_fd_sc_hd__clkbuf_8 _19704_ (.A(_06932_),
    .X(_07000_));
 sky130_fd_sc_hd__a22o_1 _19705_ (.A1(\datamem.data_ram[6][0] ),
    .A2(_06952_),
    .B1(_06973_),
    .B2(\datamem.data_ram[0][0] ),
    .X(_07001_));
 sky130_fd_sc_hd__a221o_1 _19706_ (.A1(\datamem.data_ram[2][0] ),
    .A2(_07000_),
    .B1(_06966_),
    .B2(\datamem.data_ram[3][0] ),
    .C1(_07001_),
    .X(_07002_));
 sky130_fd_sc_hd__a211o_1 _19707_ (.A1(\datamem.data_ram[1][0] ),
    .A2(_06997_),
    .B1(_06999_),
    .C1(_07002_),
    .X(_07003_));
 sky130_fd_sc_hd__a22o_1 _19708_ (.A1(\datamem.data_ram[23][0] ),
    .A2(_06926_),
    .B1(_06948_),
    .B2(\datamem.data_ram[17][0] ),
    .X(_07004_));
 sky130_fd_sc_hd__a22o_1 _19709_ (.A1(\datamem.data_ram[21][0] ),
    .A2(_06920_),
    .B1(_06954_),
    .B2(\datamem.data_ram[20][0] ),
    .X(_07005_));
 sky130_fd_sc_hd__a221o_1 _19710_ (.A1(\datamem.data_ram[22][0] ),
    .A2(_06951_),
    .B1(_06936_),
    .B2(\datamem.data_ram[16][0] ),
    .C1(_06741_),
    .X(_07006_));
 sky130_fd_sc_hd__a211o_1 _19711_ (.A1(\datamem.data_ram[18][0] ),
    .A2(_06989_),
    .B1(_07005_),
    .C1(_07006_),
    .X(_07007_));
 sky130_fd_sc_hd__a211o_1 _19712_ (.A1(\datamem.data_ram[19][0] ),
    .A2(_06966_),
    .B1(_07004_),
    .C1(_07007_),
    .X(_07008_));
 sky130_fd_sc_hd__a22o_1 _19713_ (.A1(\datamem.data_ram[30][0] ),
    .A2(_06978_),
    .B1(_06976_),
    .B2(\datamem.data_ram[28][0] ),
    .X(_07009_));
 sky130_fd_sc_hd__a22o_1 _19714_ (.A1(\datamem.data_ram[31][0] ),
    .A2(_06925_),
    .B1(_06958_),
    .B2(\datamem.data_ram[25][0] ),
    .X(_07010_));
 sky130_fd_sc_hd__a221o_1 _19715_ (.A1(\datamem.data_ram[24][0] ),
    .A2(_06936_),
    .B1(_06942_),
    .B2(\datamem.data_ram[27][0] ),
    .C1(_06769_),
    .X(_07011_));
 sky130_fd_sc_hd__a211o_1 _19716_ (.A1(\datamem.data_ram[26][0] ),
    .A2(_06989_),
    .B1(_07010_),
    .C1(_07011_),
    .X(_07012_));
 sky130_fd_sc_hd__a211o_1 _19717_ (.A1(\datamem.data_ram[29][0] ),
    .A2(_06970_),
    .B1(_07009_),
    .C1(_07012_),
    .X(_07013_));
 sky130_fd_sc_hd__a31o_1 _19718_ (.A1(_06716_),
    .A2(_07008_),
    .A3(_07013_),
    .B1(_06713_),
    .X(_07014_));
 sky130_fd_sc_hd__a31o_1 _19719_ (.A1(_06916_),
    .A2(_06996_),
    .A3(_07003_),
    .B1(_07014_),
    .X(_07015_));
 sky130_fd_sc_hd__and3_1 _19720_ (.A(_06986_),
    .B(_06988_),
    .C(_07015_),
    .X(_07016_));
 sky130_fd_sc_hd__o21ba_1 _19721_ (.A1(_06799_),
    .A2(_06915_),
    .B1_N(_07016_),
    .X(_07017_));
 sky130_fd_sc_hd__o21ai_1 _19722_ (.A1(_06590_),
    .A2(_06913_),
    .B1(_07017_),
    .Y(_04415_));
 sky130_fd_sc_hd__or2_1 _19723_ (.A(\datamem.data_ram[9][25] ),
    .B(_06659_),
    .X(_07018_));
 sky130_fd_sc_hd__buf_6 _19724_ (.A(_06865_),
    .X(_07019_));
 sky130_fd_sc_hd__buf_6 _19725_ (.A(_06784_),
    .X(_07020_));
 sky130_fd_sc_hd__buf_6 _19726_ (.A(_07020_),
    .X(_07021_));
 sky130_fd_sc_hd__o22a_1 _19727_ (.A1(\datamem.data_ram[13][25] ),
    .A2(_07019_),
    .B1(_07021_),
    .B2(\datamem.data_ram[15][25] ),
    .X(_07022_));
 sky130_fd_sc_hd__buf_8 _19728_ (.A(_06754_),
    .X(_07023_));
 sky130_fd_sc_hd__buf_6 _19729_ (.A(_06766_),
    .X(_07024_));
 sky130_fd_sc_hd__o22a_1 _19730_ (.A1(\datamem.data_ram[11][25] ),
    .A2(_06738_),
    .B1(_07024_),
    .B2(\datamem.data_ram[12][25] ),
    .X(_07025_));
 sky130_fd_sc_hd__o221a_1 _19731_ (.A1(\datamem.data_ram[14][25] ),
    .A2(_06683_),
    .B1(_07023_),
    .B2(\datamem.data_ram[10][25] ),
    .C1(_07025_),
    .X(_07026_));
 sky130_fd_sc_hd__o211a_1 _19732_ (.A1(\datamem.data_ram[8][25] ),
    .A2(_06649_),
    .B1(_07026_),
    .C1(_06603_),
    .X(_07027_));
 sky130_fd_sc_hd__buf_8 _19733_ (.A(_06683_),
    .X(_07028_));
 sky130_fd_sc_hd__o22a_1 _19734_ (.A1(\datamem.data_ram[0][25] ),
    .A2(_06698_),
    .B1(_06688_),
    .B2(\datamem.data_ram[4][25] ),
    .X(_07029_));
 sky130_fd_sc_hd__o22a_1 _19735_ (.A1(\datamem.data_ram[5][25] ),
    .A2(_06703_),
    .B1(_06707_),
    .B2(\datamem.data_ram[7][25] ),
    .X(_07030_));
 sky130_fd_sc_hd__buf_8 _19736_ (.A(_06769_),
    .X(_07031_));
 sky130_fd_sc_hd__o221a_1 _19737_ (.A1(\datamem.data_ram[3][25] ),
    .A2(_06738_),
    .B1(_06700_),
    .B2(\datamem.data_ram[1][25] ),
    .C1(_07031_),
    .X(_07032_));
 sky130_fd_sc_hd__o211a_1 _19738_ (.A1(\datamem.data_ram[2][25] ),
    .A2(_07023_),
    .B1(_07030_),
    .C1(_07032_),
    .X(_07033_));
 sky130_fd_sc_hd__o211a_1 _19739_ (.A1(\datamem.data_ram[6][25] ),
    .A2(_07028_),
    .B1(_07029_),
    .C1(_07033_),
    .X(_07034_));
 sky130_fd_sc_hd__a31o_1 _19740_ (.A1(_07018_),
    .A2(_07022_),
    .A3(_07027_),
    .B1(_07034_),
    .X(_07035_));
 sky130_fd_sc_hd__o22a_1 _19741_ (.A1(\datamem.data_ram[38][25] ),
    .A2(_06719_),
    .B1(_06687_),
    .B2(\datamem.data_ram[36][25] ),
    .X(_07036_));
 sky130_fd_sc_hd__buf_6 _19742_ (.A(_06823_),
    .X(_07037_));
 sky130_fd_sc_hd__o22a_1 _19743_ (.A1(\datamem.data_ram[39][25] ),
    .A2(_06726_),
    .B1(_06656_),
    .B2(\datamem.data_ram[33][25] ),
    .X(_07038_));
 sky130_fd_sc_hd__o221a_1 _19744_ (.A1(\datamem.data_ram[32][25] ),
    .A2(_06821_),
    .B1(_06828_),
    .B2(\datamem.data_ram[35][25] ),
    .C1(_06733_),
    .X(_07039_));
 sky130_fd_sc_hd__o211a_1 _19745_ (.A1(\datamem.data_ram[37][25] ),
    .A2(_07037_),
    .B1(_07038_),
    .C1(_07039_),
    .X(_07040_));
 sky130_fd_sc_hd__o211a_1 _19746_ (.A1(\datamem.data_ram[34][25] ),
    .A2(_07023_),
    .B1(_07036_),
    .C1(_07040_),
    .X(_07041_));
 sky130_fd_sc_hd__o22a_1 _19747_ (.A1(\datamem.data_ram[46][25] ),
    .A2(_06719_),
    .B1(_06657_),
    .B2(\datamem.data_ram[41][25] ),
    .X(_07042_));
 sky130_fd_sc_hd__o22a_1 _19748_ (.A1(\datamem.data_ram[47][25] ),
    .A2(_06725_),
    .B1(_06765_),
    .B2(\datamem.data_ram[44][25] ),
    .X(_07043_));
 sky130_fd_sc_hd__o221a_1 _19749_ (.A1(\datamem.data_ram[45][25] ),
    .A2(_06723_),
    .B1(_06807_),
    .B2(\datamem.data_ram[40][25] ),
    .C1(_07043_),
    .X(_07044_));
 sky130_fd_sc_hd__o211a_1 _19750_ (.A1(\datamem.data_ram[42][25] ),
    .A2(_06754_),
    .B1(_06810_),
    .C1(_07044_),
    .X(_07045_));
 sky130_fd_sc_hd__o211a_1 _19751_ (.A1(\datamem.data_ram[43][25] ),
    .A2(_06863_),
    .B1(_07042_),
    .C1(_07045_),
    .X(_07046_));
 sky130_fd_sc_hd__or3_1 _19752_ (.A(_06715_),
    .B(_07041_),
    .C(_07046_),
    .X(_07047_));
 sky130_fd_sc_hd__o22a_1 _19753_ (.A1(\datamem.data_ram[61][25] ),
    .A2(_07037_),
    .B1(_06657_),
    .B2(\datamem.data_ram[57][25] ),
    .X(_07048_));
 sky130_fd_sc_hd__o22a_1 _19754_ (.A1(\datamem.data_ram[59][25] ),
    .A2(_06812_),
    .B1(_06765_),
    .B2(\datamem.data_ram[60][25] ),
    .X(_07049_));
 sky130_fd_sc_hd__o221a_1 _19755_ (.A1(\datamem.data_ram[56][25] ),
    .A2(_06807_),
    .B1(_06726_),
    .B2(\datamem.data_ram[63][25] ),
    .C1(_07049_),
    .X(_07050_));
 sky130_fd_sc_hd__o211a_1 _19756_ (.A1(\datamem.data_ram[62][25] ),
    .A2(_06719_),
    .B1(_06810_),
    .C1(_07050_),
    .X(_07051_));
 sky130_fd_sc_hd__o211a_1 _19757_ (.A1(\datamem.data_ram[58][25] ),
    .A2(_07023_),
    .B1(_07048_),
    .C1(_07051_),
    .X(_07052_));
 sky130_fd_sc_hd__o22a_1 _19758_ (.A1(\datamem.data_ram[54][25] ),
    .A2(_06719_),
    .B1(_06671_),
    .B2(\datamem.data_ram[55][25] ),
    .X(_07053_));
 sky130_fd_sc_hd__o22a_1 _19759_ (.A1(\datamem.data_ram[50][25] ),
    .A2(_06803_),
    .B1(_06696_),
    .B2(\datamem.data_ram[48][25] ),
    .X(_07054_));
 sky130_fd_sc_hd__o221a_1 _19760_ (.A1(\datamem.data_ram[53][25] ),
    .A2(_06723_),
    .B1(_06731_),
    .B2(\datamem.data_ram[51][25] ),
    .C1(_06733_),
    .X(_07055_));
 sky130_fd_sc_hd__o211a_1 _19761_ (.A1(\datamem.data_ram[52][25] ),
    .A2(_06687_),
    .B1(_07054_),
    .C1(_07055_),
    .X(_07056_));
 sky130_fd_sc_hd__o211a_1 _19762_ (.A1(\datamem.data_ram[49][25] ),
    .A2(_06658_),
    .B1(_07053_),
    .C1(_07056_),
    .X(_07057_));
 sky130_fd_sc_hd__or3_1 _19763_ (.A(_06752_),
    .B(_07052_),
    .C(_07057_),
    .X(_07058_));
 sky130_fd_sc_hd__o22a_1 _19764_ (.A1(\datamem.data_ram[20][25] ),
    .A2(_07024_),
    .B1(_06700_),
    .B2(\datamem.data_ram[17][25] ),
    .X(_07059_));
 sky130_fd_sc_hd__o221a_1 _19765_ (.A1(\datamem.data_ram[21][25] ),
    .A2(_06865_),
    .B1(_06672_),
    .B2(\datamem.data_ram[23][25] ),
    .C1(_07059_),
    .X(_07060_));
 sky130_fd_sc_hd__o22a_1 _19766_ (.A1(\datamem.data_ram[18][25] ),
    .A2(_06692_),
    .B1(_06779_),
    .B2(\datamem.data_ram[16][25] ),
    .X(_07061_));
 sky130_fd_sc_hd__o221a_1 _19767_ (.A1(\datamem.data_ram[22][25] ),
    .A2(_06683_),
    .B1(_06739_),
    .B2(\datamem.data_ram[19][25] ),
    .C1(_07061_),
    .X(_07062_));
 sky130_fd_sc_hd__o22a_1 _19768_ (.A1(\datamem.data_ram[30][25] ),
    .A2(_06763_),
    .B1(_06691_),
    .B2(\datamem.data_ram[26][25] ),
    .X(_07063_));
 sky130_fd_sc_hd__o221a_1 _19769_ (.A1(\datamem.data_ram[24][25] ),
    .A2(_06697_),
    .B1(_06657_),
    .B2(\datamem.data_ram[25][25] ),
    .C1(_07063_),
    .X(_07064_));
 sky130_fd_sc_hd__o22a_1 _19770_ (.A1(\datamem.data_ram[29][25] ),
    .A2(_06768_),
    .B1(_06760_),
    .B2(\datamem.data_ram[31][25] ),
    .X(_07065_));
 sky130_fd_sc_hd__o221a_1 _19771_ (.A1(\datamem.data_ram[27][25] ),
    .A2(_06829_),
    .B1(_07024_),
    .B2(\datamem.data_ram[28][25] ),
    .C1(_07065_),
    .X(_07066_));
 sky130_fd_sc_hd__and3_1 _19772_ (.A(_06967_),
    .B(_07064_),
    .C(_07066_),
    .X(_07067_));
 sky130_fd_sc_hd__a31o_1 _19773_ (.A1(_06681_),
    .A2(_07060_),
    .A3(_07062_),
    .B1(_07067_),
    .X(_07068_));
 sky130_fd_sc_hd__a32o_1 _19774_ (.A1(_06713_),
    .A2(_07047_),
    .A3(_07058_),
    .B1(_07068_),
    .B2(_06797_),
    .X(_07069_));
 sky130_fd_sc_hd__a21oi_4 _19775_ (.A1(_06596_),
    .A2(_07035_),
    .B1(_07069_),
    .Y(_07070_));
 sky130_fd_sc_hd__clkbuf_8 _19776_ (.A(_06716_),
    .X(_07071_));
 sky130_fd_sc_hd__o22a_1 _19777_ (.A1(\datamem.data_ram[38][9] ),
    .A2(_06683_),
    .B1(_06688_),
    .B2(\datamem.data_ram[36][9] ),
    .X(_07072_));
 sky130_fd_sc_hd__o22a_1 _19778_ (.A1(\datamem.data_ram[39][9] ),
    .A2(_06761_),
    .B1(_06700_),
    .B2(\datamem.data_ram[33][9] ),
    .X(_07073_));
 sky130_fd_sc_hd__o221a_1 _19779_ (.A1(\datamem.data_ram[34][9] ),
    .A2(_06754_),
    .B1(_06738_),
    .B2(\datamem.data_ram[35][9] ),
    .C1(_07031_),
    .X(_07074_));
 sky130_fd_sc_hd__o211a_1 _19780_ (.A1(\datamem.data_ram[37][9] ),
    .A2(_06865_),
    .B1(_07073_),
    .C1(_07074_),
    .X(_07075_));
 sky130_fd_sc_hd__o211a_1 _19781_ (.A1(\datamem.data_ram[32][9] ),
    .A2(_06649_),
    .B1(_07072_),
    .C1(_07075_),
    .X(_07076_));
 sky130_fd_sc_hd__clkbuf_8 _19782_ (.A(_06863_),
    .X(_07077_));
 sky130_fd_sc_hd__o22a_1 _19783_ (.A1(\datamem.data_ram[44][9] ),
    .A2(_06688_),
    .B1(_06701_),
    .B2(\datamem.data_ram[41][9] ),
    .X(_07078_));
 sky130_fd_sc_hd__o22a_1 _19784_ (.A1(\datamem.data_ram[46][9] ),
    .A2(_06763_),
    .B1(_06611_),
    .B2(\datamem.data_ram[42][9] ),
    .X(_07079_));
 sky130_fd_sc_hd__o221a_1 _19785_ (.A1(\datamem.data_ram[45][9] ),
    .A2(_06703_),
    .B1(_06779_),
    .B2(\datamem.data_ram[40][9] ),
    .C1(_07079_),
    .X(_07080_));
 sky130_fd_sc_hd__clkbuf_8 _19786_ (.A(_06602_),
    .X(_07081_));
 sky130_fd_sc_hd__o211a_1 _19787_ (.A1(\datamem.data_ram[47][9] ),
    .A2(_06672_),
    .B1(_07080_),
    .C1(_07081_),
    .X(_07082_));
 sky130_fd_sc_hd__o211a_1 _19788_ (.A1(\datamem.data_ram[43][9] ),
    .A2(_07077_),
    .B1(_07078_),
    .C1(_07082_),
    .X(_07083_));
 sky130_fd_sc_hd__o22a_1 _19789_ (.A1(\datamem.data_ram[55][9] ),
    .A2(_06707_),
    .B1(_06783_),
    .B2(\datamem.data_ram[49][9] ),
    .X(_07084_));
 sky130_fd_sc_hd__buf_6 _19790_ (.A(_06743_),
    .X(_07085_));
 sky130_fd_sc_hd__o22a_1 _19791_ (.A1(\datamem.data_ram[54][9] ),
    .A2(_07085_),
    .B1(_06633_),
    .B2(\datamem.data_ram[51][9] ),
    .X(_07086_));
 sky130_fd_sc_hd__o221a_1 _19792_ (.A1(\datamem.data_ram[48][9] ),
    .A2(_06778_),
    .B1(_06766_),
    .B2(\datamem.data_ram[52][9] ),
    .C1(_07086_),
    .X(_07087_));
 sky130_fd_sc_hd__o211a_1 _19793_ (.A1(\datamem.data_ram[53][9] ),
    .A2(_06703_),
    .B1(_07031_),
    .C1(_07087_),
    .X(_07088_));
 sky130_fd_sc_hd__o211a_1 _19794_ (.A1(\datamem.data_ram[50][9] ),
    .A2(_07023_),
    .B1(_07084_),
    .C1(_07088_),
    .X(_07089_));
 sky130_fd_sc_hd__o22a_1 _19795_ (.A1(\datamem.data_ram[62][9] ),
    .A2(_06629_),
    .B1(_06620_),
    .B2(\datamem.data_ram[60][9] ),
    .X(_07090_));
 sky130_fd_sc_hd__o22a_1 _19796_ (.A1(\datamem.data_ram[61][9] ),
    .A2(_06663_),
    .B1(_06706_),
    .B2(\datamem.data_ram[63][9] ),
    .X(_07091_));
 sky130_fd_sc_hd__o221a_1 _19797_ (.A1(\datamem.data_ram[58][9] ),
    .A2(_06611_),
    .B1(_06647_),
    .B2(\datamem.data_ram[56][9] ),
    .C1(_06601_),
    .X(_07092_));
 sky130_fd_sc_hd__o211a_1 _19798_ (.A1(\datamem.data_ram[57][9] ),
    .A2(_06783_),
    .B1(_07091_),
    .C1(_07092_),
    .X(_07093_));
 sky130_fd_sc_hd__o211a_1 _19799_ (.A1(\datamem.data_ram[59][9] ),
    .A2(_06636_),
    .B1(_07090_),
    .C1(_07093_),
    .X(_07094_));
 sky130_fd_sc_hd__o31a_1 _19800_ (.A1(_06753_),
    .A2(_07089_),
    .A3(_07094_),
    .B1(_06713_),
    .X(_07095_));
 sky130_fd_sc_hd__o31a_1 _19801_ (.A1(_07071_),
    .A2(_07076_),
    .A3(_07083_),
    .B1(_07095_),
    .X(_07096_));
 sky130_fd_sc_hd__o22a_1 _19802_ (.A1(\datamem.data_ram[15][9] ),
    .A2(_06761_),
    .B1(_06783_),
    .B2(\datamem.data_ram[9][9] ),
    .X(_07097_));
 sky130_fd_sc_hd__o221a_1 _19803_ (.A1(\datamem.data_ram[13][9] ),
    .A2(_06865_),
    .B1(_06688_),
    .B2(\datamem.data_ram[12][9] ),
    .C1(_07097_),
    .X(_07098_));
 sky130_fd_sc_hd__o22a_1 _19804_ (.A1(\datamem.data_ram[14][9] ),
    .A2(_06764_),
    .B1(_06692_),
    .B2(\datamem.data_ram[10][9] ),
    .X(_07099_));
 sky130_fd_sc_hd__o221a_1 _19805_ (.A1(\datamem.data_ram[8][9] ),
    .A2(_06698_),
    .B1(_06739_),
    .B2(\datamem.data_ram[11][9] ),
    .C1(_07099_),
    .X(_07100_));
 sky130_fd_sc_hd__o22a_1 _19806_ (.A1(\datamem.data_ram[2][9] ),
    .A2(_06691_),
    .B1(_06760_),
    .B2(\datamem.data_ram[7][9] ),
    .X(_07101_));
 sky130_fd_sc_hd__o221a_1 _19807_ (.A1(\datamem.data_ram[6][9] ),
    .A2(_06719_),
    .B1(_06697_),
    .B2(\datamem.data_ram[0][9] ),
    .C1(_07101_),
    .X(_07102_));
 sky130_fd_sc_hd__o22a_1 _19808_ (.A1(\datamem.data_ram[4][9] ),
    .A2(_06766_),
    .B1(_06699_),
    .B2(\datamem.data_ram[1][9] ),
    .X(_07103_));
 sky130_fd_sc_hd__o221a_1 _19809_ (.A1(\datamem.data_ram[5][9] ),
    .A2(_06724_),
    .B1(_06738_),
    .B2(\datamem.data_ram[3][9] ),
    .C1(_07103_),
    .X(_07104_));
 sky130_fd_sc_hd__and3_1 _19810_ (.A(_06680_),
    .B(_07102_),
    .C(_07104_),
    .X(_07105_));
 sky130_fd_sc_hd__a31o_1 _19811_ (.A1(_06603_),
    .A2(_07098_),
    .A3(_07100_),
    .B1(_07105_),
    .X(_07106_));
 sky130_fd_sc_hd__or2_1 _19812_ (.A(\datamem.data_ram[18][9] ),
    .B(_06613_),
    .X(_07107_));
 sky130_fd_sc_hd__o22a_1 _19813_ (.A1(\datamem.data_ram[22][9] ),
    .A2(_06630_),
    .B1(_06672_),
    .B2(\datamem.data_ram[23][9] ),
    .X(_07108_));
 sky130_fd_sc_hd__o22a_1 _19814_ (.A1(\datamem.data_ram[21][9] ),
    .A2(_06702_),
    .B1(_06619_),
    .B2(\datamem.data_ram[20][9] ),
    .X(_07109_));
 sky130_fd_sc_hd__o221a_1 _19815_ (.A1(\datamem.data_ram[16][9] ),
    .A2(_06697_),
    .B1(_06700_),
    .B2(\datamem.data_ram[17][9] ),
    .C1(_07109_),
    .X(_07110_));
 sky130_fd_sc_hd__o211a_1 _19816_ (.A1(\datamem.data_ram[19][9] ),
    .A2(_06636_),
    .B1(_07110_),
    .C1(_06777_),
    .X(_07111_));
 sky130_fd_sc_hd__o22a_1 _19817_ (.A1(\datamem.data_ram[30][9] ),
    .A2(_06629_),
    .B1(_06620_),
    .B2(\datamem.data_ram[28][9] ),
    .X(_07112_));
 sky130_fd_sc_hd__o22a_1 _19818_ (.A1(\datamem.data_ram[24][9] ),
    .A2(_06647_),
    .B1(_06782_),
    .B2(\datamem.data_ram[25][9] ),
    .X(_07113_));
 sky130_fd_sc_hd__o221a_1 _19819_ (.A1(\datamem.data_ram[26][9] ),
    .A2(_06611_),
    .B1(_06634_),
    .B2(\datamem.data_ram[27][9] ),
    .C1(_06601_),
    .X(_07114_));
 sky130_fd_sc_hd__o211a_1 _19820_ (.A1(\datamem.data_ram[29][9] ),
    .A2(_06703_),
    .B1(_07113_),
    .C1(_07114_),
    .X(_07115_));
 sky130_fd_sc_hd__o211a_1 _19821_ (.A1(\datamem.data_ram[31][9] ),
    .A2(_06672_),
    .B1(_07112_),
    .C1(_07115_),
    .X(_07116_));
 sky130_fd_sc_hd__a31o_1 _19822_ (.A1(_07107_),
    .A2(_07108_),
    .A3(_07111_),
    .B1(_07116_),
    .X(_07117_));
 sky130_fd_sc_hd__a22o_1 _19823_ (.A1(_06596_),
    .A2(_07106_),
    .B1(_07117_),
    .B2(_06797_),
    .X(_07118_));
 sky130_fd_sc_hd__nor2_2 _19824_ (.A(_07096_),
    .B(_07118_),
    .Y(_07119_));
 sky130_fd_sc_hd__or2_1 _19825_ (.A(\rvcpu.dp.plem.ALUResultM[1] ),
    .B(_06588_),
    .X(_07120_));
 sky130_fd_sc_hd__o32a_1 _19826_ (.A1(_05391_),
    .A2(_06586_),
    .A3(_07070_),
    .B1(_07119_),
    .B2(_07120_),
    .X(_07121_));
 sky130_fd_sc_hd__clkbuf_8 _19827_ (.A(_06990_),
    .X(_07122_));
 sky130_fd_sc_hd__buf_4 _19828_ (.A(_06976_),
    .X(_07123_));
 sky130_fd_sc_hd__a22o_1 _19829_ (.A1(\datamem.data_ram[32][1] ),
    .A2(_07122_),
    .B1(_07123_),
    .B2(\datamem.data_ram[36][1] ),
    .X(_07124_));
 sky130_fd_sc_hd__buf_8 _19830_ (.A(_06993_),
    .X(_07125_));
 sky130_fd_sc_hd__a22o_1 _19831_ (.A1(\datamem.data_ram[34][1] ),
    .A2(_07000_),
    .B1(_06970_),
    .B2(\datamem.data_ram[37][1] ),
    .X(_07126_));
 sky130_fd_sc_hd__buf_4 _19832_ (.A(_06952_),
    .X(_07127_));
 sky130_fd_sc_hd__a221o_1 _19833_ (.A1(\datamem.data_ram[38][1] ),
    .A2(_07127_),
    .B1(_06966_),
    .B2(\datamem.data_ram[35][1] ),
    .C1(_06967_),
    .X(_07128_));
 sky130_fd_sc_hd__a211o_1 _19834_ (.A1(\datamem.data_ram[39][1] ),
    .A2(_07125_),
    .B1(_07126_),
    .C1(_07128_),
    .X(_07129_));
 sky130_fd_sc_hd__a211o_1 _19835_ (.A1(\datamem.data_ram[33][1] ),
    .A2(_06997_),
    .B1(_07124_),
    .C1(_07129_),
    .X(_07130_));
 sky130_fd_sc_hd__buf_4 _19836_ (.A(_06777_),
    .X(_07131_));
 sky130_fd_sc_hd__buf_6 _19837_ (.A(_06921_),
    .X(_07132_));
 sky130_fd_sc_hd__clkbuf_8 _19838_ (.A(_06948_),
    .X(_07133_));
 sky130_fd_sc_hd__a22o_1 _19839_ (.A1(\datamem.data_ram[47][1] ),
    .A2(_06993_),
    .B1(_06976_),
    .B2(\datamem.data_ram[44][1] ),
    .X(_07134_));
 sky130_fd_sc_hd__a221o_1 _19840_ (.A1(\datamem.data_ram[45][1] ),
    .A2(_07132_),
    .B1(_07133_),
    .B2(\datamem.data_ram[41][1] ),
    .C1(_07134_),
    .X(_07135_));
 sky130_fd_sc_hd__clkbuf_8 _19841_ (.A(_06989_),
    .X(_07136_));
 sky130_fd_sc_hd__clkbuf_8 _19842_ (.A(_06943_),
    .X(_07137_));
 sky130_fd_sc_hd__buf_4 _19843_ (.A(_06973_),
    .X(_07138_));
 sky130_fd_sc_hd__a22o_1 _19844_ (.A1(\datamem.data_ram[46][1] ),
    .A2(_06978_),
    .B1(_07138_),
    .B2(\datamem.data_ram[40][1] ),
    .X(_07139_));
 sky130_fd_sc_hd__a221o_1 _19845_ (.A1(\datamem.data_ram[42][1] ),
    .A2(_07136_),
    .B1(_07137_),
    .B2(\datamem.data_ram[43][1] ),
    .C1(_07139_),
    .X(_07140_));
 sky130_fd_sc_hd__or3_1 _19846_ (.A(_07131_),
    .B(_07135_),
    .C(_07140_),
    .X(_07141_));
 sky130_fd_sc_hd__a22o_1 _19847_ (.A1(\datamem.data_ram[54][1] ),
    .A2(_06952_),
    .B1(_06969_),
    .B2(\datamem.data_ram[53][1] ),
    .X(_07142_));
 sky130_fd_sc_hd__a221o_1 _19848_ (.A1(\datamem.data_ram[48][1] ),
    .A2(_07138_),
    .B1(_06977_),
    .B2(\datamem.data_ram[52][1] ),
    .C1(_07142_),
    .X(_07143_));
 sky130_fd_sc_hd__a221o_1 _19849_ (.A1(\datamem.data_ram[50][1] ),
    .A2(_06932_),
    .B1(_06958_),
    .B2(\datamem.data_ram[49][1] ),
    .C1(_06742_),
    .X(_07144_));
 sky130_fd_sc_hd__a221o_1 _19850_ (.A1(\datamem.data_ram[51][1] ),
    .A2(_06966_),
    .B1(_06927_),
    .B2(\datamem.data_ram[55][1] ),
    .C1(_07144_),
    .X(_07145_));
 sky130_fd_sc_hd__or2_1 _19851_ (.A(_07143_),
    .B(_07145_),
    .X(_07146_));
 sky130_fd_sc_hd__a22o_1 _19852_ (.A1(\datamem.data_ram[62][1] ),
    .A2(_07127_),
    .B1(_06970_),
    .B2(\datamem.data_ram[61][1] ),
    .X(_07147_));
 sky130_fd_sc_hd__a22o_1 _19853_ (.A1(\datamem.data_ram[58][1] ),
    .A2(_06932_),
    .B1(_06973_),
    .B2(\datamem.data_ram[56][1] ),
    .X(_07148_));
 sky130_fd_sc_hd__a221o_1 _19854_ (.A1(\datamem.data_ram[59][1] ),
    .A2(_06961_),
    .B1(_06948_),
    .B2(\datamem.data_ram[57][1] ),
    .C1(_07031_),
    .X(_07149_));
 sky130_fd_sc_hd__a211o_1 _19855_ (.A1(\datamem.data_ram[60][1] ),
    .A2(_06977_),
    .B1(_07148_),
    .C1(_07149_),
    .X(_07150_));
 sky130_fd_sc_hd__a211o_1 _19856_ (.A1(\datamem.data_ram[63][1] ),
    .A2(_07125_),
    .B1(_07147_),
    .C1(_07150_),
    .X(_07151_));
 sky130_fd_sc_hd__a31o_1 _19857_ (.A1(_07071_),
    .A2(_07146_),
    .A3(_07151_),
    .B1(_06985_),
    .X(_07152_));
 sky130_fd_sc_hd__a31o_1 _19858_ (.A1(_06916_),
    .A2(_07130_),
    .A3(_07141_),
    .B1(_07152_),
    .X(_07153_));
 sky130_fd_sc_hd__nand2_8 _19859_ (.A(_06750_),
    .B(_06860_),
    .Y(_07154_));
 sky130_fd_sc_hd__a22o_1 _19860_ (.A1(\datamem.data_ram[0][1] ),
    .A2(_06990_),
    .B1(_06966_),
    .B2(\datamem.data_ram[3][1] ),
    .X(_07155_));
 sky130_fd_sc_hd__a221o_1 _19861_ (.A1(\datamem.data_ram[5][1] ),
    .A2(_07132_),
    .B1(_07125_),
    .B2(\datamem.data_ram[7][1] ),
    .C1(_07155_),
    .X(_07156_));
 sky130_fd_sc_hd__a22o_1 _19862_ (.A1(\datamem.data_ram[6][1] ),
    .A2(_07127_),
    .B1(_06977_),
    .B2(\datamem.data_ram[4][1] ),
    .X(_07157_));
 sky130_fd_sc_hd__a221o_1 _19863_ (.A1(\datamem.data_ram[2][1] ),
    .A2(_07136_),
    .B1(_07133_),
    .B2(\datamem.data_ram[1][1] ),
    .C1(_07157_),
    .X(_07158_));
 sky130_fd_sc_hd__clkbuf_8 _19864_ (.A(_06978_),
    .X(_07159_));
 sky130_fd_sc_hd__a22o_1 _19865_ (.A1(\datamem.data_ram[14][1] ),
    .A2(_07159_),
    .B1(_06949_),
    .B2(\datamem.data_ram[9][1] ),
    .X(_07160_));
 sky130_fd_sc_hd__a22o_1 _19866_ (.A1(\datamem.data_ram[13][1] ),
    .A2(_06969_),
    .B1(_06926_),
    .B2(\datamem.data_ram[15][1] ),
    .X(_07161_));
 sky130_fd_sc_hd__a221o_1 _19867_ (.A1(\datamem.data_ram[10][1] ),
    .A2(_06932_),
    .B1(_06973_),
    .B2(\datamem.data_ram[8][1] ),
    .C1(_07031_),
    .X(_07162_));
 sky130_fd_sc_hd__a211o_1 _19868_ (.A1(\datamem.data_ram[11][1] ),
    .A2(_06966_),
    .B1(_07161_),
    .C1(_07162_),
    .X(_07163_));
 sky130_fd_sc_hd__a211o_1 _19869_ (.A1(\datamem.data_ram[12][1] ),
    .A2(_07123_),
    .B1(_07160_),
    .C1(_07163_),
    .X(_07164_));
 sky130_fd_sc_hd__o31a_1 _19870_ (.A1(_06604_),
    .A2(_07156_),
    .A3(_07158_),
    .B1(_07164_),
    .X(_07165_));
 sky130_fd_sc_hd__a22o_1 _19871_ (.A1(\datamem.data_ram[30][1] ),
    .A2(_07159_),
    .B1(_06949_),
    .B2(\datamem.data_ram[25][1] ),
    .X(_07166_));
 sky130_fd_sc_hd__a22o_1 _19872_ (.A1(\datamem.data_ram[26][1] ),
    .A2(_06989_),
    .B1(_06973_),
    .B2(\datamem.data_ram[24][1] ),
    .X(_07167_));
 sky130_fd_sc_hd__a221o_1 _19873_ (.A1(\datamem.data_ram[29][1] ),
    .A2(_06969_),
    .B1(_06943_),
    .B2(\datamem.data_ram[27][1] ),
    .C1(_07031_),
    .X(_07168_));
 sky130_fd_sc_hd__a211o_1 _19874_ (.A1(\datamem.data_ram[31][1] ),
    .A2(_06927_),
    .B1(_07167_),
    .C1(_07168_),
    .X(_07169_));
 sky130_fd_sc_hd__a211o_1 _19875_ (.A1(\datamem.data_ram[28][1] ),
    .A2(_07123_),
    .B1(_07166_),
    .C1(_07169_),
    .X(_07170_));
 sky130_fd_sc_hd__a22o_1 _19876_ (.A1(\datamem.data_ram[21][1] ),
    .A2(_06970_),
    .B1(_06977_),
    .B2(\datamem.data_ram[20][1] ),
    .X(_07171_));
 sky130_fd_sc_hd__a22o_1 _19877_ (.A1(\datamem.data_ram[18][1] ),
    .A2(_06931_),
    .B1(_06942_),
    .B2(\datamem.data_ram[19][1] ),
    .X(_07172_));
 sky130_fd_sc_hd__a221o_1 _19878_ (.A1(\datamem.data_ram[22][1] ),
    .A2(_06978_),
    .B1(_06973_),
    .B2(\datamem.data_ram[16][1] ),
    .C1(_07172_),
    .X(_07173_));
 sky130_fd_sc_hd__a211o_1 _19879_ (.A1(\datamem.data_ram[23][1] ),
    .A2(_06927_),
    .B1(_07173_),
    .C1(_07081_),
    .X(_07174_));
 sky130_fd_sc_hd__a211o_1 _19880_ (.A1(\datamem.data_ram[17][1] ),
    .A2(_06997_),
    .B1(_07171_),
    .C1(_07174_),
    .X(_07175_));
 sky130_fd_sc_hd__or2_2 _19881_ (.A(\rvcpu.dp.plem.ALUResultM[7] ),
    .B(_06750_),
    .X(_07176_));
 sky130_fd_sc_hd__clkbuf_8 _19882_ (.A(_07176_),
    .X(_07177_));
 sky130_fd_sc_hd__a21o_1 _19883_ (.A1(_07170_),
    .A2(_07175_),
    .B1(_07177_),
    .X(_07178_));
 sky130_fd_sc_hd__o211a_1 _19884_ (.A1(_07154_),
    .A2(_07165_),
    .B1(_07178_),
    .C1(_06988_),
    .X(_07179_));
 sky130_fd_sc_hd__o22a_1 _19885_ (.A1(\datamem.data_ram[24][17] ),
    .A2(_06698_),
    .B1(_07021_),
    .B2(\datamem.data_ram[31][17] ),
    .X(_07180_));
 sky130_fd_sc_hd__o221a_1 _19886_ (.A1(\datamem.data_ram[26][17] ),
    .A2(_06613_),
    .B1(_07077_),
    .B2(\datamem.data_ram[27][17] ),
    .C1(_07180_),
    .X(_07181_));
 sky130_fd_sc_hd__buf_4 _19887_ (.A(_06688_),
    .X(_07182_));
 sky130_fd_sc_hd__o22a_1 _19888_ (.A1(\datamem.data_ram[30][17] ),
    .A2(_06630_),
    .B1(_06665_),
    .B2(\datamem.data_ram[29][17] ),
    .X(_07183_));
 sky130_fd_sc_hd__o221a_1 _19889_ (.A1(\datamem.data_ram[28][17] ),
    .A2(_07182_),
    .B1(_06659_),
    .B2(\datamem.data_ram[25][17] ),
    .C1(_07183_),
    .X(_07184_));
 sky130_fd_sc_hd__o22a_1 _19890_ (.A1(\datamem.data_ram[18][17] ),
    .A2(_06612_),
    .B1(_06664_),
    .B2(\datamem.data_ram[21][17] ),
    .X(_07185_));
 sky130_fd_sc_hd__o221a_1 _19891_ (.A1(\datamem.data_ram[22][17] ),
    .A2(_06630_),
    .B1(_06701_),
    .B2(\datamem.data_ram[17][17] ),
    .C1(_07185_),
    .X(_07186_));
 sky130_fd_sc_hd__o22a_1 _19892_ (.A1(\datamem.data_ram[16][17] ),
    .A2(_06648_),
    .B1(_06707_),
    .B2(\datamem.data_ram[23][17] ),
    .X(_07187_));
 sky130_fd_sc_hd__o221a_1 _19893_ (.A1(\datamem.data_ram[19][17] ),
    .A2(_06739_),
    .B1(_06621_),
    .B2(\datamem.data_ram[20][17] ),
    .C1(_07187_),
    .X(_07188_));
 sky130_fd_sc_hd__and3_1 _19894_ (.A(_06681_),
    .B(_07186_),
    .C(_07188_),
    .X(_07189_));
 sky130_fd_sc_hd__a31o_1 _19895_ (.A1(_06604_),
    .A2(_07181_),
    .A3(_07184_),
    .B1(_07189_),
    .X(_07190_));
 sky130_fd_sc_hd__clkbuf_8 _19896_ (.A(_06698_),
    .X(_07191_));
 sky130_fd_sc_hd__o22a_1 _19897_ (.A1(\datamem.data_ram[6][17] ),
    .A2(_07028_),
    .B1(_06621_),
    .B2(\datamem.data_ram[4][17] ),
    .X(_07192_));
 sky130_fd_sc_hd__o22a_1 _19898_ (.A1(\datamem.data_ram[7][17] ),
    .A2(_07020_),
    .B1(_06658_),
    .B2(\datamem.data_ram[1][17] ),
    .X(_07193_));
 sky130_fd_sc_hd__o221a_1 _19899_ (.A1(\datamem.data_ram[2][17] ),
    .A2(_06612_),
    .B1(_06863_),
    .B2(\datamem.data_ram[3][17] ),
    .C1(_06776_),
    .X(_07194_));
 sky130_fd_sc_hd__o211a_1 _19900_ (.A1(\datamem.data_ram[5][17] ),
    .A2(_06665_),
    .B1(_07193_),
    .C1(_07194_),
    .X(_07195_));
 sky130_fd_sc_hd__o211a_1 _19901_ (.A1(\datamem.data_ram[0][17] ),
    .A2(_07191_),
    .B1(_07192_),
    .C1(_07195_),
    .X(_07196_));
 sky130_fd_sc_hd__o22a_1 _19902_ (.A1(\datamem.data_ram[10][17] ),
    .A2(_06613_),
    .B1(_06665_),
    .B2(\datamem.data_ram[13][17] ),
    .X(_07197_));
 sky130_fd_sc_hd__o22a_1 _19903_ (.A1(\datamem.data_ram[14][17] ),
    .A2(_06683_),
    .B1(_06648_),
    .B2(\datamem.data_ram[8][17] ),
    .X(_07198_));
 sky130_fd_sc_hd__o221a_1 _19904_ (.A1(\datamem.data_ram[11][17] ),
    .A2(_06863_),
    .B1(_07020_),
    .B2(\datamem.data_ram[15][17] ),
    .C1(_06602_),
    .X(_07199_));
 sky130_fd_sc_hd__o211a_1 _19905_ (.A1(\datamem.data_ram[9][17] ),
    .A2(_06659_),
    .B1(_07198_),
    .C1(_07199_),
    .X(_07200_));
 sky130_fd_sc_hd__o211a_1 _19906_ (.A1(\datamem.data_ram[12][17] ),
    .A2(_07182_),
    .B1(_07197_),
    .C1(_07200_),
    .X(_07201_));
 sky130_fd_sc_hd__o21a_1 _19907_ (.A1(_07196_),
    .A2(_07201_),
    .B1(_06596_),
    .X(_07202_));
 sky130_fd_sc_hd__clkbuf_8 _19908_ (.A(_07023_),
    .X(_07203_));
 sky130_fd_sc_hd__o22a_1 _19909_ (.A1(\datamem.data_ram[45][17] ),
    .A2(_06665_),
    .B1(_06701_),
    .B2(\datamem.data_ram[41][17] ),
    .X(_07204_));
 sky130_fd_sc_hd__o22a_1 _19910_ (.A1(\datamem.data_ram[46][17] ),
    .A2(_06628_),
    .B1(_06829_),
    .B2(\datamem.data_ram[43][17] ),
    .X(_07205_));
 sky130_fd_sc_hd__o221a_1 _19911_ (.A1(\datamem.data_ram[40][17] ),
    .A2(_06648_),
    .B1(_06707_),
    .B2(\datamem.data_ram[47][17] ),
    .C1(_07205_),
    .X(_07206_));
 sky130_fd_sc_hd__o211a_1 _19912_ (.A1(\datamem.data_ram[44][17] ),
    .A2(_06621_),
    .B1(_07206_),
    .C1(_07081_),
    .X(_07207_));
 sky130_fd_sc_hd__o211a_1 _19913_ (.A1(\datamem.data_ram[42][17] ),
    .A2(_07203_),
    .B1(_07204_),
    .C1(_07207_),
    .X(_07208_));
 sky130_fd_sc_hd__o22a_1 _19914_ (.A1(\datamem.data_ram[38][17] ),
    .A2(_06630_),
    .B1(_06621_),
    .B2(\datamem.data_ram[36][17] ),
    .X(_07209_));
 sky130_fd_sc_hd__o22a_1 _19915_ (.A1(\datamem.data_ram[37][17] ),
    .A2(_06664_),
    .B1(_06658_),
    .B2(\datamem.data_ram[33][17] ),
    .X(_07210_));
 sky130_fd_sc_hd__o221a_1 _19916_ (.A1(\datamem.data_ram[34][17] ),
    .A2(_06612_),
    .B1(_06863_),
    .B2(\datamem.data_ram[35][17] ),
    .C1(_06776_),
    .X(_07211_));
 sky130_fd_sc_hd__o211a_1 _19917_ (.A1(\datamem.data_ram[39][17] ),
    .A2(_07021_),
    .B1(_07210_),
    .C1(_07211_),
    .X(_07212_));
 sky130_fd_sc_hd__o211a_1 _19918_ (.A1(\datamem.data_ram[32][17] ),
    .A2(_07191_),
    .B1(_07209_),
    .C1(_07212_),
    .X(_07213_));
 sky130_fd_sc_hd__o22a_1 _19919_ (.A1(\datamem.data_ram[63][17] ),
    .A2(_07020_),
    .B1(_06620_),
    .B2(\datamem.data_ram[60][17] ),
    .X(_07214_));
 sky130_fd_sc_hd__o22a_1 _19920_ (.A1(\datamem.data_ram[61][17] ),
    .A2(_07037_),
    .B1(_06837_),
    .B2(\datamem.data_ram[56][17] ),
    .X(_07215_));
 sky130_fd_sc_hd__o221a_1 _19921_ (.A1(\datamem.data_ram[62][17] ),
    .A2(_06682_),
    .B1(_06790_),
    .B2(\datamem.data_ram[57][17] ),
    .C1(_06810_),
    .X(_07216_));
 sky130_fd_sc_hd__o211a_1 _19922_ (.A1(\datamem.data_ram[58][17] ),
    .A2(_06612_),
    .B1(_07215_),
    .C1(_07216_),
    .X(_07217_));
 sky130_fd_sc_hd__o211a_1 _19923_ (.A1(\datamem.data_ram[59][17] ),
    .A2(_06636_),
    .B1(_07214_),
    .C1(_07217_),
    .X(_07218_));
 sky130_fd_sc_hd__o22a_1 _19924_ (.A1(\datamem.data_ram[54][17] ),
    .A2(_06683_),
    .B1(_06664_),
    .B2(\datamem.data_ram[53][17] ),
    .X(_07219_));
 sky130_fd_sc_hd__o22a_1 _19925_ (.A1(\datamem.data_ram[48][17] ),
    .A2(_06807_),
    .B1(_06789_),
    .B2(\datamem.data_ram[49][17] ),
    .X(_07220_));
 sky130_fd_sc_hd__o221a_1 _19926_ (.A1(\datamem.data_ram[55][17] ),
    .A2(_06784_),
    .B1(_06806_),
    .B2(\datamem.data_ram[52][17] ),
    .C1(_07220_),
    .X(_07221_));
 sky130_fd_sc_hd__o211a_1 _19927_ (.A1(\datamem.data_ram[51][17] ),
    .A2(_06863_),
    .B1(_07221_),
    .C1(_06776_),
    .X(_07222_));
 sky130_fd_sc_hd__o211a_1 _19928_ (.A1(\datamem.data_ram[50][17] ),
    .A2(_06613_),
    .B1(_07219_),
    .C1(_07222_),
    .X(_07223_));
 sky130_fd_sc_hd__o31a_1 _19929_ (.A1(_06753_),
    .A2(_07218_),
    .A3(_07223_),
    .B1(_06713_),
    .X(_07224_));
 sky130_fd_sc_hd__o31a_1 _19930_ (.A1(_07071_),
    .A2(_07208_),
    .A3(_07213_),
    .B1(_07224_),
    .X(_07225_));
 sky130_fd_sc_hd__a211oi_4 _19931_ (.A1(_06797_),
    .A2(_07190_),
    .B1(_07202_),
    .C1(_07225_),
    .Y(_07226_));
 sky130_fd_sc_hd__o31a_1 _19932_ (.A1(\rvcpu.dp.plem.ALUResultM[0] ),
    .A2(_06586_),
    .A3(_06987_),
    .B1(_06915_),
    .X(_07227_));
 sky130_fd_sc_hd__o2bb2a_1 _19933_ (.A1_N(_07153_),
    .A2_N(_07179_),
    .B1(_07226_),
    .B2(_07227_),
    .X(_07228_));
 sky130_fd_sc_hd__o21ai_1 _19934_ (.A1(_06583_),
    .A2(_07121_),
    .B1(_07228_),
    .Y(_04426_));
 sky130_fd_sc_hd__o22a_1 _19935_ (.A1(\datamem.data_ram[37][18] ),
    .A2(_06703_),
    .B1(_06648_),
    .B2(\datamem.data_ram[32][18] ),
    .X(_07229_));
 sky130_fd_sc_hd__buf_6 _19936_ (.A(_06805_),
    .X(_07230_));
 sky130_fd_sc_hd__o22a_1 _19937_ (.A1(\datamem.data_ram[35][18] ),
    .A2(_06634_),
    .B1(_07230_),
    .B2(\datamem.data_ram[36][18] ),
    .X(_07231_));
 sky130_fd_sc_hd__o221a_1 _19938_ (.A1(\datamem.data_ram[39][18] ),
    .A2(_06760_),
    .B1(_06782_),
    .B2(\datamem.data_ram[33][18] ),
    .C1(_06769_),
    .X(_07232_));
 sky130_fd_sc_hd__o211a_1 _19939_ (.A1(\datamem.data_ram[38][18] ),
    .A2(_06629_),
    .B1(_07231_),
    .C1(_07232_),
    .X(_07233_));
 sky130_fd_sc_hd__o211a_1 _19940_ (.A1(\datamem.data_ram[34][18] ),
    .A2(_06613_),
    .B1(_07229_),
    .C1(_07233_),
    .X(_07234_));
 sky130_fd_sc_hd__o22a_1 _19941_ (.A1(\datamem.data_ram[45][18] ),
    .A2(_06664_),
    .B1(_06783_),
    .B2(\datamem.data_ram[41][18] ),
    .X(_07235_));
 sky130_fd_sc_hd__o22a_1 _19942_ (.A1(\datamem.data_ram[46][18] ),
    .A2(_06627_),
    .B1(_06803_),
    .B2(\datamem.data_ram[42][18] ),
    .X(_07236_));
 sky130_fd_sc_hd__o221a_1 _19943_ (.A1(\datamem.data_ram[40][18] ),
    .A2(_06778_),
    .B1(_06619_),
    .B2(\datamem.data_ram[44][18] ),
    .C1(_07236_),
    .X(_07237_));
 sky130_fd_sc_hd__o211a_1 _19944_ (.A1(\datamem.data_ram[47][18] ),
    .A2(_06707_),
    .B1(_07237_),
    .C1(_06602_),
    .X(_07238_));
 sky130_fd_sc_hd__o211a_1 _19945_ (.A1(\datamem.data_ram[43][18] ),
    .A2(_06636_),
    .B1(_07235_),
    .C1(_07238_),
    .X(_07239_));
 sky130_fd_sc_hd__o22a_1 _19946_ (.A1(\datamem.data_ram[53][18] ),
    .A2(_06702_),
    .B1(_06706_),
    .B2(\datamem.data_ram[55][18] ),
    .X(_07240_));
 sky130_fd_sc_hd__o22a_1 _19947_ (.A1(\datamem.data_ram[54][18] ),
    .A2(_07085_),
    .B1(_06646_),
    .B2(\datamem.data_ram[48][18] ),
    .X(_07241_));
 sky130_fd_sc_hd__buf_4 _19948_ (.A(_06653_),
    .X(_07242_));
 sky130_fd_sc_hd__clkbuf_8 _19949_ (.A(_07242_),
    .X(_07243_));
 sky130_fd_sc_hd__o221a_1 _19950_ (.A1(\datamem.data_ram[51][18] ),
    .A2(_06633_),
    .B1(_07243_),
    .B2(\datamem.data_ram[49][18] ),
    .C1(_06678_),
    .X(_07244_));
 sky130_fd_sc_hd__o211a_1 _19951_ (.A1(\datamem.data_ram[52][18] ),
    .A2(_06619_),
    .B1(_07241_),
    .C1(_07244_),
    .X(_07245_));
 sky130_fd_sc_hd__o211a_1 _19952_ (.A1(\datamem.data_ram[50][18] ),
    .A2(_06692_),
    .B1(_07240_),
    .C1(_07245_),
    .X(_07246_));
 sky130_fd_sc_hd__o22a_1 _19953_ (.A1(\datamem.data_ram[61][18] ),
    .A2(_06663_),
    .B1(_06782_),
    .B2(\datamem.data_ram[57][18] ),
    .X(_07247_));
 sky130_fd_sc_hd__o22a_1 _19954_ (.A1(\datamem.data_ram[59][18] ),
    .A2(_06632_),
    .B1(_06704_),
    .B2(\datamem.data_ram[63][18] ),
    .X(_07248_));
 sky130_fd_sc_hd__o221a_1 _19955_ (.A1(\datamem.data_ram[56][18] ),
    .A2(_06646_),
    .B1(_06765_),
    .B2(\datamem.data_ram[60][18] ),
    .C1(_07248_),
    .X(_07249_));
 sky130_fd_sc_hd__o211a_1 _19956_ (.A1(\datamem.data_ram[62][18] ),
    .A2(_06628_),
    .B1(_06601_),
    .C1(_07249_),
    .X(_07250_));
 sky130_fd_sc_hd__o211a_1 _19957_ (.A1(\datamem.data_ram[58][18] ),
    .A2(_06692_),
    .B1(_07247_),
    .C1(_07250_),
    .X(_07251_));
 sky130_fd_sc_hd__or3_1 _19958_ (.A(_06752_),
    .B(_07246_),
    .C(_07251_),
    .X(_07252_));
 sky130_fd_sc_hd__o311a_1 _19959_ (.A1(_06716_),
    .A2(_07234_),
    .A3(_07239_),
    .B1(_07252_),
    .C1(_06713_),
    .X(_07253_));
 sky130_fd_sc_hd__o22a_1 _19960_ (.A1(\datamem.data_ram[5][18] ),
    .A2(_06663_),
    .B1(_06784_),
    .B2(\datamem.data_ram[7][18] ),
    .X(_07254_));
 sky130_fd_sc_hd__o221a_1 _19961_ (.A1(\datamem.data_ram[2][18] ),
    .A2(_06612_),
    .B1(_06648_),
    .B2(\datamem.data_ram[0][18] ),
    .C1(_07254_),
    .X(_07255_));
 sky130_fd_sc_hd__o22a_1 _19962_ (.A1(\datamem.data_ram[6][18] ),
    .A2(_06628_),
    .B1(_06806_),
    .B2(\datamem.data_ram[4][18] ),
    .X(_07256_));
 sky130_fd_sc_hd__o221a_1 _19963_ (.A1(\datamem.data_ram[3][18] ),
    .A2(_06635_),
    .B1(_06783_),
    .B2(\datamem.data_ram[1][18] ),
    .C1(_07256_),
    .X(_07257_));
 sky130_fd_sc_hd__o22a_1 _19964_ (.A1(\datamem.data_ram[15][18] ),
    .A2(_06705_),
    .B1(_06781_),
    .B2(\datamem.data_ram[9][18] ),
    .X(_07258_));
 sky130_fd_sc_hd__o221a_1 _19965_ (.A1(\datamem.data_ram[14][18] ),
    .A2(_06763_),
    .B1(_06663_),
    .B2(\datamem.data_ram[13][18] ),
    .C1(_07258_),
    .X(_07259_));
 sky130_fd_sc_hd__o22a_1 _19966_ (.A1(\datamem.data_ram[10][18] ),
    .A2(_06610_),
    .B1(_06821_),
    .B2(\datamem.data_ram[8][18] ),
    .X(_07260_));
 sky130_fd_sc_hd__o221a_1 _19967_ (.A1(\datamem.data_ram[11][18] ),
    .A2(_06737_),
    .B1(_06619_),
    .B2(\datamem.data_ram[12][18] ),
    .C1(_07260_),
    .X(_07261_));
 sky130_fd_sc_hd__and3_1 _19968_ (.A(_06602_),
    .B(_07259_),
    .C(_07261_),
    .X(_07262_));
 sky130_fd_sc_hd__a31o_1 _19969_ (.A1(_06777_),
    .A2(_07255_),
    .A3(_07257_),
    .B1(_07262_),
    .X(_07263_));
 sky130_fd_sc_hd__o22a_1 _19970_ (.A1(\datamem.data_ram[30][18] ),
    .A2(_06763_),
    .B1(_06782_),
    .B2(\datamem.data_ram[25][18] ),
    .X(_07264_));
 sky130_fd_sc_hd__o22a_1 _19971_ (.A1(\datamem.data_ram[29][18] ),
    .A2(_06662_),
    .B1(_06646_),
    .B2(\datamem.data_ram[24][18] ),
    .X(_07265_));
 sky130_fd_sc_hd__o221a_1 _19972_ (.A1(\datamem.data_ram[26][18] ),
    .A2(_06690_),
    .B1(_06633_),
    .B2(\datamem.data_ram[27][18] ),
    .C1(_06600_),
    .X(_07266_));
 sky130_fd_sc_hd__o211a_1 _19973_ (.A1(\datamem.data_ram[28][18] ),
    .A2(_06619_),
    .B1(_07265_),
    .C1(_07266_),
    .X(_07267_));
 sky130_fd_sc_hd__o211a_1 _19974_ (.A1(\datamem.data_ram[31][18] ),
    .A2(_06707_),
    .B1(_07264_),
    .C1(_07267_),
    .X(_07268_));
 sky130_fd_sc_hd__o22a_1 _19975_ (.A1(\datamem.data_ram[23][18] ),
    .A2(_06706_),
    .B1(_07230_),
    .B2(\datamem.data_ram[20][18] ),
    .X(_07269_));
 sky130_fd_sc_hd__o22a_1 _19976_ (.A1(\datamem.data_ram[21][18] ),
    .A2(_06661_),
    .B1(_06780_),
    .B2(\datamem.data_ram[17][18] ),
    .X(_07270_));
 sky130_fd_sc_hd__o221a_1 _19977_ (.A1(\datamem.data_ram[22][18] ),
    .A2(_06744_),
    .B1(_06646_),
    .B2(\datamem.data_ram[16][18] ),
    .C1(_07270_),
    .X(_07271_));
 sky130_fd_sc_hd__o211a_1 _19978_ (.A1(\datamem.data_ram[19][18] ),
    .A2(_06634_),
    .B1(_07271_),
    .C1(_06679_),
    .X(_07272_));
 sky130_fd_sc_hd__o211a_1 _19979_ (.A1(\datamem.data_ram[18][18] ),
    .A2(_06612_),
    .B1(_07269_),
    .C1(_07272_),
    .X(_07273_));
 sky130_fd_sc_hd__or3_1 _19980_ (.A(_06752_),
    .B(_07268_),
    .C(_07273_),
    .X(_07274_));
 sky130_fd_sc_hd__o211a_1 _19981_ (.A1(_06716_),
    .A2(_07263_),
    .B1(_07274_),
    .C1(_06985_),
    .X(_07275_));
 sky130_fd_sc_hd__nor2_2 _19982_ (.A(_07253_),
    .B(_07275_),
    .Y(_07276_));
 sky130_fd_sc_hd__o21a_2 _19983_ (.A1(_06911_),
    .A2(_06580_),
    .B1(_06582_),
    .X(_07277_));
 sky130_fd_sc_hd__a22o_1 _19984_ (.A1(\datamem.data_ram[11][2] ),
    .A2(_06942_),
    .B1(_06925_),
    .B2(\datamem.data_ram[15][2] ),
    .X(_07278_));
 sky130_fd_sc_hd__a22o_1 _19985_ (.A1(\datamem.data_ram[10][2] ),
    .A2(_06930_),
    .B1(_06946_),
    .B2(\datamem.data_ram[9][2] ),
    .X(_07279_));
 sky130_fd_sc_hd__a221o_1 _19986_ (.A1(\datamem.data_ram[14][2] ),
    .A2(_06950_),
    .B1(_06919_),
    .B2(\datamem.data_ram[13][2] ),
    .C1(_07279_),
    .X(_07280_));
 sky130_fd_sc_hd__a211o_1 _19987_ (.A1(\datamem.data_ram[12][2] ),
    .A2(_06954_),
    .B1(_07280_),
    .C1(_06679_),
    .X(_07281_));
 sky130_fd_sc_hd__a211o_1 _19988_ (.A1(\datamem.data_ram[8][2] ),
    .A2(_06990_),
    .B1(_07278_),
    .C1(_07281_),
    .X(_07282_));
 sky130_fd_sc_hd__a22o_1 _19989_ (.A1(\datamem.data_ram[2][2] ),
    .A2(_06931_),
    .B1(_06920_),
    .B2(\datamem.data_ram[5][2] ),
    .X(_07283_));
 sky130_fd_sc_hd__a22o_1 _19990_ (.A1(\datamem.data_ram[4][2] ),
    .A2(_06953_),
    .B1(_06946_),
    .B2(\datamem.data_ram[1][2] ),
    .X(_07284_));
 sky130_fd_sc_hd__a221o_1 _19991_ (.A1(\datamem.data_ram[6][2] ),
    .A2(_06950_),
    .B1(_06924_),
    .B2(\datamem.data_ram[7][2] ),
    .C1(_07284_),
    .X(_07285_));
 sky130_fd_sc_hd__a211o_1 _19992_ (.A1(\datamem.data_ram[3][2] ),
    .A2(_06942_),
    .B1(_07285_),
    .C1(_06601_),
    .X(_07286_));
 sky130_fd_sc_hd__a211o_1 _19993_ (.A1(\datamem.data_ram[0][2] ),
    .A2(_06973_),
    .B1(_07283_),
    .C1(_07286_),
    .X(_07287_));
 sky130_fd_sc_hd__a22o_1 _19994_ (.A1(\datamem.data_ram[22][2] ),
    .A2(_06951_),
    .B1(_06936_),
    .B2(\datamem.data_ram[16][2] ),
    .X(_07288_));
 sky130_fd_sc_hd__a22o_1 _19995_ (.A1(\datamem.data_ram[18][2] ),
    .A2(_06930_),
    .B1(_06924_),
    .B2(\datamem.data_ram[23][2] ),
    .X(_07289_));
 sky130_fd_sc_hd__a221o_1 _19996_ (.A1(\datamem.data_ram[21][2] ),
    .A2(_06919_),
    .B1(_06953_),
    .B2(\datamem.data_ram[20][2] ),
    .C1(_07289_),
    .X(_07290_));
 sky130_fd_sc_hd__a211o_1 _19997_ (.A1(\datamem.data_ram[17][2] ),
    .A2(_06947_),
    .B1(_07290_),
    .C1(_06851_),
    .X(_07291_));
 sky130_fd_sc_hd__a211o_1 _19998_ (.A1(\datamem.data_ram[19][2] ),
    .A2(_06942_),
    .B1(_07288_),
    .C1(_07291_),
    .X(_07292_));
 sky130_fd_sc_hd__a22o_1 _19999_ (.A1(\datamem.data_ram[30][2] ),
    .A2(_06950_),
    .B1(_06947_),
    .B2(\datamem.data_ram[25][2] ),
    .X(_07293_));
 sky130_fd_sc_hd__a22o_1 _20000_ (.A1(\datamem.data_ram[29][2] ),
    .A2(_06919_),
    .B1(_06953_),
    .B2(\datamem.data_ram[28][2] ),
    .X(_07294_));
 sky130_fd_sc_hd__a221o_1 _20001_ (.A1(\datamem.data_ram[26][2] ),
    .A2(_06930_),
    .B1(_06924_),
    .B2(\datamem.data_ram[31][2] ),
    .C1(_06677_),
    .X(_07295_));
 sky130_fd_sc_hd__a211o_1 _20002_ (.A1(\datamem.data_ram[24][2] ),
    .A2(_06936_),
    .B1(_07294_),
    .C1(_07295_),
    .X(_07296_));
 sky130_fd_sc_hd__a211o_2 _20003_ (.A1(\datamem.data_ram[27][2] ),
    .A2(_06942_),
    .B1(_07293_),
    .C1(_07296_),
    .X(_07297_));
 sky130_fd_sc_hd__a31o_1 _20004_ (.A1(_06714_),
    .A2(_07292_),
    .A3(_07297_),
    .B1(_06594_),
    .X(_07298_));
 sky130_fd_sc_hd__a31o_1 _20005_ (.A1(_06752_),
    .A2(_07282_),
    .A3(_07287_),
    .B1(_07298_),
    .X(_07299_));
 sky130_fd_sc_hd__a22o_1 _20006_ (.A1(\datamem.data_ram[58][2] ),
    .A2(_06930_),
    .B1(_06924_),
    .B2(\datamem.data_ram[63][2] ),
    .X(_07300_));
 sky130_fd_sc_hd__a221o_1 _20007_ (.A1(\datamem.data_ram[61][2] ),
    .A2(_06920_),
    .B1(_06942_),
    .B2(\datamem.data_ram[59][2] ),
    .C1(_07300_),
    .X(_07301_));
 sky130_fd_sc_hd__a22o_1 _20008_ (.A1(\datamem.data_ram[56][2] ),
    .A2(_06936_),
    .B1(_06953_),
    .B2(\datamem.data_ram[60][2] ),
    .X(_07302_));
 sky130_fd_sc_hd__a211o_1 _20009_ (.A1(\datamem.data_ram[62][2] ),
    .A2(_06951_),
    .B1(_06769_),
    .C1(_07302_),
    .X(_07303_));
 sky130_fd_sc_hd__a211o_1 _20010_ (.A1(\datamem.data_ram[57][2] ),
    .A2(_06948_),
    .B1(_07301_),
    .C1(_07303_),
    .X(_07304_));
 sky130_fd_sc_hd__a22o_1 _20011_ (.A1(\datamem.data_ram[48][2] ),
    .A2(_06937_),
    .B1(_06954_),
    .B2(\datamem.data_ram[52][2] ),
    .X(_07305_));
 sky130_fd_sc_hd__a22o_1 _20012_ (.A1(\datamem.data_ram[54][2] ),
    .A2(_06950_),
    .B1(_06930_),
    .B2(\datamem.data_ram[50][2] ),
    .X(_07306_));
 sky130_fd_sc_hd__a221o_1 _20013_ (.A1(\datamem.data_ram[51][2] ),
    .A2(_06941_),
    .B1(_06947_),
    .B2(\datamem.data_ram[49][2] ),
    .C1(_06600_),
    .X(_07307_));
 sky130_fd_sc_hd__a211o_1 _20014_ (.A1(\datamem.data_ram[53][2] ),
    .A2(_06920_),
    .B1(_07306_),
    .C1(_07307_),
    .X(_07308_));
 sky130_fd_sc_hd__a211o_1 _20015_ (.A1(\datamem.data_ram[55][2] ),
    .A2(_06926_),
    .B1(_07305_),
    .C1(_07308_),
    .X(_07309_));
 sky130_fd_sc_hd__a22o_1 _20016_ (.A1(\datamem.data_ram[37][2] ),
    .A2(_06919_),
    .B1(_06947_),
    .B2(\datamem.data_ram[33][2] ),
    .X(_07310_));
 sky130_fd_sc_hd__a22o_1 _20017_ (.A1(\datamem.data_ram[35][2] ),
    .A2(_06941_),
    .B1(_06924_),
    .B2(\datamem.data_ram[39][2] ),
    .X(_07311_));
 sky130_fd_sc_hd__a221o_1 _20018_ (.A1(\datamem.data_ram[32][2] ),
    .A2(_06935_),
    .B1(_06953_),
    .B2(\datamem.data_ram[36][2] ),
    .C1(_07311_),
    .X(_07312_));
 sky130_fd_sc_hd__a211o_1 _20019_ (.A1(\datamem.data_ram[34][2] ),
    .A2(_06930_),
    .B1(_06600_),
    .C1(_07312_),
    .X(_07313_));
 sky130_fd_sc_hd__a211o_1 _20020_ (.A1(\datamem.data_ram[38][2] ),
    .A2(_06951_),
    .B1(_07310_),
    .C1(_07313_),
    .X(_07314_));
 sky130_fd_sc_hd__a22o_1 _20021_ (.A1(\datamem.data_ram[46][2] ),
    .A2(_06950_),
    .B1(_06953_),
    .B2(\datamem.data_ram[44][2] ),
    .X(_07315_));
 sky130_fd_sc_hd__a221o_1 _20022_ (.A1(\datamem.data_ram[40][2] ),
    .A2(_06935_),
    .B1(_06946_),
    .B2(\datamem.data_ram[41][2] ),
    .C1(_07315_),
    .X(_07316_));
 sky130_fd_sc_hd__a22o_1 _20023_ (.A1(\datamem.data_ram[42][2] ),
    .A2(_06930_),
    .B1(_06924_),
    .B2(\datamem.data_ram[47][2] ),
    .X(_07317_));
 sky130_fd_sc_hd__a221o_1 _20024_ (.A1(\datamem.data_ram[45][2] ),
    .A2(_06919_),
    .B1(_06941_),
    .B2(\datamem.data_ram[43][2] ),
    .C1(_07317_),
    .X(_07318_));
 sky130_fd_sc_hd__or3_1 _20025_ (.A(_06769_),
    .B(_07316_),
    .C(_07318_),
    .X(_07319_));
 sky130_fd_sc_hd__a31o_1 _20026_ (.A1(_06752_),
    .A2(_07314_),
    .A3(_07319_),
    .B1(_06860_),
    .X(_07320_));
 sky130_fd_sc_hd__a31o_1 _20027_ (.A1(_06715_),
    .A2(_07304_),
    .A3(_07309_),
    .B1(_07320_),
    .X(_07321_));
 sky130_fd_sc_hd__nand2_1 _20028_ (.A(_07299_),
    .B(_07321_),
    .Y(_07322_));
 sky130_fd_sc_hd__or3b_1 _20029_ (.A(_06911_),
    .B(_07322_),
    .C_N(_06588_),
    .X(_07323_));
 sky130_fd_sc_hd__o22a_1 _20030_ (.A1(\datamem.data_ram[30][26] ),
    .A2(_06763_),
    .B1(_06766_),
    .B2(\datamem.data_ram[28][26] ),
    .X(_07324_));
 sky130_fd_sc_hd__o22a_1 _20031_ (.A1(\datamem.data_ram[26][26] ),
    .A2(_06609_),
    .B1(_06632_),
    .B2(\datamem.data_ram[27][26] ),
    .X(_07325_));
 sky130_fd_sc_hd__o221a_1 _20032_ (.A1(\datamem.data_ram[24][26] ),
    .A2(_06695_),
    .B1(_07243_),
    .B2(\datamem.data_ram[25][26] ),
    .C1(_07325_),
    .X(_07326_));
 sky130_fd_sc_hd__o211a_1 _20033_ (.A1(\datamem.data_ram[29][26] ),
    .A2(_06702_),
    .B1(_06741_),
    .C1(_07326_),
    .X(_07327_));
 sky130_fd_sc_hd__o211a_1 _20034_ (.A1(\datamem.data_ram[31][26] ),
    .A2(_06761_),
    .B1(_07324_),
    .C1(_07327_),
    .X(_07328_));
 sky130_fd_sc_hd__o22a_1 _20035_ (.A1(\datamem.data_ram[16][26] ),
    .A2(_06778_),
    .B1(_06699_),
    .B2(\datamem.data_ram[17][26] ),
    .X(_07329_));
 sky130_fd_sc_hd__o22a_1 _20036_ (.A1(\datamem.data_ram[22][26] ),
    .A2(_07085_),
    .B1(_06705_),
    .B2(\datamem.data_ram[23][26] ),
    .X(_07330_));
 sky130_fd_sc_hd__o221a_1 _20037_ (.A1(\datamem.data_ram[18][26] ),
    .A2(_06690_),
    .B1(_06662_),
    .B2(\datamem.data_ram[21][26] ),
    .C1(_06678_),
    .X(_07331_));
 sky130_fd_sc_hd__o211a_1 _20038_ (.A1(\datamem.data_ram[20][26] ),
    .A2(_06619_),
    .B1(_07330_),
    .C1(_07331_),
    .X(_07332_));
 sky130_fd_sc_hd__o211a_1 _20039_ (.A1(\datamem.data_ram[19][26] ),
    .A2(_06635_),
    .B1(_07329_),
    .C1(_07332_),
    .X(_07333_));
 sky130_fd_sc_hd__o22a_1 _20040_ (.A1(\datamem.data_ram[6][26] ),
    .A2(_06744_),
    .B1(_06765_),
    .B2(\datamem.data_ram[4][26] ),
    .X(_07334_));
 sky130_fd_sc_hd__o22a_1 _20041_ (.A1(\datamem.data_ram[0][26] ),
    .A2(_06645_),
    .B1(_07242_),
    .B2(\datamem.data_ram[1][26] ),
    .X(_07335_));
 sky130_fd_sc_hd__o221a_1 _20042_ (.A1(\datamem.data_ram[3][26] ),
    .A2(_06729_),
    .B1(_06668_),
    .B2(\datamem.data_ram[7][26] ),
    .C1(_06677_),
    .X(_07336_));
 sky130_fd_sc_hd__o211a_1 _20043_ (.A1(\datamem.data_ram[5][26] ),
    .A2(_06722_),
    .B1(_07335_),
    .C1(_07336_),
    .X(_07337_));
 sky130_fd_sc_hd__o211a_1 _20044_ (.A1(\datamem.data_ram[2][26] ),
    .A2(_06691_),
    .B1(_07334_),
    .C1(_07337_),
    .X(_07338_));
 sky130_fd_sc_hd__o22a_1 _20045_ (.A1(\datamem.data_ram[14][26] ),
    .A2(_06744_),
    .B1(_07243_),
    .B2(\datamem.data_ram[9][26] ),
    .X(_07339_));
 sky130_fd_sc_hd__o22a_1 _20046_ (.A1(\datamem.data_ram[8][26] ),
    .A2(_06820_),
    .B1(_06632_),
    .B2(\datamem.data_ram[11][26] ),
    .X(_07340_));
 sky130_fd_sc_hd__o221a_1 _20047_ (.A1(\datamem.data_ram[10][26] ),
    .A2(_06609_),
    .B1(_06617_),
    .B2(\datamem.data_ram[12][26] ),
    .C1(_06598_),
    .X(_07341_));
 sky130_fd_sc_hd__o211a_1 _20048_ (.A1(\datamem.data_ram[13][26] ),
    .A2(_06662_),
    .B1(_07340_),
    .C1(_07341_),
    .X(_07342_));
 sky130_fd_sc_hd__o211a_1 _20049_ (.A1(\datamem.data_ram[15][26] ),
    .A2(_06760_),
    .B1(_07339_),
    .C1(_07342_),
    .X(_07343_));
 sky130_fd_sc_hd__o22a_1 _20050_ (.A1(\datamem.data_ram[34][26] ),
    .A2(_06608_),
    .B1(_06644_),
    .B2(\datamem.data_ram[32][26] ),
    .X(_07344_));
 sky130_fd_sc_hd__o221a_1 _20051_ (.A1(\datamem.data_ram[37][26] ),
    .A2(_06721_),
    .B1(_06668_),
    .B2(\datamem.data_ram[39][26] ),
    .C1(_07344_),
    .X(_07345_));
 sky130_fd_sc_hd__o22a_1 _20052_ (.A1(\datamem.data_ram[38][26] ),
    .A2(_06624_),
    .B1(_06616_),
    .B2(\datamem.data_ram[36][26] ),
    .X(_07346_));
 sky130_fd_sc_hd__o221a_1 _20053_ (.A1(\datamem.data_ram[35][26] ),
    .A2(_06729_),
    .B1(_07242_),
    .B2(\datamem.data_ram[33][26] ),
    .C1(_07346_),
    .X(_07347_));
 sky130_fd_sc_hd__and3_1 _20054_ (.A(_06678_),
    .B(_07345_),
    .C(_07347_),
    .X(_07348_));
 sky130_fd_sc_hd__o22a_1 _20055_ (.A1(\datamem.data_ram[43][26] ),
    .A2(_06631_),
    .B1(_06684_),
    .B2(\datamem.data_ram[44][26] ),
    .X(_07349_));
 sky130_fd_sc_hd__o221a_1 _20056_ (.A1(\datamem.data_ram[42][26] ),
    .A2(_06609_),
    .B1(_06704_),
    .B2(\datamem.data_ram[47][26] ),
    .C1(_07349_),
    .X(_07350_));
 sky130_fd_sc_hd__o22a_1 _20057_ (.A1(\datamem.data_ram[45][26] ),
    .A2(_06660_),
    .B1(_06644_),
    .B2(\datamem.data_ram[40][26] ),
    .X(_07351_));
 sky130_fd_sc_hd__o221a_1 _20058_ (.A1(\datamem.data_ram[46][26] ),
    .A2(_06743_),
    .B1(_07242_),
    .B2(\datamem.data_ram[41][26] ),
    .C1(_07351_),
    .X(_07352_));
 sky130_fd_sc_hd__a31o_1 _20059_ (.A1(_06600_),
    .A2(_07350_),
    .A3(_07352_),
    .B1(_06592_),
    .X(_07353_));
 sky130_fd_sc_hd__o221a_1 _20060_ (.A1(\datamem.data_ram[62][26] ),
    .A2(_06743_),
    .B1(_06704_),
    .B2(\datamem.data_ram[63][26] ),
    .C1(_06598_),
    .X(_07354_));
 sky130_fd_sc_hd__or2_1 _20061_ (.A(\datamem.data_ram[59][26] ),
    .B(_06631_),
    .X(_07355_));
 sky130_fd_sc_hd__o221a_1 _20062_ (.A1(\datamem.data_ram[60][26] ),
    .A2(_06684_),
    .B1(_07242_),
    .B2(\datamem.data_ram[57][26] ),
    .C1(_07355_),
    .X(_07356_));
 sky130_fd_sc_hd__or2_1 _20063_ (.A(\datamem.data_ram[58][26] ),
    .B(_06608_),
    .X(_07357_));
 sky130_fd_sc_hd__o221a_1 _20064_ (.A1(\datamem.data_ram[61][26] ),
    .A2(_06721_),
    .B1(_06645_),
    .B2(\datamem.data_ram[56][26] ),
    .C1(_07357_),
    .X(_07358_));
 sky130_fd_sc_hd__and3_1 _20065_ (.A(_07354_),
    .B(_07356_),
    .C(_07358_),
    .X(_07359_));
 sky130_fd_sc_hd__o22a_1 _20066_ (.A1(\datamem.data_ram[50][26] ),
    .A2(_06608_),
    .B1(_06660_),
    .B2(\datamem.data_ram[53][26] ),
    .X(_07360_));
 sky130_fd_sc_hd__o221a_1 _20067_ (.A1(\datamem.data_ram[48][26] ),
    .A2(_06645_),
    .B1(_06617_),
    .B2(\datamem.data_ram[52][26] ),
    .C1(_07360_),
    .X(_07361_));
 sky130_fd_sc_hd__o22a_1 _20068_ (.A1(\datamem.data_ram[54][26] ),
    .A2(_06625_),
    .B1(_06631_),
    .B2(\datamem.data_ram[51][26] ),
    .X(_07362_));
 sky130_fd_sc_hd__o221a_1 _20069_ (.A1(\datamem.data_ram[55][26] ),
    .A2(_06704_),
    .B1(_07242_),
    .B2(\datamem.data_ram[49][26] ),
    .C1(_07362_),
    .X(_07363_));
 sky130_fd_sc_hd__a31o_1 _20070_ (.A1(_06678_),
    .A2(_07361_),
    .A3(_07363_),
    .B1(_06750_),
    .X(_07364_));
 sky130_fd_sc_hd__o22a_1 _20071_ (.A1(_07348_),
    .A2(_07353_),
    .B1(_07359_),
    .B2(_07364_),
    .X(_07365_));
 sky130_fd_sc_hd__o32a_1 _20072_ (.A1(_07154_),
    .A2(_07338_),
    .A3(_07343_),
    .B1(_07365_),
    .B2(_06860_),
    .X(_07366_));
 sky130_fd_sc_hd__o31a_4 _20073_ (.A1(_07177_),
    .A2(_07328_),
    .A3(_07333_),
    .B1(_07366_),
    .X(_07367_));
 sky130_fd_sc_hd__inv_2 _20074_ (.A(_07367_),
    .Y(_07368_));
 sky130_fd_sc_hd__o22a_1 _20075_ (.A1(\datamem.data_ram[46][10] ),
    .A2(_06718_),
    .B1(_06656_),
    .B2(\datamem.data_ram[41][10] ),
    .X(_07369_));
 sky130_fd_sc_hd__o221a_1 _20076_ (.A1(\datamem.data_ram[45][10] ),
    .A2(_07037_),
    .B1(_06837_),
    .B2(\datamem.data_ram[40][10] ),
    .C1(_07369_),
    .X(_07370_));
 sky130_fd_sc_hd__o22a_1 _20077_ (.A1(\datamem.data_ram[42][10] ),
    .A2(_06803_),
    .B1(_06726_),
    .B2(\datamem.data_ram[47][10] ),
    .X(_07371_));
 sky130_fd_sc_hd__o221a_1 _20078_ (.A1(\datamem.data_ram[43][10] ),
    .A2(_06829_),
    .B1(_06806_),
    .B2(\datamem.data_ram[44][10] ),
    .C1(_07371_),
    .X(_07372_));
 sky130_fd_sc_hd__o22a_1 _20079_ (.A1(\datamem.data_ram[38][10] ),
    .A2(_06717_),
    .B1(_06812_),
    .B2(\datamem.data_ram[35][10] ),
    .X(_07373_));
 sky130_fd_sc_hd__o221a_1 _20080_ (.A1(\datamem.data_ram[34][10] ),
    .A2(_06803_),
    .B1(_06805_),
    .B2(\datamem.data_ram[36][10] ),
    .C1(_07373_),
    .X(_07374_));
 sky130_fd_sc_hd__o22a_1 _20081_ (.A1(\datamem.data_ram[37][10] ),
    .A2(_06722_),
    .B1(_06669_),
    .B2(\datamem.data_ram[39][10] ),
    .X(_07375_));
 sky130_fd_sc_hd__o221a_1 _20082_ (.A1(\datamem.data_ram[32][10] ),
    .A2(_06821_),
    .B1(_06789_),
    .B2(\datamem.data_ram[33][10] ),
    .C1(_07375_),
    .X(_07376_));
 sky130_fd_sc_hd__and3_1 _20083_ (.A(_06679_),
    .B(_07374_),
    .C(_07376_),
    .X(_07377_));
 sky130_fd_sc_hd__a31o_1 _20084_ (.A1(_06602_),
    .A2(_07370_),
    .A3(_07372_),
    .B1(_07377_),
    .X(_07378_));
 sky130_fd_sc_hd__o22a_1 _20085_ (.A1(\datamem.data_ram[53][10] ),
    .A2(_06823_),
    .B1(_06670_),
    .B2(\datamem.data_ram[55][10] ),
    .X(_07379_));
 sky130_fd_sc_hd__o22a_1 _20086_ (.A1(\datamem.data_ram[54][10] ),
    .A2(_06626_),
    .B1(_06811_),
    .B2(\datamem.data_ram[48][10] ),
    .X(_07380_));
 sky130_fd_sc_hd__o221a_1 _20087_ (.A1(\datamem.data_ram[50][10] ),
    .A2(_06802_),
    .B1(_06780_),
    .B2(\datamem.data_ram[49][10] ),
    .C1(_06732_),
    .X(_07381_));
 sky130_fd_sc_hd__o211a_1 _20088_ (.A1(\datamem.data_ram[52][10] ),
    .A2(_06805_),
    .B1(_07380_),
    .C1(_07381_),
    .X(_07382_));
 sky130_fd_sc_hd__o211a_1 _20089_ (.A1(\datamem.data_ram[51][10] ),
    .A2(_06829_),
    .B1(_07379_),
    .C1(_07382_),
    .X(_07383_));
 sky130_fd_sc_hd__o22a_1 _20090_ (.A1(\datamem.data_ram[62][10] ),
    .A2(_06627_),
    .B1(_06723_),
    .B2(\datamem.data_ram[61][10] ),
    .X(_07384_));
 sky130_fd_sc_hd__o22a_1 _20091_ (.A1(\datamem.data_ram[58][10] ),
    .A2(_06689_),
    .B1(_06668_),
    .B2(\datamem.data_ram[63][10] ),
    .X(_07385_));
 sky130_fd_sc_hd__o221a_1 _20092_ (.A1(\datamem.data_ram[56][10] ),
    .A2(_06811_),
    .B1(_06685_),
    .B2(\datamem.data_ram[60][10] ),
    .C1(_07385_),
    .X(_07386_));
 sky130_fd_sc_hd__o211a_1 _20093_ (.A1(\datamem.data_ram[59][10] ),
    .A2(_06828_),
    .B1(_07386_),
    .C1(_06851_),
    .X(_07387_));
 sky130_fd_sc_hd__o211a_1 _20094_ (.A1(\datamem.data_ram[57][10] ),
    .A2(_06790_),
    .B1(_07384_),
    .C1(_07387_),
    .X(_07388_));
 sky130_fd_sc_hd__or3_1 _20095_ (.A(_06751_),
    .B(_07383_),
    .C(_07388_),
    .X(_07389_));
 sky130_fd_sc_hd__o211a_1 _20096_ (.A1(_06715_),
    .A2(_07378_),
    .B1(_07389_),
    .C1(_06712_),
    .X(_07390_));
 sky130_fd_sc_hd__o22a_1 _20097_ (.A1(\datamem.data_ram[2][10] ),
    .A2(_06804_),
    .B1(_06687_),
    .B2(\datamem.data_ram[4][10] ),
    .X(_07391_));
 sky130_fd_sc_hd__o22a_1 _20098_ (.A1(\datamem.data_ram[6][10] ),
    .A2(_06718_),
    .B1(_06656_),
    .B2(\datamem.data_ram[1][10] ),
    .X(_07392_));
 sky130_fd_sc_hd__o221a_1 _20099_ (.A1(\datamem.data_ram[5][10] ),
    .A2(_06723_),
    .B1(_06828_),
    .B2(\datamem.data_ram[3][10] ),
    .C1(_06733_),
    .X(_07393_));
 sky130_fd_sc_hd__o211a_1 _20100_ (.A1(\datamem.data_ram[0][10] ),
    .A2(_06837_),
    .B1(_07392_),
    .C1(_07393_),
    .X(_07394_));
 sky130_fd_sc_hd__o211a_1 _20101_ (.A1(\datamem.data_ram[7][10] ),
    .A2(_07020_),
    .B1(_07391_),
    .C1(_07394_),
    .X(_07395_));
 sky130_fd_sc_hd__o22a_1 _20102_ (.A1(\datamem.data_ram[13][10] ),
    .A2(_06724_),
    .B1(_06697_),
    .B2(\datamem.data_ram[8][10] ),
    .X(_07396_));
 sky130_fd_sc_hd__o22a_1 _20103_ (.A1(\datamem.data_ram[14][10] ),
    .A2(_06717_),
    .B1(_06730_),
    .B2(\datamem.data_ram[11][10] ),
    .X(_07397_));
 sky130_fd_sc_hd__o221a_1 _20104_ (.A1(\datamem.data_ram[12][10] ),
    .A2(_06686_),
    .B1(_06656_),
    .B2(\datamem.data_ram[9][10] ),
    .C1(_07397_),
    .X(_07398_));
 sky130_fd_sc_hd__o211a_1 _20105_ (.A1(\datamem.data_ram[10][10] ),
    .A2(_06754_),
    .B1(_06810_),
    .C1(_07398_),
    .X(_07399_));
 sky130_fd_sc_hd__o211a_1 _20106_ (.A1(\datamem.data_ram[15][10] ),
    .A2(_06672_),
    .B1(_07396_),
    .C1(_07399_),
    .X(_07400_));
 sky130_fd_sc_hd__o22a_1 _20107_ (.A1(\datamem.data_ram[16][10] ),
    .A2(_06696_),
    .B1(_06656_),
    .B2(\datamem.data_ram[17][10] ),
    .X(_07401_));
 sky130_fd_sc_hd__o22a_1 _20108_ (.A1(\datamem.data_ram[22][10] ),
    .A2(_06717_),
    .B1(_06669_),
    .B2(\datamem.data_ram[23][10] ),
    .X(_07402_));
 sky130_fd_sc_hd__o221a_1 _20109_ (.A1(\datamem.data_ram[19][10] ),
    .A2(_06812_),
    .B1(_06685_),
    .B2(\datamem.data_ram[20][10] ),
    .C1(_06732_),
    .X(_07403_));
 sky130_fd_sc_hd__o211a_1 _20110_ (.A1(\datamem.data_ram[21][10] ),
    .A2(_06723_),
    .B1(_07402_),
    .C1(_07403_),
    .X(_07404_));
 sky130_fd_sc_hd__o211a_1 _20111_ (.A1(\datamem.data_ram[18][10] ),
    .A2(_06804_),
    .B1(_07401_),
    .C1(_07404_),
    .X(_07405_));
 sky130_fd_sc_hd__o22a_1 _20112_ (.A1(\datamem.data_ram[29][10] ),
    .A2(_06723_),
    .B1(_06686_),
    .B2(\datamem.data_ram[28][10] ),
    .X(_07406_));
 sky130_fd_sc_hd__o22a_1 _20113_ (.A1(\datamem.data_ram[26][10] ),
    .A2(_06689_),
    .B1(_06645_),
    .B2(\datamem.data_ram[24][10] ),
    .X(_07407_));
 sky130_fd_sc_hd__o221a_1 _20114_ (.A1(\datamem.data_ram[30][10] ),
    .A2(_06626_),
    .B1(_06669_),
    .B2(\datamem.data_ram[31][10] ),
    .C1(_07407_),
    .X(_07408_));
 sky130_fd_sc_hd__o211a_1 _20115_ (.A1(\datamem.data_ram[27][10] ),
    .A2(_06731_),
    .B1(_07408_),
    .C1(_06741_),
    .X(_07409_));
 sky130_fd_sc_hd__o211a_1 _20116_ (.A1(\datamem.data_ram[25][10] ),
    .A2(_06657_),
    .B1(_07406_),
    .C1(_07409_),
    .X(_07410_));
 sky130_fd_sc_hd__or3_1 _20117_ (.A(_06752_),
    .B(_07405_),
    .C(_07410_),
    .X(_07411_));
 sky130_fd_sc_hd__o311a_1 _20118_ (.A1(_06715_),
    .A2(_07395_),
    .A3(_07400_),
    .B1(_06860_),
    .C1(_07411_),
    .X(_07412_));
 sky130_fd_sc_hd__nor2_4 _20119_ (.A(_07390_),
    .B(_07412_),
    .Y(_07413_));
 sky130_fd_sc_hd__o32a_1 _20120_ (.A1(_05391_),
    .A2(_06586_),
    .A3(_07368_),
    .B1(_07413_),
    .B2(_07120_),
    .X(_07414_));
 sky130_fd_sc_hd__o211a_1 _20121_ (.A1(_06912_),
    .A2(_07276_),
    .B1(_07323_),
    .C1(_07414_),
    .X(_07415_));
 sky130_fd_sc_hd__o22a_1 _20122_ (.A1(_07277_),
    .A2(_07322_),
    .B1(_07415_),
    .B2(_06583_),
    .X(_07416_));
 sky130_fd_sc_hd__o21ai_1 _20123_ (.A1(_06915_),
    .A2(_07276_),
    .B1(_07416_),
    .Y(_04437_));
 sky130_fd_sc_hd__o22a_1 _20124_ (.A1(\datamem.data_ram[6][27] ),
    .A2(_06719_),
    .B1(_06754_),
    .B2(\datamem.data_ram[2][27] ),
    .X(_07417_));
 sky130_fd_sc_hd__o221a_1 _20125_ (.A1(\datamem.data_ram[5][27] ),
    .A2(_06664_),
    .B1(_06648_),
    .B2(\datamem.data_ram[0][27] ),
    .C1(_07417_),
    .X(_07418_));
 sky130_fd_sc_hd__o22a_1 _20126_ (.A1(\datamem.data_ram[7][27] ),
    .A2(_06671_),
    .B1(_06657_),
    .B2(\datamem.data_ram[1][27] ),
    .X(_07419_));
 sky130_fd_sc_hd__o221a_1 _20127_ (.A1(\datamem.data_ram[3][27] ),
    .A2(_06863_),
    .B1(_06620_),
    .B2(\datamem.data_ram[4][27] ),
    .C1(_07419_),
    .X(_07420_));
 sky130_fd_sc_hd__o22a_1 _20128_ (.A1(\datamem.data_ram[11][27] ),
    .A2(_06828_),
    .B1(_06656_),
    .B2(\datamem.data_ram[9][27] ),
    .X(_07421_));
 sky130_fd_sc_hd__o221a_1 _20129_ (.A1(\datamem.data_ram[10][27] ),
    .A2(_06804_),
    .B1(_07037_),
    .B2(\datamem.data_ram[13][27] ),
    .C1(_07421_),
    .X(_07422_));
 sky130_fd_sc_hd__o22a_1 _20130_ (.A1(\datamem.data_ram[8][27] ),
    .A2(_06696_),
    .B1(_06686_),
    .B2(\datamem.data_ram[12][27] ),
    .X(_07423_));
 sky130_fd_sc_hd__o221a_1 _20131_ (.A1(\datamem.data_ram[14][27] ),
    .A2(_06682_),
    .B1(_06671_),
    .B2(\datamem.data_ram[15][27] ),
    .C1(_07423_),
    .X(_07424_));
 sky130_fd_sc_hd__and3_1 _20132_ (.A(_06602_),
    .B(_07422_),
    .C(_07424_),
    .X(_07425_));
 sky130_fd_sc_hd__a31o_1 _20133_ (.A1(_06777_),
    .A2(_07418_),
    .A3(_07420_),
    .B1(_07425_),
    .X(_07426_));
 sky130_fd_sc_hd__o22a_1 _20134_ (.A1(\datamem.data_ram[34][27] ),
    .A2(_06610_),
    .B1(_06805_),
    .B2(\datamem.data_ram[36][27] ),
    .X(_07427_));
 sky130_fd_sc_hd__o22a_1 _20135_ (.A1(\datamem.data_ram[38][27] ),
    .A2(_06626_),
    .B1(_06820_),
    .B2(\datamem.data_ram[32][27] ),
    .X(_07428_));
 sky130_fd_sc_hd__o221a_1 _20136_ (.A1(\datamem.data_ram[35][27] ),
    .A2(_06632_),
    .B1(_06704_),
    .B2(\datamem.data_ram[39][27] ),
    .C1(_06677_),
    .X(_07429_));
 sky130_fd_sc_hd__o211a_1 _20137_ (.A1(\datamem.data_ram[37][27] ),
    .A2(_06815_),
    .B1(_07428_),
    .C1(_07429_),
    .X(_07430_));
 sky130_fd_sc_hd__o211a_1 _20138_ (.A1(\datamem.data_ram[33][27] ),
    .A2(_06782_),
    .B1(_07427_),
    .C1(_07430_),
    .X(_07431_));
 sky130_fd_sc_hd__o22a_1 _20139_ (.A1(\datamem.data_ram[46][27] ),
    .A2(_06627_),
    .B1(_06821_),
    .B2(\datamem.data_ram[40][27] ),
    .X(_07432_));
 sky130_fd_sc_hd__o22a_1 _20140_ (.A1(\datamem.data_ram[45][27] ),
    .A2(_06721_),
    .B1(_06654_),
    .B2(\datamem.data_ram[41][27] ),
    .X(_07433_));
 sky130_fd_sc_hd__o221a_1 _20141_ (.A1(\datamem.data_ram[47][27] ),
    .A2(_06704_),
    .B1(_06617_),
    .B2(\datamem.data_ram[44][27] ),
    .C1(_07433_),
    .X(_07434_));
 sky130_fd_sc_hd__o211a_1 _20142_ (.A1(\datamem.data_ram[43][27] ),
    .A2(_06828_),
    .B1(_07434_),
    .C1(_06851_),
    .X(_07435_));
 sky130_fd_sc_hd__o211a_1 _20143_ (.A1(\datamem.data_ram[42][27] ),
    .A2(_06611_),
    .B1(_07432_),
    .C1(_07435_),
    .X(_07436_));
 sky130_fd_sc_hd__or3_2 _20144_ (.A(_06714_),
    .B(_07431_),
    .C(_07436_),
    .X(_07437_));
 sky130_fd_sc_hd__o22a_1 _20145_ (.A1(\datamem.data_ram[61][27] ),
    .A2(_06815_),
    .B1(_06781_),
    .B2(\datamem.data_ram[57][27] ),
    .X(_07438_));
 sky130_fd_sc_hd__o22a_1 _20146_ (.A1(\datamem.data_ram[59][27] ),
    .A2(_06729_),
    .B1(_06668_),
    .B2(\datamem.data_ram[63][27] ),
    .X(_07439_));
 sky130_fd_sc_hd__o221a_1 _20147_ (.A1(\datamem.data_ram[56][27] ),
    .A2(_06820_),
    .B1(_06617_),
    .B2(\datamem.data_ram[60][27] ),
    .C1(_07439_),
    .X(_07440_));
 sky130_fd_sc_hd__o211a_1 _20148_ (.A1(\datamem.data_ram[62][27] ),
    .A2(_06627_),
    .B1(_06600_),
    .C1(_07440_),
    .X(_07441_));
 sky130_fd_sc_hd__o211a_1 _20149_ (.A1(\datamem.data_ram[58][27] ),
    .A2(_06611_),
    .B1(_07438_),
    .C1(_07441_),
    .X(_07442_));
 sky130_fd_sc_hd__o22a_1 _20150_ (.A1(\datamem.data_ram[53][27] ),
    .A2(_06815_),
    .B1(_06670_),
    .B2(\datamem.data_ram[55][27] ),
    .X(_07443_));
 sky130_fd_sc_hd__o22a_1 _20151_ (.A1(\datamem.data_ram[54][27] ),
    .A2(_06626_),
    .B1(_06811_),
    .B2(\datamem.data_ram[48][27] ),
    .X(_07444_));
 sky130_fd_sc_hd__o221a_1 _20152_ (.A1(\datamem.data_ram[50][27] ),
    .A2(_06609_),
    .B1(_06632_),
    .B2(\datamem.data_ram[51][27] ),
    .C1(_06677_),
    .X(_07445_));
 sky130_fd_sc_hd__o211a_1 _20153_ (.A1(\datamem.data_ram[49][27] ),
    .A2(_06781_),
    .B1(_07444_),
    .C1(_07445_),
    .X(_07446_));
 sky130_fd_sc_hd__o211a_1 _20154_ (.A1(\datamem.data_ram[52][27] ),
    .A2(_07230_),
    .B1(_07443_),
    .C1(_07446_),
    .X(_07447_));
 sky130_fd_sc_hd__or3_1 _20155_ (.A(_06751_),
    .B(_07442_),
    .C(_07447_),
    .X(_07448_));
 sky130_fd_sc_hd__or2_1 _20156_ (.A(\datamem.data_ram[25][27] ),
    .B(_06657_),
    .X(_07449_));
 sky130_fd_sc_hd__o22a_1 _20157_ (.A1(\datamem.data_ram[31][27] ),
    .A2(_06671_),
    .B1(_06687_),
    .B2(\datamem.data_ram[28][27] ),
    .X(_07450_));
 sky130_fd_sc_hd__o22a_1 _20158_ (.A1(\datamem.data_ram[26][27] ),
    .A2(_06690_),
    .B1(_06730_),
    .B2(\datamem.data_ram[27][27] ),
    .X(_07451_));
 sky130_fd_sc_hd__o221a_1 _20159_ (.A1(\datamem.data_ram[30][27] ),
    .A2(_06718_),
    .B1(_06696_),
    .B2(\datamem.data_ram[24][27] ),
    .C1(_07451_),
    .X(_07452_));
 sky130_fd_sc_hd__o211a_1 _20160_ (.A1(\datamem.data_ram[29][27] ),
    .A2(_06724_),
    .B1(_06810_),
    .C1(_07452_),
    .X(_07453_));
 sky130_fd_sc_hd__o22a_1 _20161_ (.A1(\datamem.data_ram[18][27] ),
    .A2(_06728_),
    .B1(_06768_),
    .B2(\datamem.data_ram[21][27] ),
    .X(_07454_));
 sky130_fd_sc_hd__o22a_1 _20162_ (.A1(\datamem.data_ram[16][27] ),
    .A2(_06695_),
    .B1(_06725_),
    .B2(\datamem.data_ram[23][27] ),
    .X(_07455_));
 sky130_fd_sc_hd__o221a_1 _20163_ (.A1(\datamem.data_ram[19][27] ),
    .A2(_06730_),
    .B1(_06765_),
    .B2(\datamem.data_ram[20][27] ),
    .C1(_06732_),
    .X(_07456_));
 sky130_fd_sc_hd__o211a_1 _20164_ (.A1(\datamem.data_ram[22][27] ),
    .A2(_06718_),
    .B1(_07455_),
    .C1(_07456_),
    .X(_07457_));
 sky130_fd_sc_hd__o211a_1 _20165_ (.A1(\datamem.data_ram[17][27] ),
    .A2(_06657_),
    .B1(_07454_),
    .C1(_07457_),
    .X(_07458_));
 sky130_fd_sc_hd__a31o_1 _20166_ (.A1(_07449_),
    .A2(_07450_),
    .A3(_07453_),
    .B1(_07458_),
    .X(_07459_));
 sky130_fd_sc_hd__a32o_1 _20167_ (.A1(_06712_),
    .A2(_07437_),
    .A3(_07448_),
    .B1(_07459_),
    .B2(_06797_),
    .X(_07460_));
 sky130_fd_sc_hd__a21oi_4 _20168_ (.A1(_06596_),
    .A2(_07426_),
    .B1(_07460_),
    .Y(_07461_));
 sky130_fd_sc_hd__o22a_1 _20169_ (.A1(\datamem.data_ram[26][11] ),
    .A2(_06754_),
    .B1(_06697_),
    .B2(\datamem.data_ram[24][11] ),
    .X(_07462_));
 sky130_fd_sc_hd__o221a_1 _20170_ (.A1(\datamem.data_ram[28][11] ),
    .A2(_06688_),
    .B1(_06658_),
    .B2(\datamem.data_ram[25][11] ),
    .C1(_07462_),
    .X(_07463_));
 sky130_fd_sc_hd__o22a_1 _20171_ (.A1(\datamem.data_ram[30][11] ),
    .A2(_06764_),
    .B1(_06761_),
    .B2(\datamem.data_ram[31][11] ),
    .X(_07464_));
 sky130_fd_sc_hd__o221a_1 _20172_ (.A1(\datamem.data_ram[29][11] ),
    .A2(_06865_),
    .B1(_06863_),
    .B2(\datamem.data_ram[27][11] ),
    .C1(_07464_),
    .X(_07465_));
 sky130_fd_sc_hd__o22a_1 _20173_ (.A1(\datamem.data_ram[19][11] ),
    .A2(_06731_),
    .B1(_06656_),
    .B2(\datamem.data_ram[17][11] ),
    .X(_07466_));
 sky130_fd_sc_hd__o221a_1 _20174_ (.A1(\datamem.data_ram[16][11] ),
    .A2(_06837_),
    .B1(_06687_),
    .B2(\datamem.data_ram[20][11] ),
    .C1(_07466_),
    .X(_07467_));
 sky130_fd_sc_hd__o22a_1 _20175_ (.A1(\datamem.data_ram[21][11] ),
    .A2(_06768_),
    .B1(_06726_),
    .B2(\datamem.data_ram[23][11] ),
    .X(_07468_));
 sky130_fd_sc_hd__o221a_1 _20176_ (.A1(\datamem.data_ram[22][11] ),
    .A2(_06719_),
    .B1(_06754_),
    .B2(\datamem.data_ram[18][11] ),
    .C1(_07468_),
    .X(_07469_));
 sky130_fd_sc_hd__and3_1 _20177_ (.A(_06680_),
    .B(_07467_),
    .C(_07469_),
    .X(_07470_));
 sky130_fd_sc_hd__a31o_1 _20178_ (.A1(_06603_),
    .A2(_07463_),
    .A3(_07465_),
    .B1(_07470_),
    .X(_07471_));
 sky130_fd_sc_hd__o22a_1 _20179_ (.A1(\datamem.data_ram[15][11] ),
    .A2(_06761_),
    .B1(_07024_),
    .B2(\datamem.data_ram[12][11] ),
    .X(_07472_));
 sky130_fd_sc_hd__o22a_1 _20180_ (.A1(\datamem.data_ram[13][11] ),
    .A2(_06702_),
    .B1(_06778_),
    .B2(\datamem.data_ram[8][11] ),
    .X(_07473_));
 sky130_fd_sc_hd__o221a_1 _20181_ (.A1(\datamem.data_ram[14][11] ),
    .A2(_06763_),
    .B1(_06737_),
    .B2(\datamem.data_ram[11][11] ),
    .C1(_06741_),
    .X(_07474_));
 sky130_fd_sc_hd__o211a_1 _20182_ (.A1(\datamem.data_ram[10][11] ),
    .A2(_06692_),
    .B1(_07473_),
    .C1(_07474_),
    .X(_07475_));
 sky130_fd_sc_hd__o211a_1 _20183_ (.A1(\datamem.data_ram[9][11] ),
    .A2(_06701_),
    .B1(_07472_),
    .C1(_07475_),
    .X(_07476_));
 sky130_fd_sc_hd__o22a_1 _20184_ (.A1(\datamem.data_ram[0][11] ),
    .A2(_06779_),
    .B1(_06620_),
    .B2(\datamem.data_ram[4][11] ),
    .X(_07477_));
 sky130_fd_sc_hd__o22a_1 _20185_ (.A1(\datamem.data_ram[6][11] ),
    .A2(_07085_),
    .B1(_07243_),
    .B2(\datamem.data_ram[1][11] ),
    .X(_07478_));
 sky130_fd_sc_hd__o221a_1 _20186_ (.A1(\datamem.data_ram[5][11] ),
    .A2(_06768_),
    .B1(_06760_),
    .B2(\datamem.data_ram[7][11] ),
    .C1(_07478_),
    .X(_07479_));
 sky130_fd_sc_hd__o211a_1 _20187_ (.A1(\datamem.data_ram[2][11] ),
    .A2(_06692_),
    .B1(_07031_),
    .C1(_07479_),
    .X(_07480_));
 sky130_fd_sc_hd__o211a_1 _20188_ (.A1(\datamem.data_ram[3][11] ),
    .A2(_06739_),
    .B1(_07477_),
    .C1(_07480_),
    .X(_07481_));
 sky130_fd_sc_hd__o21a_1 _20189_ (.A1(_07476_),
    .A2(_07481_),
    .B1(_06596_),
    .X(_07482_));
 sky130_fd_sc_hd__o22a_1 _20190_ (.A1(\datamem.data_ram[40][11] ),
    .A2(_06697_),
    .B1(_07024_),
    .B2(\datamem.data_ram[44][11] ),
    .X(_07483_));
 sky130_fd_sc_hd__o22a_1 _20191_ (.A1(\datamem.data_ram[46][11] ),
    .A2(_06717_),
    .B1(_06730_),
    .B2(\datamem.data_ram[43][11] ),
    .X(_07484_));
 sky130_fd_sc_hd__o221a_1 _20192_ (.A1(\datamem.data_ram[42][11] ),
    .A2(_06728_),
    .B1(_06656_),
    .B2(\datamem.data_ram[41][11] ),
    .C1(_07484_),
    .X(_07485_));
 sky130_fd_sc_hd__o211a_1 _20193_ (.A1(\datamem.data_ram[47][11] ),
    .A2(_06761_),
    .B1(_07485_),
    .C1(_06742_),
    .X(_07486_));
 sky130_fd_sc_hd__o211a_1 _20194_ (.A1(\datamem.data_ram[45][11] ),
    .A2(_06865_),
    .B1(_07483_),
    .C1(_07486_),
    .X(_07487_));
 sky130_fd_sc_hd__o22a_1 _20195_ (.A1(\datamem.data_ram[38][11] ),
    .A2(_06764_),
    .B1(_07024_),
    .B2(\datamem.data_ram[36][11] ),
    .X(_07488_));
 sky130_fd_sc_hd__o22a_1 _20196_ (.A1(\datamem.data_ram[39][11] ),
    .A2(_06760_),
    .B1(_06699_),
    .B2(\datamem.data_ram[33][11] ),
    .X(_07489_));
 sky130_fd_sc_hd__o221a_1 _20197_ (.A1(\datamem.data_ram[32][11] ),
    .A2(_06778_),
    .B1(_06737_),
    .B2(\datamem.data_ram[35][11] ),
    .C1(_06769_),
    .X(_07490_));
 sky130_fd_sc_hd__o211a_1 _20198_ (.A1(\datamem.data_ram[37][11] ),
    .A2(_06703_),
    .B1(_07489_),
    .C1(_07490_),
    .X(_07491_));
 sky130_fd_sc_hd__o211a_1 _20199_ (.A1(\datamem.data_ram[34][11] ),
    .A2(_07023_),
    .B1(_07488_),
    .C1(_07491_),
    .X(_07492_));
 sky130_fd_sc_hd__o22a_1 _20200_ (.A1(\datamem.data_ram[62][11] ),
    .A2(_06763_),
    .B1(_06702_),
    .B2(\datamem.data_ram[61][11] ),
    .X(_07493_));
 sky130_fd_sc_hd__o22a_1 _20201_ (.A1(\datamem.data_ram[59][11] ),
    .A2(_06730_),
    .B1(_06765_),
    .B2(\datamem.data_ram[60][11] ),
    .X(_07494_));
 sky130_fd_sc_hd__o221a_1 _20202_ (.A1(\datamem.data_ram[58][11] ),
    .A2(_06690_),
    .B1(_07243_),
    .B2(\datamem.data_ram[57][11] ),
    .C1(_06600_),
    .X(_07495_));
 sky130_fd_sc_hd__o211a_1 _20203_ (.A1(\datamem.data_ram[56][11] ),
    .A2(_06778_),
    .B1(_07494_),
    .C1(_07495_),
    .X(_07496_));
 sky130_fd_sc_hd__o211a_1 _20204_ (.A1(\datamem.data_ram[63][11] ),
    .A2(_06761_),
    .B1(_07493_),
    .C1(_07496_),
    .X(_07497_));
 sky130_fd_sc_hd__o22a_1 _20205_ (.A1(\datamem.data_ram[50][11] ),
    .A2(_06691_),
    .B1(_06760_),
    .B2(\datamem.data_ram[55][11] ),
    .X(_07498_));
 sky130_fd_sc_hd__o22a_1 _20206_ (.A1(\datamem.data_ram[54][11] ),
    .A2(_06743_),
    .B1(_07242_),
    .B2(\datamem.data_ram[49][11] ),
    .X(_07499_));
 sky130_fd_sc_hd__o221a_1 _20207_ (.A1(\datamem.data_ram[53][11] ),
    .A2(_06722_),
    .B1(_06695_),
    .B2(\datamem.data_ram[48][11] ),
    .C1(_07499_),
    .X(_07500_));
 sky130_fd_sc_hd__o211a_1 _20208_ (.A1(\datamem.data_ram[52][11] ),
    .A2(_06766_),
    .B1(_07500_),
    .C1(_06769_),
    .X(_07501_));
 sky130_fd_sc_hd__o211a_1 _20209_ (.A1(\datamem.data_ram[51][11] ),
    .A2(_06738_),
    .B1(_07498_),
    .C1(_07501_),
    .X(_07502_));
 sky130_fd_sc_hd__o31a_1 _20210_ (.A1(_06752_),
    .A2(_07497_),
    .A3(_07502_),
    .B1(_06712_),
    .X(_07503_));
 sky130_fd_sc_hd__o31a_1 _20211_ (.A1(_06716_),
    .A2(_07487_),
    .A3(_07492_),
    .B1(_07503_),
    .X(_07504_));
 sky130_fd_sc_hd__a211oi_1 _20212_ (.A1(_06797_),
    .A2(_07471_),
    .B1(_07482_),
    .C1(_07504_),
    .Y(_07505_));
 sky130_fd_sc_hd__o32a_1 _20213_ (.A1(_05391_),
    .A2(_06586_),
    .A3(_07461_),
    .B1(net37),
    .B2(_07120_),
    .X(_07506_));
 sky130_fd_sc_hd__nor2_1 _20214_ (.A(_06590_),
    .B(_07506_),
    .Y(_07507_));
 sky130_fd_sc_hd__a22o_1 _20215_ (.A1(\datamem.data_ram[30][3] ),
    .A2(_07127_),
    .B1(_06977_),
    .B2(\datamem.data_ram[28][3] ),
    .X(_07508_));
 sky130_fd_sc_hd__a22o_1 _20216_ (.A1(\datamem.data_ram[27][3] ),
    .A2(_06941_),
    .B1(_06925_),
    .B2(\datamem.data_ram[31][3] ),
    .X(_07509_));
 sky130_fd_sc_hd__a221o_1 _20217_ (.A1(\datamem.data_ram[29][3] ),
    .A2(_06920_),
    .B1(_06937_),
    .B2(\datamem.data_ram[24][3] ),
    .C1(_07509_),
    .X(_07510_));
 sky130_fd_sc_hd__a211o_1 _20218_ (.A1(\datamem.data_ram[25][3] ),
    .A2(_06949_),
    .B1(_07510_),
    .C1(_06680_),
    .X(_07511_));
 sky130_fd_sc_hd__a211o_1 _20219_ (.A1(\datamem.data_ram[26][3] ),
    .A2(_07136_),
    .B1(_07508_),
    .C1(_07511_),
    .X(_07512_));
 sky130_fd_sc_hd__a22o_1 _20220_ (.A1(\datamem.data_ram[22][3] ),
    .A2(_07127_),
    .B1(_06976_),
    .B2(\datamem.data_ram[20][3] ),
    .X(_07513_));
 sky130_fd_sc_hd__a22o_1 _20221_ (.A1(\datamem.data_ram[19][3] ),
    .A2(_06961_),
    .B1(_06948_),
    .B2(\datamem.data_ram[17][3] ),
    .X(_07514_));
 sky130_fd_sc_hd__a221o_1 _20222_ (.A1(\datamem.data_ram[18][3] ),
    .A2(_06931_),
    .B1(_06926_),
    .B2(\datamem.data_ram[23][3] ),
    .C1(_06742_),
    .X(_07515_));
 sky130_fd_sc_hd__a211o_1 _20223_ (.A1(\datamem.data_ram[16][3] ),
    .A2(_07138_),
    .B1(_07514_),
    .C1(_07515_),
    .X(_07516_));
 sky130_fd_sc_hd__a211o_1 _20224_ (.A1(\datamem.data_ram[21][3] ),
    .A2(_07132_),
    .B1(_07513_),
    .C1(_07516_),
    .X(_07517_));
 sky130_fd_sc_hd__a22o_1 _20225_ (.A1(\datamem.data_ram[10][3] ),
    .A2(_06932_),
    .B1(_06955_),
    .B2(\datamem.data_ram[12][3] ),
    .X(_07518_));
 sky130_fd_sc_hd__a22o_1 _20226_ (.A1(\datamem.data_ram[8][3] ),
    .A2(_06935_),
    .B1(_06946_),
    .B2(\datamem.data_ram[9][3] ),
    .X(_07519_));
 sky130_fd_sc_hd__a221o_1 _20227_ (.A1(\datamem.data_ram[13][3] ),
    .A2(_06919_),
    .B1(_06925_),
    .B2(\datamem.data_ram[15][3] ),
    .C1(_07519_),
    .X(_07520_));
 sky130_fd_sc_hd__a211o_1 _20228_ (.A1(\datamem.data_ram[11][3] ),
    .A2(_06943_),
    .B1(_07520_),
    .C1(_07031_),
    .X(_07521_));
 sky130_fd_sc_hd__a211o_1 _20229_ (.A1(\datamem.data_ram[14][3] ),
    .A2(_07127_),
    .B1(_07518_),
    .C1(_07521_),
    .X(_07522_));
 sky130_fd_sc_hd__a22o_1 _20230_ (.A1(\datamem.data_ram[3][3] ),
    .A2(_06961_),
    .B1(_06955_),
    .B2(\datamem.data_ram[4][3] ),
    .X(_07523_));
 sky130_fd_sc_hd__a22o_1 _20231_ (.A1(\datamem.data_ram[7][3] ),
    .A2(_06925_),
    .B1(_06947_),
    .B2(\datamem.data_ram[1][3] ),
    .X(_07524_));
 sky130_fd_sc_hd__a221o_1 _20232_ (.A1(\datamem.data_ram[5][3] ),
    .A2(_06919_),
    .B1(_06936_),
    .B2(\datamem.data_ram[0][3] ),
    .C1(_06741_),
    .X(_07525_));
 sky130_fd_sc_hd__a211o_1 _20233_ (.A1(\datamem.data_ram[6][3] ),
    .A2(_06952_),
    .B1(_07524_),
    .C1(_07525_),
    .X(_07526_));
 sky130_fd_sc_hd__a211o_1 _20234_ (.A1(\datamem.data_ram[2][3] ),
    .A2(_07000_),
    .B1(_07523_),
    .C1(_07526_),
    .X(_07527_));
 sky130_fd_sc_hd__a31o_1 _20235_ (.A1(_06753_),
    .A2(_07522_),
    .A3(_07527_),
    .B1(_06713_),
    .X(_07528_));
 sky130_fd_sc_hd__a31o_1 _20236_ (.A1(_07071_),
    .A2(_07512_),
    .A3(_07517_),
    .B1(_07528_),
    .X(_07529_));
 sky130_fd_sc_hd__a22o_1 _20237_ (.A1(\datamem.data_ram[54][3] ),
    .A2(_07127_),
    .B1(_06966_),
    .B2(\datamem.data_ram[51][3] ),
    .X(_07530_));
 sky130_fd_sc_hd__a22o_1 _20238_ (.A1(\datamem.data_ram[52][3] ),
    .A2(_06954_),
    .B1(_06947_),
    .B2(\datamem.data_ram[49][3] ),
    .X(_07531_));
 sky130_fd_sc_hd__a221o_1 _20239_ (.A1(\datamem.data_ram[53][3] ),
    .A2(_06920_),
    .B1(_06937_),
    .B2(\datamem.data_ram[48][3] ),
    .C1(_07531_),
    .X(_07532_));
 sky130_fd_sc_hd__a211o_1 _20240_ (.A1(\datamem.data_ram[55][3] ),
    .A2(_06927_),
    .B1(_07532_),
    .C1(_06967_),
    .X(_07533_));
 sky130_fd_sc_hd__a211o_1 _20241_ (.A1(\datamem.data_ram[50][3] ),
    .A2(_07136_),
    .B1(_07530_),
    .C1(_07533_),
    .X(_07534_));
 sky130_fd_sc_hd__a22o_1 _20242_ (.A1(\datamem.data_ram[62][3] ),
    .A2(_07127_),
    .B1(_06976_),
    .B2(\datamem.data_ram[60][3] ),
    .X(_07535_));
 sky130_fd_sc_hd__a22o_1 _20243_ (.A1(\datamem.data_ram[56][3] ),
    .A2(_06937_),
    .B1(_06926_),
    .B2(\datamem.data_ram[63][3] ),
    .X(_07536_));
 sky130_fd_sc_hd__a22o_1 _20244_ (.A1(\datamem.data_ram[59][3] ),
    .A2(_06961_),
    .B1(_06948_),
    .B2(\datamem.data_ram[57][3] ),
    .X(_07537_));
 sky130_fd_sc_hd__a2111o_1 _20245_ (.A1(\datamem.data_ram[61][3] ),
    .A2(_06921_),
    .B1(_06680_),
    .C1(_07536_),
    .D1(_07537_),
    .X(_07538_));
 sky130_fd_sc_hd__a211o_1 _20246_ (.A1(\datamem.data_ram[58][3] ),
    .A2(_07136_),
    .B1(_07535_),
    .C1(_07538_),
    .X(_07539_));
 sky130_fd_sc_hd__a22o_1 _20247_ (.A1(\datamem.data_ram[34][3] ),
    .A2(_06931_),
    .B1(_06924_),
    .B2(\datamem.data_ram[39][3] ),
    .X(_07540_));
 sky130_fd_sc_hd__a221o_1 _20248_ (.A1(\datamem.data_ram[38][3] ),
    .A2(_06952_),
    .B1(_06958_),
    .B2(\datamem.data_ram[33][3] ),
    .C1(_07540_),
    .X(_07541_));
 sky130_fd_sc_hd__a22o_1 _20249_ (.A1(\datamem.data_ram[37][3] ),
    .A2(_06919_),
    .B1(_06954_),
    .B2(\datamem.data_ram[36][3] ),
    .X(_07542_));
 sky130_fd_sc_hd__a221o_1 _20250_ (.A1(\datamem.data_ram[32][3] ),
    .A2(_06937_),
    .B1(_06961_),
    .B2(\datamem.data_ram[35][3] ),
    .C1(_07542_),
    .X(_07543_));
 sky130_fd_sc_hd__or3_1 _20251_ (.A(_06967_),
    .B(_07541_),
    .C(_07543_),
    .X(_07544_));
 sky130_fd_sc_hd__a22o_1 _20252_ (.A1(\datamem.data_ram[46][3] ),
    .A2(_06951_),
    .B1(_06954_),
    .B2(\datamem.data_ram[44][3] ),
    .X(_07545_));
 sky130_fd_sc_hd__a221o_1 _20253_ (.A1(\datamem.data_ram[40][3] ),
    .A2(_06937_),
    .B1(_06958_),
    .B2(\datamem.data_ram[41][3] ),
    .C1(_07545_),
    .X(_07546_));
 sky130_fd_sc_hd__a22o_1 _20254_ (.A1(\datamem.data_ram[42][3] ),
    .A2(_06931_),
    .B1(_06924_),
    .B2(\datamem.data_ram[47][3] ),
    .X(_07547_));
 sky130_fd_sc_hd__a221o_1 _20255_ (.A1(\datamem.data_ram[45][3] ),
    .A2(_06920_),
    .B1(_06961_),
    .B2(\datamem.data_ram[43][3] ),
    .C1(_07547_),
    .X(_07548_));
 sky130_fd_sc_hd__or3_2 _20256_ (.A(_06680_),
    .B(_07546_),
    .C(_07548_),
    .X(_07549_));
 sky130_fd_sc_hd__a31o_1 _20257_ (.A1(_06753_),
    .A2(_07544_),
    .A3(_07549_),
    .B1(_06985_),
    .X(_07550_));
 sky130_fd_sc_hd__a31o_1 _20258_ (.A1(_07071_),
    .A2(_07534_),
    .A3(_07539_),
    .B1(_07550_),
    .X(_07551_));
 sky130_fd_sc_hd__and3_1 _20259_ (.A(_06988_),
    .B(_07529_),
    .C(_07551_),
    .X(_07552_));
 sky130_fd_sc_hd__o22a_1 _20260_ (.A1(\datamem.data_ram[51][19] ),
    .A2(_06635_),
    .B1(_06620_),
    .B2(\datamem.data_ram[52][19] ),
    .X(_07553_));
 sky130_fd_sc_hd__o221a_1 _20261_ (.A1(\datamem.data_ram[54][19] ),
    .A2(_06683_),
    .B1(_07023_),
    .B2(\datamem.data_ram[50][19] ),
    .C1(_07553_),
    .X(_07554_));
 sky130_fd_sc_hd__o22a_1 _20262_ (.A1(\datamem.data_ram[53][19] ),
    .A2(_06703_),
    .B1(_06707_),
    .B2(\datamem.data_ram[55][19] ),
    .X(_07555_));
 sky130_fd_sc_hd__o221a_1 _20263_ (.A1(\datamem.data_ram[48][19] ),
    .A2(_06698_),
    .B1(_06658_),
    .B2(\datamem.data_ram[49][19] ),
    .C1(_07555_),
    .X(_07556_));
 sky130_fd_sc_hd__o22a_1 _20264_ (.A1(\datamem.data_ram[63][19] ),
    .A2(_06760_),
    .B1(_06766_),
    .B2(\datamem.data_ram[60][19] ),
    .X(_07557_));
 sky130_fd_sc_hd__o221a_1 _20265_ (.A1(\datamem.data_ram[56][19] ),
    .A2(_06697_),
    .B1(_06657_),
    .B2(\datamem.data_ram[57][19] ),
    .C1(_07557_),
    .X(_07558_));
 sky130_fd_sc_hd__o22a_1 _20266_ (.A1(\datamem.data_ram[58][19] ),
    .A2(_06691_),
    .B1(_06768_),
    .B2(\datamem.data_ram[61][19] ),
    .X(_07559_));
 sky130_fd_sc_hd__o221a_1 _20267_ (.A1(\datamem.data_ram[62][19] ),
    .A2(_06719_),
    .B1(_06738_),
    .B2(\datamem.data_ram[59][19] ),
    .C1(_07559_),
    .X(_07560_));
 sky130_fd_sc_hd__and3_1 _20268_ (.A(_06967_),
    .B(_07558_),
    .C(_07560_),
    .X(_07561_));
 sky130_fd_sc_hd__a31o_1 _20269_ (.A1(_06681_),
    .A2(_07554_),
    .A3(_07556_),
    .B1(_07561_),
    .X(_07562_));
 sky130_fd_sc_hd__o22a_1 _20270_ (.A1(\datamem.data_ram[38][19] ),
    .A2(_06764_),
    .B1(_07024_),
    .B2(\datamem.data_ram[36][19] ),
    .X(_07563_));
 sky130_fd_sc_hd__o22a_1 _20271_ (.A1(\datamem.data_ram[39][19] ),
    .A2(_06760_),
    .B1(_06699_),
    .B2(\datamem.data_ram[33][19] ),
    .X(_07564_));
 sky130_fd_sc_hd__o221a_1 _20272_ (.A1(\datamem.data_ram[34][19] ),
    .A2(_06728_),
    .B1(_06737_),
    .B2(\datamem.data_ram[35][19] ),
    .C1(_06733_),
    .X(_07565_));
 sky130_fd_sc_hd__o211a_1 _20273_ (.A1(\datamem.data_ram[37][19] ),
    .A2(_06724_),
    .B1(_07564_),
    .C1(_07565_),
    .X(_07566_));
 sky130_fd_sc_hd__o211a_1 _20274_ (.A1(\datamem.data_ram[32][19] ),
    .A2(_06698_),
    .B1(_07563_),
    .C1(_07566_),
    .X(_07567_));
 sky130_fd_sc_hd__o22a_1 _20275_ (.A1(\datamem.data_ram[46][19] ),
    .A2(_06764_),
    .B1(_06700_),
    .B2(\datamem.data_ram[41][19] ),
    .X(_07568_));
 sky130_fd_sc_hd__o22a_1 _20276_ (.A1(\datamem.data_ram[47][19] ),
    .A2(_06725_),
    .B1(_06765_),
    .B2(\datamem.data_ram[44][19] ),
    .X(_07569_));
 sky130_fd_sc_hd__o221a_1 _20277_ (.A1(\datamem.data_ram[45][19] ),
    .A2(_06768_),
    .B1(_06696_),
    .B2(\datamem.data_ram[40][19] ),
    .C1(_07569_),
    .X(_07570_));
 sky130_fd_sc_hd__o211a_1 _20278_ (.A1(\datamem.data_ram[43][19] ),
    .A2(_06738_),
    .B1(_07570_),
    .C1(_06742_),
    .X(_07571_));
 sky130_fd_sc_hd__o211a_1 _20279_ (.A1(\datamem.data_ram[42][19] ),
    .A2(_07023_),
    .B1(_07568_),
    .C1(_07571_),
    .X(_07572_));
 sky130_fd_sc_hd__or3_1 _20280_ (.A(_06716_),
    .B(_07567_),
    .C(_07572_),
    .X(_07573_));
 sky130_fd_sc_hd__o211a_1 _20281_ (.A1(_06916_),
    .A2(_07562_),
    .B1(_07573_),
    .C1(_06713_),
    .X(_07574_));
 sky130_fd_sc_hd__o22a_1 _20282_ (.A1(\datamem.data_ram[29][19] ),
    .A2(_06865_),
    .B1(_06672_),
    .B2(\datamem.data_ram[31][19] ),
    .X(_07575_));
 sky130_fd_sc_hd__o22a_1 _20283_ (.A1(\datamem.data_ram[30][19] ),
    .A2(_06763_),
    .B1(_06699_),
    .B2(\datamem.data_ram[25][19] ),
    .X(_07576_));
 sky130_fd_sc_hd__o221a_1 _20284_ (.A1(\datamem.data_ram[24][19] ),
    .A2(_06697_),
    .B1(_07024_),
    .B2(\datamem.data_ram[28][19] ),
    .C1(_07576_),
    .X(_07577_));
 sky130_fd_sc_hd__o211a_1 _20285_ (.A1(\datamem.data_ram[27][19] ),
    .A2(_06739_),
    .B1(_07577_),
    .C1(_06967_),
    .X(_07578_));
 sky130_fd_sc_hd__o211a_1 _20286_ (.A1(\datamem.data_ram[26][19] ),
    .A2(_06613_),
    .B1(_07575_),
    .C1(_07578_),
    .X(_07579_));
 sky130_fd_sc_hd__o22a_1 _20287_ (.A1(\datamem.data_ram[21][19] ),
    .A2(_06865_),
    .B1(_06672_),
    .B2(\datamem.data_ram[23][19] ),
    .X(_07580_));
 sky130_fd_sc_hd__o22a_1 _20288_ (.A1(\datamem.data_ram[22][19] ),
    .A2(_06629_),
    .B1(_06779_),
    .B2(\datamem.data_ram[16][19] ),
    .X(_07581_));
 sky130_fd_sc_hd__o221a_1 _20289_ (.A1(\datamem.data_ram[18][19] ),
    .A2(_06692_),
    .B1(_06635_),
    .B2(\datamem.data_ram[19][19] ),
    .C1(_07031_),
    .X(_07582_));
 sky130_fd_sc_hd__o211a_1 _20290_ (.A1(\datamem.data_ram[20][19] ),
    .A2(_06688_),
    .B1(_07581_),
    .C1(_07582_),
    .X(_07583_));
 sky130_fd_sc_hd__o211a_1 _20291_ (.A1(\datamem.data_ram[17][19] ),
    .A2(_06659_),
    .B1(_07580_),
    .C1(_07583_),
    .X(_07584_));
 sky130_fd_sc_hd__o22a_1 _20292_ (.A1(\datamem.data_ram[14][19] ),
    .A2(_06764_),
    .B1(_06700_),
    .B2(\datamem.data_ram[9][19] ),
    .X(_07585_));
 sky130_fd_sc_hd__o22a_1 _20293_ (.A1(\datamem.data_ram[13][19] ),
    .A2(_06662_),
    .B1(_06646_),
    .B2(\datamem.data_ram[8][19] ),
    .X(_07586_));
 sky130_fd_sc_hd__o221a_1 _20294_ (.A1(\datamem.data_ram[15][19] ),
    .A2(_06726_),
    .B1(_06766_),
    .B2(\datamem.data_ram[12][19] ),
    .C1(_07586_),
    .X(_07587_));
 sky130_fd_sc_hd__o211a_1 _20295_ (.A1(\datamem.data_ram[10][19] ),
    .A2(_06754_),
    .B1(_06742_),
    .C1(_07587_),
    .X(_07588_));
 sky130_fd_sc_hd__o211a_1 _20296_ (.A1(\datamem.data_ram[11][19] ),
    .A2(_06739_),
    .B1(_07585_),
    .C1(_07588_),
    .X(_07589_));
 sky130_fd_sc_hd__o22a_1 _20297_ (.A1(\datamem.data_ram[6][19] ),
    .A2(_06764_),
    .B1(_07024_),
    .B2(\datamem.data_ram[4][19] ),
    .X(_07590_));
 sky130_fd_sc_hd__o22a_1 _20298_ (.A1(\datamem.data_ram[5][19] ),
    .A2(_06768_),
    .B1(_06699_),
    .B2(\datamem.data_ram[1][19] ),
    .X(_07591_));
 sky130_fd_sc_hd__o221a_1 _20299_ (.A1(\datamem.data_ram[2][19] ),
    .A2(_06691_),
    .B1(_06737_),
    .B2(\datamem.data_ram[3][19] ),
    .C1(_06769_),
    .X(_07592_));
 sky130_fd_sc_hd__o211a_1 _20300_ (.A1(\datamem.data_ram[7][19] ),
    .A2(_06761_),
    .B1(_07591_),
    .C1(_07592_),
    .X(_07593_));
 sky130_fd_sc_hd__o211a_1 _20301_ (.A1(\datamem.data_ram[0][19] ),
    .A2(_06698_),
    .B1(_07590_),
    .C1(_07593_),
    .X(_07594_));
 sky130_fd_sc_hd__or3_1 _20302_ (.A(_06716_),
    .B(_07589_),
    .C(_07594_),
    .X(_07595_));
 sky130_fd_sc_hd__o311a_1 _20303_ (.A1(_06916_),
    .A2(_07579_),
    .A3(_07584_),
    .B1(_07595_),
    .C1(_06985_),
    .X(_07596_));
 sky130_fd_sc_hd__nor2_2 _20304_ (.A(_07574_),
    .B(_07596_),
    .Y(_07597_));
 sky130_fd_sc_hd__nor2_1 _20305_ (.A(_07227_),
    .B(_07597_),
    .Y(_07598_));
 sky130_fd_sc_hd__or3_1 _20306_ (.A(_07507_),
    .B(_07552_),
    .C(_07598_),
    .X(_07599_));
 sky130_fd_sc_hd__clkbuf_1 _20307_ (.A(_07599_),
    .X(_04440_));
 sky130_fd_sc_hd__a22o_1 _20308_ (.A1(\datamem.data_ram[7][4] ),
    .A2(_06927_),
    .B1(_07133_),
    .B2(\datamem.data_ram[1][4] ),
    .X(_07600_));
 sky130_fd_sc_hd__a22o_1 _20309_ (.A1(\datamem.data_ram[2][4] ),
    .A2(_06932_),
    .B1(_06976_),
    .B2(\datamem.data_ram[4][4] ),
    .X(_07601_));
 sky130_fd_sc_hd__a22o_1 _20310_ (.A1(\datamem.data_ram[6][4] ),
    .A2(_06978_),
    .B1(_06943_),
    .B2(\datamem.data_ram[3][4] ),
    .X(_07602_));
 sky130_fd_sc_hd__a2111o_1 _20311_ (.A1(\datamem.data_ram[0][4] ),
    .A2(_07138_),
    .B1(_07601_),
    .C1(_07602_),
    .D1(_07081_),
    .X(_07603_));
 sky130_fd_sc_hd__a211o_1 _20312_ (.A1(\datamem.data_ram[5][4] ),
    .A2(_07132_),
    .B1(_07600_),
    .C1(_07603_),
    .X(_07604_));
 sky130_fd_sc_hd__a22o_1 _20313_ (.A1(\datamem.data_ram[10][4] ),
    .A2(_07000_),
    .B1(_07133_),
    .B2(\datamem.data_ram[9][4] ),
    .X(_07605_));
 sky130_fd_sc_hd__a22o_1 _20314_ (.A1(\datamem.data_ram[11][4] ),
    .A2(_06943_),
    .B1(_06993_),
    .B2(\datamem.data_ram[15][4] ),
    .X(_07606_));
 sky130_fd_sc_hd__a221o_1 _20315_ (.A1(\datamem.data_ram[13][4] ),
    .A2(_06969_),
    .B1(_06976_),
    .B2(\datamem.data_ram[12][4] ),
    .C1(_06776_),
    .X(_07607_));
 sky130_fd_sc_hd__a211o_1 _20316_ (.A1(\datamem.data_ram[8][4] ),
    .A2(_07138_),
    .B1(_07606_),
    .C1(_07607_),
    .X(_07608_));
 sky130_fd_sc_hd__a211o_1 _20317_ (.A1(\datamem.data_ram[14][4] ),
    .A2(_07159_),
    .B1(_07605_),
    .C1(_07608_),
    .X(_07609_));
 sky130_fd_sc_hd__and3_1 _20318_ (.A(_06916_),
    .B(_07604_),
    .C(_07609_),
    .X(_07610_));
 sky130_fd_sc_hd__a22o_1 _20319_ (.A1(\datamem.data_ram[24][4] ),
    .A2(_07122_),
    .B1(_07133_),
    .B2(\datamem.data_ram[25][4] ),
    .X(_07611_));
 sky130_fd_sc_hd__a22o_1 _20320_ (.A1(\datamem.data_ram[26][4] ),
    .A2(_06989_),
    .B1(_06921_),
    .B2(\datamem.data_ram[29][4] ),
    .X(_07612_));
 sky130_fd_sc_hd__a221o_1 _20321_ (.A1(\datamem.data_ram[27][4] ),
    .A2(_06943_),
    .B1(_06926_),
    .B2(\datamem.data_ram[31][4] ),
    .C1(_06776_),
    .X(_07613_));
 sky130_fd_sc_hd__a211o_1 _20322_ (.A1(\datamem.data_ram[30][4] ),
    .A2(_07159_),
    .B1(_07612_),
    .C1(_07613_),
    .X(_07614_));
 sky130_fd_sc_hd__a211o_1 _20323_ (.A1(\datamem.data_ram[28][4] ),
    .A2(_07123_),
    .B1(_07611_),
    .C1(_07614_),
    .X(_07615_));
 sky130_fd_sc_hd__a22o_1 _20324_ (.A1(\datamem.data_ram[18][4] ),
    .A2(_06989_),
    .B1(_06921_),
    .B2(\datamem.data_ram[21][4] ),
    .X(_07616_));
 sky130_fd_sc_hd__a211o_1 _20325_ (.A1(\datamem.data_ram[22][4] ),
    .A2(_07159_),
    .B1(_07081_),
    .C1(_07616_),
    .X(_07617_));
 sky130_fd_sc_hd__a22o_1 _20326_ (.A1(\datamem.data_ram[19][4] ),
    .A2(_06943_),
    .B1(_06993_),
    .B2(\datamem.data_ram[23][4] ),
    .X(_07618_));
 sky130_fd_sc_hd__a221o_1 _20327_ (.A1(\datamem.data_ram[16][4] ),
    .A2(_07138_),
    .B1(_06977_),
    .B2(\datamem.data_ram[20][4] ),
    .C1(_07618_),
    .X(_07619_));
 sky130_fd_sc_hd__a211o_1 _20328_ (.A1(\datamem.data_ram[17][4] ),
    .A2(_06997_),
    .B1(_07617_),
    .C1(_07619_),
    .X(_07620_));
 sky130_fd_sc_hd__a31o_1 _20329_ (.A1(_07071_),
    .A2(_07615_),
    .A3(_07620_),
    .B1(_06713_),
    .X(_07621_));
 sky130_fd_sc_hd__a22o_1 _20330_ (.A1(\datamem.data_ram[45][4] ),
    .A2(_06921_),
    .B1(_06993_),
    .B2(\datamem.data_ram[47][4] ),
    .X(_07622_));
 sky130_fd_sc_hd__a221o_1 _20331_ (.A1(\datamem.data_ram[46][4] ),
    .A2(_07159_),
    .B1(_06949_),
    .B2(\datamem.data_ram[41][4] ),
    .C1(_07622_),
    .X(_07623_));
 sky130_fd_sc_hd__a22o_1 _20332_ (.A1(\datamem.data_ram[42][4] ),
    .A2(_06989_),
    .B1(_06990_),
    .B2(\datamem.data_ram[40][4] ),
    .X(_07624_));
 sky130_fd_sc_hd__a221o_1 _20333_ (.A1(\datamem.data_ram[43][4] ),
    .A2(_06966_),
    .B1(_06977_),
    .B2(\datamem.data_ram[44][4] ),
    .C1(_07624_),
    .X(_07625_));
 sky130_fd_sc_hd__a22o_1 _20334_ (.A1(\datamem.data_ram[37][4] ),
    .A2(_06921_),
    .B1(_06993_),
    .B2(\datamem.data_ram[39][4] ),
    .X(_07626_));
 sky130_fd_sc_hd__a22o_1 _20335_ (.A1(\datamem.data_ram[34][4] ),
    .A2(_06930_),
    .B1(_06941_),
    .B2(\datamem.data_ram[35][4] ),
    .X(_07627_));
 sky130_fd_sc_hd__a221o_1 _20336_ (.A1(\datamem.data_ram[38][4] ),
    .A2(_06951_),
    .B1(_06954_),
    .B2(\datamem.data_ram[36][4] ),
    .C1(_07627_),
    .X(_07628_));
 sky130_fd_sc_hd__a211o_1 _20337_ (.A1(\datamem.data_ram[32][4] ),
    .A2(_06990_),
    .B1(_07628_),
    .C1(_06967_),
    .X(_07629_));
 sky130_fd_sc_hd__a211o_1 _20338_ (.A1(\datamem.data_ram[33][4] ),
    .A2(_07133_),
    .B1(_07626_),
    .C1(_07629_),
    .X(_07630_));
 sky130_fd_sc_hd__o31a_1 _20339_ (.A1(_07131_),
    .A2(_07623_),
    .A3(_07625_),
    .B1(_07630_),
    .X(_07631_));
 sky130_fd_sc_hd__a22o_1 _20340_ (.A1(\datamem.data_ram[58][4] ),
    .A2(_06989_),
    .B1(_06990_),
    .B2(\datamem.data_ram[56][4] ),
    .X(_07632_));
 sky130_fd_sc_hd__a221o_1 _20341_ (.A1(\datamem.data_ram[61][4] ),
    .A2(_06970_),
    .B1(_06977_),
    .B2(\datamem.data_ram[60][4] ),
    .C1(_07632_),
    .X(_07633_));
 sky130_fd_sc_hd__a22o_1 _20342_ (.A1(\datamem.data_ram[62][4] ),
    .A2(_06978_),
    .B1(_06948_),
    .B2(\datamem.data_ram[57][4] ),
    .X(_07634_));
 sky130_fd_sc_hd__clkbuf_8 _20343_ (.A(_06666_),
    .X(_07635_));
 sky130_fd_sc_hd__buf_6 _20344_ (.A(_06607_),
    .X(_07636_));
 sky130_fd_sc_hd__a31o_1 _20345_ (.A1(_07635_),
    .A2(\datamem.data_ram[59][4] ),
    .A3(_07636_),
    .B1(_06776_),
    .X(_07637_));
 sky130_fd_sc_hd__a211o_1 _20346_ (.A1(\datamem.data_ram[63][4] ),
    .A2(_07125_),
    .B1(_07634_),
    .C1(_07637_),
    .X(_07638_));
 sky130_fd_sc_hd__a22o_1 _20347_ (.A1(\datamem.data_ram[48][4] ),
    .A2(_06990_),
    .B1(_06976_),
    .B2(\datamem.data_ram[52][4] ),
    .X(_07639_));
 sky130_fd_sc_hd__a22o_1 _20348_ (.A1(\datamem.data_ram[51][4] ),
    .A2(_06942_),
    .B1(_06958_),
    .B2(\datamem.data_ram[49][4] ),
    .X(_07640_));
 sky130_fd_sc_hd__a221o_1 _20349_ (.A1(\datamem.data_ram[54][4] ),
    .A2(_06951_),
    .B1(_06931_),
    .B2(\datamem.data_ram[50][4] ),
    .C1(_06601_),
    .X(_07641_));
 sky130_fd_sc_hd__a211o_1 _20350_ (.A1(\datamem.data_ram[55][4] ),
    .A2(_06993_),
    .B1(_07640_),
    .C1(_07641_),
    .X(_07642_));
 sky130_fd_sc_hd__a211o_1 _20351_ (.A1(\datamem.data_ram[53][4] ),
    .A2(_06970_),
    .B1(_07639_),
    .C1(_07642_),
    .X(_07643_));
 sky130_fd_sc_hd__o211a_1 _20352_ (.A1(_07633_),
    .A2(_07638_),
    .B1(_07643_),
    .C1(_06716_),
    .X(_07644_));
 sky130_fd_sc_hd__a211o_1 _20353_ (.A1(_06916_),
    .A2(_07631_),
    .B1(_07644_),
    .C1(_06985_),
    .X(_07645_));
 sky130_fd_sc_hd__o21ai_2 _20354_ (.A1(_07610_),
    .A2(_07621_),
    .B1(_07645_),
    .Y(_07646_));
 sky130_fd_sc_hd__or2_1 _20355_ (.A(\datamem.data_ram[11][28] ),
    .B(_06738_),
    .X(_07647_));
 sky130_fd_sc_hd__o22a_1 _20356_ (.A1(\datamem.data_ram[14][28] ),
    .A2(_06764_),
    .B1(_06700_),
    .B2(\datamem.data_ram[9][28] ),
    .X(_07648_));
 sky130_fd_sc_hd__o22a_1 _20357_ (.A1(\datamem.data_ram[10][28] ),
    .A2(_06690_),
    .B1(_06725_),
    .B2(\datamem.data_ram[15][28] ),
    .X(_07649_));
 sky130_fd_sc_hd__o221a_1 _20358_ (.A1(\datamem.data_ram[8][28] ),
    .A2(_06696_),
    .B1(_06686_),
    .B2(\datamem.data_ram[12][28] ),
    .C1(_07649_),
    .X(_07650_));
 sky130_fd_sc_hd__o211a_1 _20359_ (.A1(\datamem.data_ram[13][28] ),
    .A2(_06724_),
    .B1(_06742_),
    .C1(_07650_),
    .X(_07651_));
 sky130_fd_sc_hd__o22a_1 _20360_ (.A1(\datamem.data_ram[6][28] ),
    .A2(_06763_),
    .B1(_06766_),
    .B2(\datamem.data_ram[4][28] ),
    .X(_07652_));
 sky130_fd_sc_hd__o22a_1 _20361_ (.A1(\datamem.data_ram[7][28] ),
    .A2(_06725_),
    .B1(_07243_),
    .B2(\datamem.data_ram[1][28] ),
    .X(_07653_));
 sky130_fd_sc_hd__o221a_1 _20362_ (.A1(\datamem.data_ram[0][28] ),
    .A2(_06695_),
    .B1(_06730_),
    .B2(\datamem.data_ram[3][28] ),
    .C1(_06678_),
    .X(_07654_));
 sky130_fd_sc_hd__o211a_1 _20363_ (.A1(\datamem.data_ram[5][28] ),
    .A2(_06702_),
    .B1(_07653_),
    .C1(_07654_),
    .X(_07655_));
 sky130_fd_sc_hd__o211a_1 _20364_ (.A1(\datamem.data_ram[2][28] ),
    .A2(_06692_),
    .B1(_07652_),
    .C1(_07655_),
    .X(_07656_));
 sky130_fd_sc_hd__a31o_1 _20365_ (.A1(_07647_),
    .A2(_07648_),
    .A3(_07651_),
    .B1(_07656_),
    .X(_07657_));
 sky130_fd_sc_hd__o22a_1 _20366_ (.A1(\datamem.data_ram[38][28] ),
    .A2(_06717_),
    .B1(_06685_),
    .B2(\datamem.data_ram[36][28] ),
    .X(_07658_));
 sky130_fd_sc_hd__o22a_1 _20367_ (.A1(\datamem.data_ram[39][28] ),
    .A2(_06668_),
    .B1(_06654_),
    .B2(\datamem.data_ram[33][28] ),
    .X(_07659_));
 sky130_fd_sc_hd__o221a_1 _20368_ (.A1(\datamem.data_ram[34][28] ),
    .A2(_06689_),
    .B1(_06729_),
    .B2(\datamem.data_ram[35][28] ),
    .C1(_06676_),
    .X(_07660_));
 sky130_fd_sc_hd__o211a_1 _20369_ (.A1(\datamem.data_ram[37][28] ),
    .A2(_06722_),
    .B1(_07659_),
    .C1(_07660_),
    .X(_07661_));
 sky130_fd_sc_hd__o211a_1 _20370_ (.A1(\datamem.data_ram[32][28] ),
    .A2(_06807_),
    .B1(_07658_),
    .C1(_07661_),
    .X(_07662_));
 sky130_fd_sc_hd__o22a_1 _20371_ (.A1(\datamem.data_ram[44][28] ),
    .A2(_06685_),
    .B1(_06655_),
    .B2(\datamem.data_ram[41][28] ),
    .X(_07663_));
 sky130_fd_sc_hd__o22a_1 _20372_ (.A1(\datamem.data_ram[42][28] ),
    .A2(_06608_),
    .B1(_06667_),
    .B2(\datamem.data_ram[47][28] ),
    .X(_07664_));
 sky130_fd_sc_hd__o221a_1 _20373_ (.A1(\datamem.data_ram[46][28] ),
    .A2(_06625_),
    .B1(_06645_),
    .B2(\datamem.data_ram[40][28] ),
    .C1(_07664_),
    .X(_07665_));
 sky130_fd_sc_hd__o211a_1 _20374_ (.A1(\datamem.data_ram[45][28] ),
    .A2(_06722_),
    .B1(_06599_),
    .C1(_07665_),
    .X(_07666_));
 sky130_fd_sc_hd__o211a_1 _20375_ (.A1(\datamem.data_ram[43][28] ),
    .A2(_06828_),
    .B1(_07663_),
    .C1(_07666_),
    .X(_07667_));
 sky130_fd_sc_hd__or3_2 _20376_ (.A(_06714_),
    .B(_07662_),
    .C(_07667_),
    .X(_07668_));
 sky130_fd_sc_hd__o22a_1 _20377_ (.A1(\datamem.data_ram[58][28] ),
    .A2(_06802_),
    .B1(_06695_),
    .B2(\datamem.data_ram[56][28] ),
    .X(_07669_));
 sky130_fd_sc_hd__o22a_1 _20378_ (.A1(\datamem.data_ram[61][28] ),
    .A2(_06660_),
    .B1(_06653_),
    .B2(\datamem.data_ram[57][28] ),
    .X(_07670_));
 sky130_fd_sc_hd__o221a_1 _20379_ (.A1(\datamem.data_ram[62][28] ),
    .A2(_06625_),
    .B1(_06684_),
    .B2(\datamem.data_ram[60][28] ),
    .C1(_07670_),
    .X(_07671_));
 sky130_fd_sc_hd__o211a_1 _20380_ (.A1(\datamem.data_ram[63][28] ),
    .A2(_06669_),
    .B1(_07671_),
    .C1(_06599_),
    .X(_07672_));
 sky130_fd_sc_hd__o211a_1 _20381_ (.A1(\datamem.data_ram[59][28] ),
    .A2(_06828_),
    .B1(_07669_),
    .C1(_07672_),
    .X(_07673_));
 sky130_fd_sc_hd__o22a_1 _20382_ (.A1(\datamem.data_ram[54][28] ),
    .A2(_06717_),
    .B1(_06695_),
    .B2(\datamem.data_ram[48][28] ),
    .X(_07674_));
 sky130_fd_sc_hd__o22a_1 _20383_ (.A1(\datamem.data_ram[53][28] ),
    .A2(_06721_),
    .B1(_07242_),
    .B2(\datamem.data_ram[49][28] ),
    .X(_07675_));
 sky130_fd_sc_hd__o221a_1 _20384_ (.A1(\datamem.data_ram[51][28] ),
    .A2(_06729_),
    .B1(_06668_),
    .B2(\datamem.data_ram[55][28] ),
    .C1(_06676_),
    .X(_07676_));
 sky130_fd_sc_hd__o211a_1 _20385_ (.A1(\datamem.data_ram[52][28] ),
    .A2(_06685_),
    .B1(_07675_),
    .C1(_07676_),
    .X(_07677_));
 sky130_fd_sc_hd__o211a_1 _20386_ (.A1(\datamem.data_ram[50][28] ),
    .A2(_06803_),
    .B1(_07674_),
    .C1(_07677_),
    .X(_07678_));
 sky130_fd_sc_hd__or3_1 _20387_ (.A(_06751_),
    .B(_07673_),
    .C(_07678_),
    .X(_07679_));
 sky130_fd_sc_hd__o22a_1 _20388_ (.A1(\datamem.data_ram[22][28] ),
    .A2(_06744_),
    .B1(_07243_),
    .B2(\datamem.data_ram[17][28] ),
    .X(_07680_));
 sky130_fd_sc_hd__o221a_1 _20389_ (.A1(\datamem.data_ram[21][28] ),
    .A2(_06768_),
    .B1(_06737_),
    .B2(\datamem.data_ram[19][28] ),
    .C1(_07680_),
    .X(_07681_));
 sky130_fd_sc_hd__o22a_1 _20390_ (.A1(\datamem.data_ram[16][28] ),
    .A2(_06646_),
    .B1(_06705_),
    .B2(\datamem.data_ram[23][28] ),
    .X(_07682_));
 sky130_fd_sc_hd__o221a_1 _20391_ (.A1(\datamem.data_ram[18][28] ),
    .A2(_06728_),
    .B1(_06766_),
    .B2(\datamem.data_ram[20][28] ),
    .C1(_07682_),
    .X(_07683_));
 sky130_fd_sc_hd__o22a_1 _20392_ (.A1(\datamem.data_ram[26][28] ),
    .A2(_06689_),
    .B1(_06661_),
    .B2(\datamem.data_ram[29][28] ),
    .X(_07684_));
 sky130_fd_sc_hd__o221a_1 _20393_ (.A1(\datamem.data_ram[31][28] ),
    .A2(_06725_),
    .B1(_06655_),
    .B2(\datamem.data_ram[25][28] ),
    .C1(_07684_),
    .X(_07685_));
 sky130_fd_sc_hd__o22a_1 _20394_ (.A1(\datamem.data_ram[30][28] ),
    .A2(_06625_),
    .B1(_06684_),
    .B2(\datamem.data_ram[28][28] ),
    .X(_07686_));
 sky130_fd_sc_hd__o221a_1 _20395_ (.A1(\datamem.data_ram[24][28] ),
    .A2(_06695_),
    .B1(_06730_),
    .B2(\datamem.data_ram[27][28] ),
    .C1(_07686_),
    .X(_07687_));
 sky130_fd_sc_hd__and3_1 _20396_ (.A(_06741_),
    .B(_07685_),
    .C(_07687_),
    .X(_07688_));
 sky130_fd_sc_hd__a31o_1 _20397_ (.A1(_07031_),
    .A2(_07681_),
    .A3(_07683_),
    .B1(_07688_),
    .X(_07689_));
 sky130_fd_sc_hd__a32o_1 _20398_ (.A1(_06712_),
    .A2(_07668_),
    .A3(_07679_),
    .B1(_07689_),
    .B2(_06796_),
    .X(_07690_));
 sky130_fd_sc_hd__a21oi_4 _20399_ (.A1(_06595_),
    .A2(_07657_),
    .B1(_07690_),
    .Y(_07691_));
 sky130_fd_sc_hd__or3_1 _20400_ (.A(_05391_),
    .B(_06586_),
    .C(_07691_),
    .X(_07692_));
 sky130_fd_sc_hd__o22a_1 _20401_ (.A1(\datamem.data_ram[37][12] ),
    .A2(_06815_),
    .B1(_06705_),
    .B2(\datamem.data_ram[39][12] ),
    .X(_07693_));
 sky130_fd_sc_hd__o221a_1 _20402_ (.A1(\datamem.data_ram[34][12] ),
    .A2(_06691_),
    .B1(_06778_),
    .B2(\datamem.data_ram[32][12] ),
    .C1(_07693_),
    .X(_07694_));
 sky130_fd_sc_hd__o22a_1 _20403_ (.A1(\datamem.data_ram[38][12] ),
    .A2(_07085_),
    .B1(_06618_),
    .B2(\datamem.data_ram[36][12] ),
    .X(_07695_));
 sky130_fd_sc_hd__o221a_1 _20404_ (.A1(\datamem.data_ram[35][12] ),
    .A2(_06737_),
    .B1(_06782_),
    .B2(\datamem.data_ram[33][12] ),
    .C1(_07695_),
    .X(_07696_));
 sky130_fd_sc_hd__o22a_1 _20405_ (.A1(\datamem.data_ram[40][12] ),
    .A2(_06820_),
    .B1(_06617_),
    .B2(\datamem.data_ram[44][12] ),
    .X(_07697_));
 sky130_fd_sc_hd__o221a_1 _20406_ (.A1(\datamem.data_ram[46][12] ),
    .A2(_06744_),
    .B1(_06690_),
    .B2(\datamem.data_ram[42][12] ),
    .C1(_07697_),
    .X(_07698_));
 sky130_fd_sc_hd__o22a_1 _20407_ (.A1(\datamem.data_ram[47][12] ),
    .A2(_06704_),
    .B1(_06780_),
    .B2(\datamem.data_ram[41][12] ),
    .X(_07699_));
 sky130_fd_sc_hd__o221a_1 _20408_ (.A1(\datamem.data_ram[45][12] ),
    .A2(_06662_),
    .B1(_06633_),
    .B2(\datamem.data_ram[43][12] ),
    .C1(_07699_),
    .X(_07700_));
 sky130_fd_sc_hd__and3_1 _20409_ (.A(_06601_),
    .B(_07698_),
    .C(_07700_),
    .X(_07701_));
 sky130_fd_sc_hd__a31o_1 _20410_ (.A1(_06776_),
    .A2(_07694_),
    .A3(_07696_),
    .B1(_07701_),
    .X(_07702_));
 sky130_fd_sc_hd__o22a_1 _20411_ (.A1(\datamem.data_ram[62][12] ),
    .A2(_06744_),
    .B1(_07243_),
    .B2(\datamem.data_ram[57][12] ),
    .X(_07703_));
 sky130_fd_sc_hd__o22a_1 _20412_ (.A1(\datamem.data_ram[61][12] ),
    .A2(_06661_),
    .B1(_06820_),
    .B2(\datamem.data_ram[56][12] ),
    .X(_07704_));
 sky130_fd_sc_hd__o221a_1 _20413_ (.A1(\datamem.data_ram[58][12] ),
    .A2(_06609_),
    .B1(_06617_),
    .B2(\datamem.data_ram[60][12] ),
    .C1(_06598_),
    .X(_07705_));
 sky130_fd_sc_hd__o211a_1 _20414_ (.A1(\datamem.data_ram[63][12] ),
    .A2(_06705_),
    .B1(_07704_),
    .C1(_07705_),
    .X(_07706_));
 sky130_fd_sc_hd__o211a_1 _20415_ (.A1(\datamem.data_ram[59][12] ),
    .A2(_06737_),
    .B1(_07703_),
    .C1(_07706_),
    .X(_07707_));
 sky130_fd_sc_hd__o22a_1 _20416_ (.A1(\datamem.data_ram[53][12] ),
    .A2(_06662_),
    .B1(_07243_),
    .B2(\datamem.data_ram[49][12] ),
    .X(_07708_));
 sky130_fd_sc_hd__o22a_1 _20417_ (.A1(\datamem.data_ram[55][12] ),
    .A2(_06667_),
    .B1(_06684_),
    .B2(\datamem.data_ram[52][12] ),
    .X(_07709_));
 sky130_fd_sc_hd__o221a_1 _20418_ (.A1(\datamem.data_ram[54][12] ),
    .A2(_06743_),
    .B1(_06645_),
    .B2(\datamem.data_ram[48][12] ),
    .C1(_07709_),
    .X(_07710_));
 sky130_fd_sc_hd__o211a_1 _20419_ (.A1(\datamem.data_ram[51][12] ),
    .A2(_06633_),
    .B1(_07710_),
    .C1(_06678_),
    .X(_07711_));
 sky130_fd_sc_hd__o211a_1 _20420_ (.A1(\datamem.data_ram[50][12] ),
    .A2(_06691_),
    .B1(_07708_),
    .C1(_07711_),
    .X(_07712_));
 sky130_fd_sc_hd__or3_1 _20421_ (.A(_06751_),
    .B(_07707_),
    .C(_07712_),
    .X(_07713_));
 sky130_fd_sc_hd__o211a_1 _20422_ (.A1(_06715_),
    .A2(_07702_),
    .B1(_07713_),
    .C1(_06712_),
    .X(_07714_));
 sky130_fd_sc_hd__o22a_1 _20423_ (.A1(\datamem.data_ram[7][12] ),
    .A2(_06706_),
    .B1(_07230_),
    .B2(\datamem.data_ram[4][12] ),
    .X(_07715_));
 sky130_fd_sc_hd__o22a_1 _20424_ (.A1(\datamem.data_ram[2][12] ),
    .A2(_06610_),
    .B1(_06815_),
    .B2(\datamem.data_ram[5][12] ),
    .X(_07716_));
 sky130_fd_sc_hd__o221a_1 _20425_ (.A1(\datamem.data_ram[3][12] ),
    .A2(_06633_),
    .B1(_07243_),
    .B2(\datamem.data_ram[1][12] ),
    .C1(_06678_),
    .X(_07717_));
 sky130_fd_sc_hd__o211a_1 _20426_ (.A1(\datamem.data_ram[0][12] ),
    .A2(_06647_),
    .B1(_07716_),
    .C1(_07717_),
    .X(_07718_));
 sky130_fd_sc_hd__o211a_1 _20427_ (.A1(\datamem.data_ram[6][12] ),
    .A2(_06629_),
    .B1(_07715_),
    .C1(_07718_),
    .X(_07719_));
 sky130_fd_sc_hd__o22a_1 _20428_ (.A1(\datamem.data_ram[13][12] ),
    .A2(_06663_),
    .B1(_06647_),
    .B2(\datamem.data_ram[8][12] ),
    .X(_07720_));
 sky130_fd_sc_hd__o22a_1 _20429_ (.A1(\datamem.data_ram[11][12] ),
    .A2(_06632_),
    .B1(_06780_),
    .B2(\datamem.data_ram[9][12] ),
    .X(_07721_));
 sky130_fd_sc_hd__o221a_1 _20430_ (.A1(\datamem.data_ram[14][12] ),
    .A2(_07085_),
    .B1(_06618_),
    .B2(\datamem.data_ram[12][12] ),
    .C1(_07721_),
    .X(_07722_));
 sky130_fd_sc_hd__o211a_1 _20431_ (.A1(\datamem.data_ram[15][12] ),
    .A2(_06784_),
    .B1(_07722_),
    .C1(_06601_),
    .X(_07723_));
 sky130_fd_sc_hd__o211a_1 _20432_ (.A1(\datamem.data_ram[10][12] ),
    .A2(_06612_),
    .B1(_07720_),
    .C1(_07723_),
    .X(_07724_));
 sky130_fd_sc_hd__o22a_1 _20433_ (.A1(\datamem.data_ram[16][12] ),
    .A2(_06646_),
    .B1(_06618_),
    .B2(\datamem.data_ram[20][12] ),
    .X(_07725_));
 sky130_fd_sc_hd__o22a_1 _20434_ (.A1(\datamem.data_ram[21][12] ),
    .A2(_06661_),
    .B1(_06704_),
    .B2(\datamem.data_ram[23][12] ),
    .X(_07726_));
 sky130_fd_sc_hd__o221a_1 _20435_ (.A1(\datamem.data_ram[19][12] ),
    .A2(_06632_),
    .B1(_06780_),
    .B2(\datamem.data_ram[17][12] ),
    .C1(_06677_),
    .X(_07727_));
 sky130_fd_sc_hd__o211a_1 _20436_ (.A1(\datamem.data_ram[22][12] ),
    .A2(_07085_),
    .B1(_07726_),
    .C1(_07727_),
    .X(_07728_));
 sky130_fd_sc_hd__o211a_1 _20437_ (.A1(\datamem.data_ram[18][12] ),
    .A2(_06611_),
    .B1(_07725_),
    .C1(_07728_),
    .X(_07729_));
 sky130_fd_sc_hd__o22a_1 _20438_ (.A1(\datamem.data_ram[26][12] ),
    .A2(_06610_),
    .B1(_06821_),
    .B2(\datamem.data_ram[24][12] ),
    .X(_07730_));
 sky130_fd_sc_hd__o22a_1 _20439_ (.A1(\datamem.data_ram[29][12] ),
    .A2(_06721_),
    .B1(_06654_),
    .B2(\datamem.data_ram[25][12] ),
    .X(_07731_));
 sky130_fd_sc_hd__o221a_1 _20440_ (.A1(\datamem.data_ram[30][12] ),
    .A2(_06743_),
    .B1(_06617_),
    .B2(\datamem.data_ram[28][12] ),
    .C1(_07731_),
    .X(_07732_));
 sky130_fd_sc_hd__o211a_1 _20441_ (.A1(\datamem.data_ram[31][12] ),
    .A2(_06705_),
    .B1(_07732_),
    .C1(_06600_),
    .X(_07733_));
 sky130_fd_sc_hd__o211a_1 _20442_ (.A1(\datamem.data_ram[27][12] ),
    .A2(_06634_),
    .B1(_07730_),
    .C1(_07733_),
    .X(_07734_));
 sky130_fd_sc_hd__or3_1 _20443_ (.A(_06751_),
    .B(_07729_),
    .C(_07734_),
    .X(_07735_));
 sky130_fd_sc_hd__o311a_1 _20444_ (.A1(_06715_),
    .A2(_07719_),
    .A3(_07724_),
    .B1(_06860_),
    .C1(_07735_),
    .X(_07736_));
 sky130_fd_sc_hd__nor2_4 _20445_ (.A(_07714_),
    .B(_07736_),
    .Y(_07737_));
 sky130_fd_sc_hd__o22a_1 _20446_ (.A1(\datamem.data_ram[5][20] ),
    .A2(_06702_),
    .B1(_06706_),
    .B2(\datamem.data_ram[7][20] ),
    .X(_07738_));
 sky130_fd_sc_hd__o221a_1 _20447_ (.A1(\datamem.data_ram[6][20] ),
    .A2(_06764_),
    .B1(_06779_),
    .B2(\datamem.data_ram[0][20] ),
    .C1(_07738_),
    .X(_07739_));
 sky130_fd_sc_hd__o22a_1 _20448_ (.A1(\datamem.data_ram[2][20] ),
    .A2(_06691_),
    .B1(_06619_),
    .B2(\datamem.data_ram[4][20] ),
    .X(_07740_));
 sky130_fd_sc_hd__o221a_1 _20449_ (.A1(\datamem.data_ram[3][20] ),
    .A2(_06738_),
    .B1(_06700_),
    .B2(\datamem.data_ram[1][20] ),
    .C1(_07740_),
    .X(_07741_));
 sky130_fd_sc_hd__o22a_1 _20450_ (.A1(\datamem.data_ram[11][20] ),
    .A2(_06730_),
    .B1(_06705_),
    .B2(\datamem.data_ram[15][20] ),
    .X(_07742_));
 sky130_fd_sc_hd__o221a_1 _20451_ (.A1(\datamem.data_ram[13][20] ),
    .A2(_06768_),
    .B1(_06699_),
    .B2(\datamem.data_ram[9][20] ),
    .C1(_07742_),
    .X(_07743_));
 sky130_fd_sc_hd__o22a_1 _20452_ (.A1(\datamem.data_ram[14][20] ),
    .A2(_06744_),
    .B1(_06765_),
    .B2(\datamem.data_ram[12][20] ),
    .X(_07744_));
 sky130_fd_sc_hd__o221a_1 _20453_ (.A1(\datamem.data_ram[10][20] ),
    .A2(_06728_),
    .B1(_06778_),
    .B2(\datamem.data_ram[8][20] ),
    .C1(_07744_),
    .X(_07745_));
 sky130_fd_sc_hd__and3_1 _20454_ (.A(_06742_),
    .B(_07743_),
    .C(_07745_),
    .X(_07746_));
 sky130_fd_sc_hd__a31o_1 _20455_ (.A1(_06680_),
    .A2(_07739_),
    .A3(_07741_),
    .B1(_07746_),
    .X(_07747_));
 sky130_fd_sc_hd__o22a_1 _20456_ (.A1(\datamem.data_ram[30][20] ),
    .A2(_06628_),
    .B1(_07230_),
    .B2(\datamem.data_ram[28][20] ),
    .X(_07748_));
 sky130_fd_sc_hd__o22a_1 _20457_ (.A1(\datamem.data_ram[24][20] ),
    .A2(_06821_),
    .B1(_06781_),
    .B2(\datamem.data_ram[25][20] ),
    .X(_07749_));
 sky130_fd_sc_hd__o221a_1 _20458_ (.A1(\datamem.data_ram[26][20] ),
    .A2(_06690_),
    .B1(_06633_),
    .B2(\datamem.data_ram[27][20] ),
    .C1(_06600_),
    .X(_07750_));
 sky130_fd_sc_hd__o211a_1 _20459_ (.A1(\datamem.data_ram[29][20] ),
    .A2(_06663_),
    .B1(_07749_),
    .C1(_07750_),
    .X(_07751_));
 sky130_fd_sc_hd__o211a_1 _20460_ (.A1(\datamem.data_ram[31][20] ),
    .A2(_06707_),
    .B1(_07748_),
    .C1(_07751_),
    .X(_07752_));
 sky130_fd_sc_hd__o22a_1 _20461_ (.A1(\datamem.data_ram[18][20] ),
    .A2(_06611_),
    .B1(_06782_),
    .B2(\datamem.data_ram[17][20] ),
    .X(_07753_));
 sky130_fd_sc_hd__o22a_1 _20462_ (.A1(\datamem.data_ram[21][20] ),
    .A2(_06661_),
    .B1(_06704_),
    .B2(\datamem.data_ram[23][20] ),
    .X(_07754_));
 sky130_fd_sc_hd__o221a_1 _20463_ (.A1(\datamem.data_ram[22][20] ),
    .A2(_07085_),
    .B1(_06646_),
    .B2(\datamem.data_ram[16][20] ),
    .C1(_07754_),
    .X(_07755_));
 sky130_fd_sc_hd__o211a_1 _20464_ (.A1(\datamem.data_ram[20][20] ),
    .A2(_07230_),
    .B1(_07755_),
    .C1(_06679_),
    .X(_07756_));
 sky130_fd_sc_hd__o211a_1 _20465_ (.A1(\datamem.data_ram[19][20] ),
    .A2(_06635_),
    .B1(_07753_),
    .C1(_07756_),
    .X(_07757_));
 sky130_fd_sc_hd__o21a_1 _20466_ (.A1(_07752_),
    .A2(_07757_),
    .B1(_06796_),
    .X(_07758_));
 sky130_fd_sc_hd__o22a_1 _20467_ (.A1(\datamem.data_ram[45][20] ),
    .A2(_06702_),
    .B1(_06619_),
    .B2(\datamem.data_ram[44][20] ),
    .X(_07759_));
 sky130_fd_sc_hd__o22a_1 _20468_ (.A1(\datamem.data_ram[42][20] ),
    .A2(_06609_),
    .B1(_07242_),
    .B2(\datamem.data_ram[41][20] ),
    .X(_07760_));
 sky130_fd_sc_hd__o221a_1 _20469_ (.A1(\datamem.data_ram[46][20] ),
    .A2(_06744_),
    .B1(_06725_),
    .B2(\datamem.data_ram[47][20] ),
    .C1(_07760_),
    .X(_07761_));
 sky130_fd_sc_hd__o211a_1 _20470_ (.A1(\datamem.data_ram[40][20] ),
    .A2(_06778_),
    .B1(_07761_),
    .C1(_06601_),
    .X(_07762_));
 sky130_fd_sc_hd__o211a_1 _20471_ (.A1(\datamem.data_ram[43][20] ),
    .A2(_06635_),
    .B1(_07759_),
    .C1(_07762_),
    .X(_07763_));
 sky130_fd_sc_hd__o22a_1 _20472_ (.A1(\datamem.data_ram[38][20] ),
    .A2(_06628_),
    .B1(_07230_),
    .B2(\datamem.data_ram[36][20] ),
    .X(_07764_));
 sky130_fd_sc_hd__o22a_1 _20473_ (.A1(\datamem.data_ram[37][20] ),
    .A2(_06662_),
    .B1(_06781_),
    .B2(\datamem.data_ram[33][20] ),
    .X(_07765_));
 sky130_fd_sc_hd__o221a_1 _20474_ (.A1(\datamem.data_ram[34][20] ),
    .A2(_06690_),
    .B1(_06633_),
    .B2(\datamem.data_ram[35][20] ),
    .C1(_06678_),
    .X(_07766_));
 sky130_fd_sc_hd__o211a_1 _20475_ (.A1(\datamem.data_ram[39][20] ),
    .A2(_06706_),
    .B1(_07765_),
    .C1(_07766_),
    .X(_07767_));
 sky130_fd_sc_hd__o211a_1 _20476_ (.A1(\datamem.data_ram[32][20] ),
    .A2(_06779_),
    .B1(_07764_),
    .C1(_07767_),
    .X(_07768_));
 sky130_fd_sc_hd__o22a_1 _20477_ (.A1(\datamem.data_ram[53][20] ),
    .A2(_06662_),
    .B1(_06705_),
    .B2(\datamem.data_ram[55][20] ),
    .X(_07769_));
 sky130_fd_sc_hd__o22a_1 _20478_ (.A1(\datamem.data_ram[54][20] ),
    .A2(_06743_),
    .B1(_06820_),
    .B2(\datamem.data_ram[48][20] ),
    .X(_07770_));
 sky130_fd_sc_hd__o221a_1 _20479_ (.A1(\datamem.data_ram[50][20] ),
    .A2(_06609_),
    .B1(_06632_),
    .B2(\datamem.data_ram[51][20] ),
    .C1(_06677_),
    .X(_07771_));
 sky130_fd_sc_hd__o211a_1 _20480_ (.A1(\datamem.data_ram[52][20] ),
    .A2(_06618_),
    .B1(_07770_),
    .C1(_07771_),
    .X(_07772_));
 sky130_fd_sc_hd__o211a_1 _20481_ (.A1(\datamem.data_ram[49][20] ),
    .A2(_06782_),
    .B1(_07769_),
    .C1(_07772_),
    .X(_07773_));
 sky130_fd_sc_hd__o22a_1 _20482_ (.A1(\datamem.data_ram[62][20] ),
    .A2(_06627_),
    .B1(_06815_),
    .B2(\datamem.data_ram[61][20] ),
    .X(_07774_));
 sky130_fd_sc_hd__o22a_1 _20483_ (.A1(\datamem.data_ram[63][20] ),
    .A2(_06668_),
    .B1(_06654_),
    .B2(\datamem.data_ram[57][20] ),
    .X(_07775_));
 sky130_fd_sc_hd__o221a_1 _20484_ (.A1(\datamem.data_ram[56][20] ),
    .A2(_06820_),
    .B1(_06617_),
    .B2(\datamem.data_ram[60][20] ),
    .C1(_07775_),
    .X(_07776_));
 sky130_fd_sc_hd__o211a_1 _20485_ (.A1(\datamem.data_ram[58][20] ),
    .A2(_06610_),
    .B1(_06600_),
    .C1(_07776_),
    .X(_07777_));
 sky130_fd_sc_hd__o211a_1 _20486_ (.A1(\datamem.data_ram[59][20] ),
    .A2(_06634_),
    .B1(_07774_),
    .C1(_07777_),
    .X(_07778_));
 sky130_fd_sc_hd__o31a_1 _20487_ (.A1(_06751_),
    .A2(_07773_),
    .A3(_07778_),
    .B1(_06594_),
    .X(_07779_));
 sky130_fd_sc_hd__o31a_1 _20488_ (.A1(_06715_),
    .A2(_07763_),
    .A3(_07768_),
    .B1(_07779_),
    .X(_07780_));
 sky130_fd_sc_hd__a211oi_4 _20489_ (.A1(_06596_),
    .A2(_07747_),
    .B1(_07758_),
    .C1(_07780_),
    .Y(_07781_));
 sky130_fd_sc_hd__o22a_1 _20490_ (.A1(\rvcpu.dp.plem.ALUResultM[1] ),
    .A2(_07737_),
    .B1(_07781_),
    .B2(\rvcpu.dp.plem.ALUResultM[0] ),
    .X(_07782_));
 sky130_fd_sc_hd__and3b_1 _20491_ (.A_N(_06589_),
    .B(_07692_),
    .C(_07782_),
    .X(_07783_));
 sky130_fd_sc_hd__a211o_1 _20492_ (.A1(_06589_),
    .A2(_07646_),
    .B1(_07783_),
    .C1(_06583_),
    .X(_07784_));
 sky130_fd_sc_hd__o22a_1 _20493_ (.A1(_06915_),
    .A2(_07781_),
    .B1(_07646_),
    .B2(_07277_),
    .X(_07785_));
 sky130_fd_sc_hd__nand2_1 _20494_ (.A(_07784_),
    .B(_07785_),
    .Y(_04441_));
 sky130_fd_sc_hd__o22a_1 _20495_ (.A1(\datamem.data_ram[34][21] ),
    .A2(_06613_),
    .B1(_06701_),
    .B2(\datamem.data_ram[33][21] ),
    .X(_07786_));
 sky130_fd_sc_hd__o221a_1 _20496_ (.A1(\datamem.data_ram[37][21] ),
    .A2(_06665_),
    .B1(_07021_),
    .B2(\datamem.data_ram[39][21] ),
    .C1(_07786_),
    .X(_07787_));
 sky130_fd_sc_hd__o22a_1 _20497_ (.A1(\datamem.data_ram[38][21] ),
    .A2(_06630_),
    .B1(_06688_),
    .B2(\datamem.data_ram[36][21] ),
    .X(_07788_));
 sky130_fd_sc_hd__o221a_1 _20498_ (.A1(\datamem.data_ram[32][21] ),
    .A2(_06649_),
    .B1(_07077_),
    .B2(\datamem.data_ram[35][21] ),
    .C1(_07788_),
    .X(_07789_));
 sky130_fd_sc_hd__and3_1 _20499_ (.A(_07131_),
    .B(_07787_),
    .C(_07789_),
    .X(_07790_));
 sky130_fd_sc_hd__buf_4 _20500_ (.A(_07021_),
    .X(_07791_));
 sky130_fd_sc_hd__o22a_1 _20501_ (.A1(\datamem.data_ram[47][21] ),
    .A2(_07791_),
    .B1(_07182_),
    .B2(\datamem.data_ram[44][21] ),
    .X(_07792_));
 sky130_fd_sc_hd__o22a_1 _20502_ (.A1(\datamem.data_ram[46][21] ),
    .A2(_06630_),
    .B1(_06701_),
    .B2(\datamem.data_ram[41][21] ),
    .X(_07793_));
 sky130_fd_sc_hd__o221a_1 _20503_ (.A1(\datamem.data_ram[40][21] ),
    .A2(_06698_),
    .B1(_06636_),
    .B2(\datamem.data_ram[43][21] ),
    .C1(_07081_),
    .X(_07794_));
 sky130_fd_sc_hd__o211a_1 _20504_ (.A1(\datamem.data_ram[42][21] ),
    .A2(_07203_),
    .B1(_07793_),
    .C1(_07794_),
    .X(_07795_));
 sky130_fd_sc_hd__o211a_1 _20505_ (.A1(\datamem.data_ram[45][21] ),
    .A2(_07019_),
    .B1(_07792_),
    .C1(_07795_),
    .X(_07796_));
 sky130_fd_sc_hd__o22a_1 _20506_ (.A1(\datamem.data_ram[55][21] ),
    .A2(_07021_),
    .B1(_06701_),
    .B2(\datamem.data_ram[49][21] ),
    .X(_07797_));
 sky130_fd_sc_hd__o221a_1 _20507_ (.A1(\datamem.data_ram[48][21] ),
    .A2(_07191_),
    .B1(_07182_),
    .B2(\datamem.data_ram[52][21] ),
    .C1(_07797_),
    .X(_07798_));
 sky130_fd_sc_hd__o22a_1 _20508_ (.A1(\datamem.data_ram[54][21] ),
    .A2(_06630_),
    .B1(_06665_),
    .B2(\datamem.data_ram[53][21] ),
    .X(_07799_));
 sky130_fd_sc_hd__o221a_1 _20509_ (.A1(\datamem.data_ram[50][21] ),
    .A2(_06613_),
    .B1(_07077_),
    .B2(\datamem.data_ram[51][21] ),
    .C1(_07799_),
    .X(_07800_));
 sky130_fd_sc_hd__and3_1 _20510_ (.A(_07131_),
    .B(_07798_),
    .C(_07800_),
    .X(_07801_));
 sky130_fd_sc_hd__o22a_1 _20511_ (.A1(\datamem.data_ram[61][21] ),
    .A2(_06665_),
    .B1(_06636_),
    .B2(\datamem.data_ram[59][21] ),
    .X(_07802_));
 sky130_fd_sc_hd__o221a_1 _20512_ (.A1(\datamem.data_ram[62][21] ),
    .A2(_07028_),
    .B1(_06659_),
    .B2(\datamem.data_ram[57][21] ),
    .C1(_07802_),
    .X(_07803_));
 sky130_fd_sc_hd__o22a_1 _20513_ (.A1(\datamem.data_ram[56][21] ),
    .A2(_06649_),
    .B1(_06621_),
    .B2(\datamem.data_ram[60][21] ),
    .X(_07804_));
 sky130_fd_sc_hd__o221a_1 _20514_ (.A1(\datamem.data_ram[58][21] ),
    .A2(_06613_),
    .B1(_07791_),
    .B2(\datamem.data_ram[63][21] ),
    .C1(_07804_),
    .X(_07805_));
 sky130_fd_sc_hd__a31o_1 _20515_ (.A1(_06604_),
    .A2(_07803_),
    .A3(_07805_),
    .B1(_06916_),
    .X(_07806_));
 sky130_fd_sc_hd__o32a_2 _20516_ (.A1(_07071_),
    .A2(_07790_),
    .A3(_07796_),
    .B1(_07801_),
    .B2(_07806_),
    .X(_07807_));
 sky130_fd_sc_hd__clkbuf_8 _20517_ (.A(_06659_),
    .X(_07808_));
 sky130_fd_sc_hd__o22a_1 _20518_ (.A1(\datamem.data_ram[30][21] ),
    .A2(_07028_),
    .B1(_07808_),
    .B2(\datamem.data_ram[25][21] ),
    .X(_07809_));
 sky130_fd_sc_hd__o22a_1 _20519_ (.A1(\datamem.data_ram[29][21] ),
    .A2(_06865_),
    .B1(_06672_),
    .B2(\datamem.data_ram[31][21] ),
    .X(_07810_));
 sky130_fd_sc_hd__o221a_1 _20520_ (.A1(\datamem.data_ram[24][21] ),
    .A2(_06649_),
    .B1(_06621_),
    .B2(\datamem.data_ram[28][21] ),
    .C1(_07810_),
    .X(_07811_));
 sky130_fd_sc_hd__o211a_1 _20521_ (.A1(\datamem.data_ram[26][21] ),
    .A2(_07203_),
    .B1(_06604_),
    .C1(_07811_),
    .X(_07812_));
 sky130_fd_sc_hd__o211a_1 _20522_ (.A1(\datamem.data_ram[27][21] ),
    .A2(_07077_),
    .B1(_07809_),
    .C1(_07812_),
    .X(_07813_));
 sky130_fd_sc_hd__o22a_1 _20523_ (.A1(\datamem.data_ram[22][21] ),
    .A2(_07028_),
    .B1(_07182_),
    .B2(\datamem.data_ram[20][21] ),
    .X(_07814_));
 sky130_fd_sc_hd__o22a_1 _20524_ (.A1(\datamem.data_ram[23][21] ),
    .A2(_07021_),
    .B1(_06659_),
    .B2(\datamem.data_ram[17][21] ),
    .X(_07815_));
 sky130_fd_sc_hd__o221a_1 _20525_ (.A1(\datamem.data_ram[16][21] ),
    .A2(_06649_),
    .B1(_06636_),
    .B2(\datamem.data_ram[19][21] ),
    .C1(_06777_),
    .X(_07816_));
 sky130_fd_sc_hd__o211a_1 _20526_ (.A1(\datamem.data_ram[21][21] ),
    .A2(_07019_),
    .B1(_07815_),
    .C1(_07816_),
    .X(_07817_));
 sky130_fd_sc_hd__o211a_1 _20527_ (.A1(\datamem.data_ram[18][21] ),
    .A2(_07203_),
    .B1(_07814_),
    .C1(_07817_),
    .X(_07818_));
 sky130_fd_sc_hd__clkbuf_8 _20528_ (.A(_06640_),
    .X(_07819_));
 sky130_fd_sc_hd__buf_8 _20529_ (.A(_07819_),
    .X(_07820_));
 sky130_fd_sc_hd__buf_6 _20530_ (.A(_07820_),
    .X(_07821_));
 sky130_fd_sc_hd__buf_8 _20531_ (.A(_07821_),
    .X(_07822_));
 sky130_fd_sc_hd__clkbuf_8 _20532_ (.A(_06605_),
    .X(_07823_));
 sky130_fd_sc_hd__buf_8 _20533_ (.A(_06652_),
    .X(_07824_));
 sky130_fd_sc_hd__buf_6 _20534_ (.A(_07824_),
    .X(_07825_));
 sky130_fd_sc_hd__buf_6 _20535_ (.A(_07825_),
    .X(_07826_));
 sky130_fd_sc_hd__buf_6 _20536_ (.A(_07826_),
    .X(_07827_));
 sky130_fd_sc_hd__buf_6 _20537_ (.A(_07827_),
    .X(_07828_));
 sky130_fd_sc_hd__buf_6 _20538_ (.A(_07828_),
    .X(_07829_));
 sky130_fd_sc_hd__a22o_1 _20539_ (.A1(_07823_),
    .A2(\datamem.data_ram[6][21] ),
    .B1(\datamem.data_ram[7][21] ),
    .B2(_07829_),
    .X(_07830_));
 sky130_fd_sc_hd__buf_6 _20540_ (.A(_06944_),
    .X(_07831_));
 sky130_fd_sc_hd__buf_6 _20541_ (.A(_07831_),
    .X(_07832_));
 sky130_fd_sc_hd__buf_6 _20542_ (.A(_07832_),
    .X(_07833_));
 sky130_fd_sc_hd__or2_1 _20543_ (.A(\datamem.data_ram[5][21] ),
    .B(_07833_),
    .X(_07834_));
 sky130_fd_sc_hd__buf_6 _20544_ (.A(_07826_),
    .X(_07835_));
 sky130_fd_sc_hd__buf_8 _20545_ (.A(_07835_),
    .X(_07836_));
 sky130_fd_sc_hd__buf_6 _20546_ (.A(_07836_),
    .X(_07837_));
 sky130_fd_sc_hd__buf_8 _20547_ (.A(_06606_),
    .X(_07838_));
 sky130_fd_sc_hd__buf_6 _20548_ (.A(_07838_),
    .X(_07839_));
 sky130_fd_sc_hd__buf_6 _20549_ (.A(_07839_),
    .X(_07840_));
 sky130_fd_sc_hd__o21a_1 _20550_ (.A1(\datamem.data_ram[4][21] ),
    .A2(_07837_),
    .B1(_07840_),
    .X(_07841_));
 sky130_fd_sc_hd__a22o_1 _20551_ (.A1(_07822_),
    .A2(_07830_),
    .B1(_07834_),
    .B2(_07841_),
    .X(_07842_));
 sky130_fd_sc_hd__mux4_1 _20552_ (.A0(\datamem.data_ram[0][21] ),
    .A1(\datamem.data_ram[1][21] ),
    .A2(\datamem.data_ram[2][21] ),
    .A3(\datamem.data_ram[3][21] ),
    .S0(_07837_),
    .S1(_07822_),
    .X(_07843_));
 sky130_fd_sc_hd__buf_6 _20553_ (.A(_06614_),
    .X(_07844_));
 sky130_fd_sc_hd__buf_6 _20554_ (.A(_07844_),
    .X(_07845_));
 sky130_fd_sc_hd__mux2_1 _20555_ (.A0(_07842_),
    .A1(_07843_),
    .S(_07845_),
    .X(_07846_));
 sky130_fd_sc_hd__o22a_1 _20556_ (.A1(\datamem.data_ram[14][21] ),
    .A2(_07028_),
    .B1(_06649_),
    .B2(\datamem.data_ram[8][21] ),
    .X(_07847_));
 sky130_fd_sc_hd__o22a_1 _20557_ (.A1(\datamem.data_ram[15][21] ),
    .A2(_07020_),
    .B1(_06688_),
    .B2(\datamem.data_ram[12][21] ),
    .X(_07848_));
 sky130_fd_sc_hd__clkbuf_8 _20558_ (.A(_07835_),
    .X(_07849_));
 sky130_fd_sc_hd__a22o_1 _20559_ (.A1(_07823_),
    .A2(\datamem.data_ram[10][21] ),
    .B1(\datamem.data_ram[11][21] ),
    .B2(_07849_),
    .X(_07850_));
 sky130_fd_sc_hd__buf_6 _20560_ (.A(_06940_),
    .X(_07851_));
 sky130_fd_sc_hd__o22a_1 _20561_ (.A1(\datamem.data_ram[13][21] ),
    .A2(_06664_),
    .B1(_07850_),
    .B2(_07851_),
    .X(_07852_));
 sky130_fd_sc_hd__and3_1 _20562_ (.A(_06603_),
    .B(_07848_),
    .C(_07852_),
    .X(_07853_));
 sky130_fd_sc_hd__o211a_1 _20563_ (.A1(\datamem.data_ram[9][21] ),
    .A2(_07808_),
    .B1(_07847_),
    .C1(_07853_),
    .X(_07854_));
 sky130_fd_sc_hd__a211o_1 _20564_ (.A1(_07131_),
    .A2(_07846_),
    .B1(_07854_),
    .C1(_07154_),
    .X(_07855_));
 sky130_fd_sc_hd__o31a_1 _20565_ (.A1(_07177_),
    .A2(_07813_),
    .A3(_07818_),
    .B1(_07855_),
    .X(_07856_));
 sky130_fd_sc_hd__o21ai_2 _20566_ (.A1(_06985_),
    .A2(_07807_),
    .B1(_07856_),
    .Y(_07857_));
 sky130_fd_sc_hd__nor2_4 _20567_ (.A(\rvcpu.dp.plem.ALUResultM[6] ),
    .B(_06860_),
    .Y(_07858_));
 sky130_fd_sc_hd__buf_4 _20568_ (.A(_06922_),
    .X(_07859_));
 sky130_fd_sc_hd__buf_6 _20569_ (.A(_07859_),
    .X(_07860_));
 sky130_fd_sc_hd__mux2_1 _20570_ (.A0(\datamem.data_ram[38][13] ),
    .A1(\datamem.data_ram[39][13] ),
    .S(_07829_),
    .X(_07861_));
 sky130_fd_sc_hd__buf_4 _20571_ (.A(_06917_),
    .X(_07862_));
 sky130_fd_sc_hd__clkbuf_8 _20572_ (.A(_07862_),
    .X(_07863_));
 sky130_fd_sc_hd__mux2_1 _20573_ (.A0(\datamem.data_ram[36][13] ),
    .A1(\datamem.data_ram[37][13] ),
    .S(_07828_),
    .X(_07864_));
 sky130_fd_sc_hd__mux4_1 _20574_ (.A0(\datamem.data_ram[32][13] ),
    .A1(\datamem.data_ram[33][13] ),
    .A2(\datamem.data_ram[34][13] ),
    .A3(\datamem.data_ram[35][13] ),
    .S0(_07835_),
    .S1(_07821_),
    .X(_07865_));
 sky130_fd_sc_hd__buf_6 _20575_ (.A(_06641_),
    .X(_07866_));
 sky130_fd_sc_hd__clkbuf_8 _20576_ (.A(_07866_),
    .X(_07867_));
 sky130_fd_sc_hd__clkbuf_8 _20577_ (.A(_07867_),
    .X(_07868_));
 sky130_fd_sc_hd__o22a_1 _20578_ (.A1(_07863_),
    .A2(_07864_),
    .B1(_07865_),
    .B2(_07868_),
    .X(_07869_));
 sky130_fd_sc_hd__o21ai_1 _20579_ (.A1(_07860_),
    .A2(_07861_),
    .B1(_07869_),
    .Y(_07870_));
 sky130_fd_sc_hd__a21oi_1 _20580_ (.A1(_07858_),
    .A2(_07870_),
    .B1(_06603_),
    .Y(_07871_));
 sky130_fd_sc_hd__nand2_8 _20581_ (.A(\rvcpu.dp.plem.ALUResultM[7] ),
    .B(_06592_),
    .Y(_07872_));
 sky130_fd_sc_hd__a22o_1 _20582_ (.A1(_07635_),
    .A2(\datamem.data_ram[51][13] ),
    .B1(_07831_),
    .B2(\datamem.data_ram[50][13] ),
    .X(_07873_));
 sky130_fd_sc_hd__buf_8 _20583_ (.A(_07824_),
    .X(_07874_));
 sky130_fd_sc_hd__mux2_1 _20584_ (.A0(\datamem.data_ram[48][13] ),
    .A1(\datamem.data_ram[49][13] ),
    .S(_07874_),
    .X(_07875_));
 sky130_fd_sc_hd__or2_1 _20585_ (.A(_07867_),
    .B(_07875_),
    .X(_07876_));
 sky130_fd_sc_hd__a22o_1 _20586_ (.A1(_07821_),
    .A2(_07873_),
    .B1(_07876_),
    .B2(_06940_),
    .X(_07877_));
 sky130_fd_sc_hd__o221a_1 _20587_ (.A1(\datamem.data_ram[54][13] ),
    .A2(_06628_),
    .B1(_06706_),
    .B2(\datamem.data_ram[55][13] ),
    .C1(_07877_),
    .X(_07878_));
 sky130_fd_sc_hd__o221a_1 _20588_ (.A1(\datamem.data_ram[53][13] ),
    .A2(_06703_),
    .B1(_06620_),
    .B2(\datamem.data_ram[52][13] ),
    .C1(_07878_),
    .X(_07879_));
 sky130_fd_sc_hd__mux2_1 _20589_ (.A0(\datamem.data_ram[16][13] ),
    .A1(\datamem.data_ram[17][13] ),
    .S(_07826_),
    .X(_07880_));
 sky130_fd_sc_hd__or2_1 _20590_ (.A(_06666_),
    .B(\datamem.data_ram[18][13] ),
    .X(_07881_));
 sky130_fd_sc_hd__o211a_1 _20591_ (.A1(\datamem.data_ram[19][13] ),
    .A2(_07831_),
    .B1(_07881_),
    .C1(_07820_),
    .X(_07882_));
 sky130_fd_sc_hd__a211o_1 _20592_ (.A1(_07839_),
    .A2(_07880_),
    .B1(_07882_),
    .C1(_07867_),
    .X(_07883_));
 sky130_fd_sc_hd__o221a_1 _20593_ (.A1(\datamem.data_ram[22][13] ),
    .A2(_06628_),
    .B1(_07230_),
    .B2(\datamem.data_ram[20][13] ),
    .C1(_07883_),
    .X(_07884_));
 sky130_fd_sc_hd__o221a_1 _20594_ (.A1(\datamem.data_ram[21][13] ),
    .A2(_06664_),
    .B1(_07020_),
    .B2(\datamem.data_ram[23][13] ),
    .C1(_07884_),
    .X(_07885_));
 sky130_fd_sc_hd__mux2_1 _20595_ (.A0(\datamem.data_ram[0][13] ),
    .A1(\datamem.data_ram[1][13] ),
    .S(_07827_),
    .X(_07886_));
 sky130_fd_sc_hd__or2_1 _20596_ (.A(\datamem.data_ram[2][13] ),
    .B(_07826_),
    .X(_07887_));
 sky130_fd_sc_hd__o211a_1 _20597_ (.A1(_07823_),
    .A2(\datamem.data_ram[3][13] ),
    .B1(_07821_),
    .C1(_07887_),
    .X(_07888_));
 sky130_fd_sc_hd__a211o_1 _20598_ (.A1(_07839_),
    .A2(_07886_),
    .B1(_07888_),
    .C1(_07868_),
    .X(_07889_));
 sky130_fd_sc_hd__o22a_1 _20599_ (.A1(\datamem.data_ram[5][13] ),
    .A2(_07037_),
    .B1(_06687_),
    .B2(\datamem.data_ram[4][13] ),
    .X(_07890_));
 sky130_fd_sc_hd__o22a_1 _20600_ (.A1(\datamem.data_ram[6][13] ),
    .A2(_06682_),
    .B1(_06671_),
    .B2(\datamem.data_ram[7][13] ),
    .X(_07891_));
 sky130_fd_sc_hd__a31o_1 _20601_ (.A1(_07889_),
    .A2(_07890_),
    .A3(_07891_),
    .B1(_07154_),
    .X(_07892_));
 sky130_fd_sc_hd__o221a_1 _20602_ (.A1(_07872_),
    .A2(_07879_),
    .B1(_07885_),
    .B2(_07177_),
    .C1(_07892_),
    .X(_07893_));
 sky130_fd_sc_hd__o22a_1 _20603_ (.A1(\datamem.data_ram[61][13] ),
    .A2(_06723_),
    .B1(_06731_),
    .B2(\datamem.data_ram[59][13] ),
    .X(_07894_));
 sky130_fd_sc_hd__o221a_1 _20604_ (.A1(\datamem.data_ram[56][13] ),
    .A2(_06837_),
    .B1(_06657_),
    .B2(\datamem.data_ram[57][13] ),
    .C1(_07894_),
    .X(_07895_));
 sky130_fd_sc_hd__o22a_1 _20605_ (.A1(\datamem.data_ram[58][13] ),
    .A2(_06728_),
    .B1(_06686_),
    .B2(\datamem.data_ram[60][13] ),
    .X(_07896_));
 sky130_fd_sc_hd__o221a_1 _20606_ (.A1(\datamem.data_ram[62][13] ),
    .A2(_06682_),
    .B1(_06671_),
    .B2(\datamem.data_ram[63][13] ),
    .C1(_07896_),
    .X(_07897_));
 sky130_fd_sc_hd__a21o_1 _20607_ (.A1(_07895_),
    .A2(_07897_),
    .B1(_07872_),
    .X(_07898_));
 sky130_fd_sc_hd__o22a_1 _20608_ (.A1(\datamem.data_ram[40][13] ),
    .A2(_06807_),
    .B1(_06731_),
    .B2(\datamem.data_ram[43][13] ),
    .X(_07899_));
 sky130_fd_sc_hd__o221a_1 _20609_ (.A1(\datamem.data_ram[47][13] ),
    .A2(_06784_),
    .B1(_06790_),
    .B2(\datamem.data_ram[41][13] ),
    .C1(_07899_),
    .X(_07900_));
 sky130_fd_sc_hd__o22a_1 _20610_ (.A1(\datamem.data_ram[42][13] ),
    .A2(_06804_),
    .B1(_07037_),
    .B2(\datamem.data_ram[45][13] ),
    .X(_07901_));
 sky130_fd_sc_hd__o22a_1 _20611_ (.A1(\datamem.data_ram[46][13] ),
    .A2(_06682_),
    .B1(_06806_),
    .B2(\datamem.data_ram[44][13] ),
    .X(_07902_));
 sky130_fd_sc_hd__nand2_8 _20612_ (.A(_05347_),
    .B(_06594_),
    .Y(_07903_));
 sky130_fd_sc_hd__a31o_1 _20613_ (.A1(_07900_),
    .A2(_07901_),
    .A3(_07902_),
    .B1(_07903_),
    .X(_07904_));
 sky130_fd_sc_hd__o22a_1 _20614_ (.A1(\datamem.data_ram[26][13] ),
    .A2(_06802_),
    .B1(_06661_),
    .B2(\datamem.data_ram[29][13] ),
    .X(_07905_));
 sky130_fd_sc_hd__o221a_1 _20615_ (.A1(\datamem.data_ram[31][13] ),
    .A2(_06705_),
    .B1(_06618_),
    .B2(\datamem.data_ram[28][13] ),
    .C1(_07905_),
    .X(_07906_));
 sky130_fd_sc_hd__o22a_1 _20616_ (.A1(\datamem.data_ram[24][13] ),
    .A2(_06820_),
    .B1(_06780_),
    .B2(\datamem.data_ram[25][13] ),
    .X(_07907_));
 sky130_fd_sc_hd__o221a_1 _20617_ (.A1(\datamem.data_ram[30][13] ),
    .A2(_07085_),
    .B1(_06633_),
    .B2(\datamem.data_ram[27][13] ),
    .C1(_07907_),
    .X(_07908_));
 sky130_fd_sc_hd__and2_1 _20618_ (.A(_07906_),
    .B(_07908_),
    .X(_07909_));
 sky130_fd_sc_hd__mux2_1 _20619_ (.A0(\datamem.data_ram[12][13] ),
    .A1(\datamem.data_ram[13][13] ),
    .S(_07874_),
    .X(_07910_));
 sky130_fd_sc_hd__buf_6 _20620_ (.A(_06652_),
    .X(_07911_));
 sky130_fd_sc_hd__buf_6 _20621_ (.A(_07911_),
    .X(_07912_));
 sky130_fd_sc_hd__or2_1 _20622_ (.A(\datamem.data_ram[14][13] ),
    .B(_07912_),
    .X(_07913_));
 sky130_fd_sc_hd__o211a_1 _20623_ (.A1(\datamem.data_ram[15][13] ),
    .A2(_06944_),
    .B1(_07913_),
    .C1(\rvcpu.dp.plem.ALUResultM[3] ),
    .X(_07914_));
 sky130_fd_sc_hd__a211o_1 _20624_ (.A1(_07839_),
    .A2(_07910_),
    .B1(_07914_),
    .C1(_07844_),
    .X(_07915_));
 sky130_fd_sc_hd__o221a_1 _20625_ (.A1(\datamem.data_ram[10][13] ),
    .A2(_06610_),
    .B1(_06781_),
    .B2(\datamem.data_ram[9][13] ),
    .C1(_07915_),
    .X(_07916_));
 sky130_fd_sc_hd__o221a_1 _20626_ (.A1(\datamem.data_ram[8][13] ),
    .A2(_06647_),
    .B1(_06634_),
    .B2(\datamem.data_ram[11][13] ),
    .C1(_07916_),
    .X(_07917_));
 sky130_fd_sc_hd__o221a_1 _20627_ (.A1(_07177_),
    .A2(_07909_),
    .B1(_07917_),
    .B2(_07154_),
    .C1(_06602_),
    .X(_07918_));
 sky130_fd_sc_hd__and3_1 _20628_ (.A(_07898_),
    .B(_07904_),
    .C(_07918_),
    .X(_07919_));
 sky130_fd_sc_hd__a21oi_4 _20629_ (.A1(_07871_),
    .A2(_07893_),
    .B1(_07919_),
    .Y(_07920_));
 sky130_fd_sc_hd__o22a_1 _20630_ (.A1(\datamem.data_ram[5][29] ),
    .A2(_06663_),
    .B1(_06784_),
    .B2(\datamem.data_ram[7][29] ),
    .X(_07921_));
 sky130_fd_sc_hd__o221a_1 _20631_ (.A1(\datamem.data_ram[2][29] ),
    .A2(_06612_),
    .B1(_06779_),
    .B2(\datamem.data_ram[0][29] ),
    .C1(_07921_),
    .X(_07922_));
 sky130_fd_sc_hd__o22a_1 _20632_ (.A1(\datamem.data_ram[6][29] ),
    .A2(_06628_),
    .B1(_07230_),
    .B2(\datamem.data_ram[4][29] ),
    .X(_07923_));
 sky130_fd_sc_hd__o221a_1 _20633_ (.A1(\datamem.data_ram[3][29] ),
    .A2(_06635_),
    .B1(_06783_),
    .B2(\datamem.data_ram[1][29] ),
    .C1(_07923_),
    .X(_07924_));
 sky130_fd_sc_hd__o22a_1 _20634_ (.A1(\datamem.data_ram[14][29] ),
    .A2(_06627_),
    .B1(_06781_),
    .B2(\datamem.data_ram[9][29] ),
    .X(_07925_));
 sky130_fd_sc_hd__o221a_1 _20635_ (.A1(\datamem.data_ram[13][29] ),
    .A2(_06702_),
    .B1(_06706_),
    .B2(\datamem.data_ram[15][29] ),
    .C1(_07925_),
    .X(_07926_));
 sky130_fd_sc_hd__o22a_1 _20636_ (.A1(\datamem.data_ram[10][29] ),
    .A2(_06610_),
    .B1(_06821_),
    .B2(\datamem.data_ram[8][29] ),
    .X(_07927_));
 sky130_fd_sc_hd__o221a_1 _20637_ (.A1(\datamem.data_ram[11][29] ),
    .A2(_06737_),
    .B1(_06619_),
    .B2(\datamem.data_ram[12][29] ),
    .C1(_07927_),
    .X(_07928_));
 sky130_fd_sc_hd__and3_1 _20638_ (.A(_06602_),
    .B(_07926_),
    .C(_07928_),
    .X(_07929_));
 sky130_fd_sc_hd__a31o_1 _20639_ (.A1(_06777_),
    .A2(_07922_),
    .A3(_07924_),
    .B1(_07929_),
    .X(_07930_));
 sky130_fd_sc_hd__o22a_1 _20640_ (.A1(\datamem.data_ram[22][29] ),
    .A2(_06682_),
    .B1(_06806_),
    .B2(\datamem.data_ram[20][29] ),
    .X(_07931_));
 sky130_fd_sc_hd__o22a_1 _20641_ (.A1(\datamem.data_ram[16][29] ),
    .A2(_06807_),
    .B1(_06789_),
    .B2(\datamem.data_ram[17][29] ),
    .X(_07932_));
 sky130_fd_sc_hd__o221a_1 _20642_ (.A1(\datamem.data_ram[18][29] ),
    .A2(_06803_),
    .B1(_06823_),
    .B2(\datamem.data_ram[21][29] ),
    .C1(_06733_),
    .X(_07933_));
 sky130_fd_sc_hd__o211a_1 _20643_ (.A1(\datamem.data_ram[19][29] ),
    .A2(_06829_),
    .B1(_07932_),
    .C1(_07933_),
    .X(_07934_));
 sky130_fd_sc_hd__o211a_1 _20644_ (.A1(\datamem.data_ram[23][29] ),
    .A2(_07020_),
    .B1(_07931_),
    .C1(_07934_),
    .X(_07935_));
 sky130_fd_sc_hd__o22a_1 _20645_ (.A1(\datamem.data_ram[31][29] ),
    .A2(_06671_),
    .B1(_06806_),
    .B2(\datamem.data_ram[28][29] ),
    .X(_07936_));
 sky130_fd_sc_hd__o22a_1 _20646_ (.A1(\datamem.data_ram[29][29] ),
    .A2(_06823_),
    .B1(_06807_),
    .B2(\datamem.data_ram[24][29] ),
    .X(_07937_));
 sky130_fd_sc_hd__o221a_1 _20647_ (.A1(\datamem.data_ram[26][29] ),
    .A2(_06803_),
    .B1(_06789_),
    .B2(\datamem.data_ram[25][29] ),
    .C1(_06851_),
    .X(_07938_));
 sky130_fd_sc_hd__o211a_1 _20648_ (.A1(\datamem.data_ram[30][29] ),
    .A2(_06682_),
    .B1(_07937_),
    .C1(_07938_),
    .X(_07939_));
 sky130_fd_sc_hd__o211a_1 _20649_ (.A1(\datamem.data_ram[27][29] ),
    .A2(_06863_),
    .B1(_07936_),
    .C1(_07939_),
    .X(_07940_));
 sky130_fd_sc_hd__o21a_1 _20650_ (.A1(_07935_),
    .A2(_07940_),
    .B1(_06797_),
    .X(_07941_));
 sky130_fd_sc_hd__o22a_1 _20651_ (.A1(\datamem.data_ram[37][29] ),
    .A2(_07037_),
    .B1(_06784_),
    .B2(\datamem.data_ram[39][29] ),
    .X(_07942_));
 sky130_fd_sc_hd__o22a_1 _20652_ (.A1(\datamem.data_ram[38][29] ),
    .A2(_06626_),
    .B1(_06812_),
    .B2(\datamem.data_ram[35][29] ),
    .X(_07943_));
 sky130_fd_sc_hd__o221a_1 _20653_ (.A1(\datamem.data_ram[34][29] ),
    .A2(_06610_),
    .B1(_06618_),
    .B2(\datamem.data_ram[36][29] ),
    .C1(_07943_),
    .X(_07944_));
 sky130_fd_sc_hd__o211a_1 _20654_ (.A1(\datamem.data_ram[32][29] ),
    .A2(_06647_),
    .B1(_07944_),
    .C1(_06679_),
    .X(_07945_));
 sky130_fd_sc_hd__o211a_1 _20655_ (.A1(\datamem.data_ram[33][29] ),
    .A2(_06783_),
    .B1(_07942_),
    .C1(_07945_),
    .X(_07946_));
 sky130_fd_sc_hd__o22a_1 _20656_ (.A1(\datamem.data_ram[42][29] ),
    .A2(_06804_),
    .B1(_06837_),
    .B2(\datamem.data_ram[40][29] ),
    .X(_07947_));
 sky130_fd_sc_hd__o22a_1 _20657_ (.A1(\datamem.data_ram[46][29] ),
    .A2(_06627_),
    .B1(_06805_),
    .B2(\datamem.data_ram[44][29] ),
    .X(_07948_));
 sky130_fd_sc_hd__o221a_1 _20658_ (.A1(\datamem.data_ram[43][29] ),
    .A2(_06828_),
    .B1(_06789_),
    .B2(\datamem.data_ram[41][29] ),
    .C1(_06851_),
    .X(_07949_));
 sky130_fd_sc_hd__o211a_1 _20659_ (.A1(\datamem.data_ram[45][29] ),
    .A2(_07037_),
    .B1(_07948_),
    .C1(_07949_),
    .X(_07950_));
 sky130_fd_sc_hd__o211a_1 _20660_ (.A1(\datamem.data_ram[47][29] ),
    .A2(_07020_),
    .B1(_07947_),
    .C1(_07950_),
    .X(_07951_));
 sky130_fd_sc_hd__o22a_1 _20661_ (.A1(\datamem.data_ram[62][29] ),
    .A2(_06627_),
    .B1(_06805_),
    .B2(\datamem.data_ram[60][29] ),
    .X(_07952_));
 sky130_fd_sc_hd__o22a_1 _20662_ (.A1(\datamem.data_ram[61][29] ),
    .A2(_06661_),
    .B1(_06811_),
    .B2(\datamem.data_ram[56][29] ),
    .X(_07953_));
 sky130_fd_sc_hd__o221a_1 _20663_ (.A1(\datamem.data_ram[58][29] ),
    .A2(_06802_),
    .B1(_06812_),
    .B2(\datamem.data_ram[59][29] ),
    .C1(_06599_),
    .X(_07954_));
 sky130_fd_sc_hd__o211a_1 _20664_ (.A1(\datamem.data_ram[57][29] ),
    .A2(_06789_),
    .B1(_07953_),
    .C1(_07954_),
    .X(_07955_));
 sky130_fd_sc_hd__o211a_1 _20665_ (.A1(\datamem.data_ram[63][29] ),
    .A2(_06784_),
    .B1(_07952_),
    .C1(_07955_),
    .X(_07956_));
 sky130_fd_sc_hd__o22a_1 _20666_ (.A1(\datamem.data_ram[54][29] ),
    .A2(_06718_),
    .B1(_06670_),
    .B2(\datamem.data_ram[55][29] ),
    .X(_07957_));
 sky130_fd_sc_hd__o22a_1 _20667_ (.A1(\datamem.data_ram[51][29] ),
    .A2(_06729_),
    .B1(_06684_),
    .B2(\datamem.data_ram[52][29] ),
    .X(_07958_));
 sky130_fd_sc_hd__o221a_1 _20668_ (.A1(\datamem.data_ram[48][29] ),
    .A2(_06811_),
    .B1(_06655_),
    .B2(\datamem.data_ram[49][29] ),
    .C1(_07958_),
    .X(_07959_));
 sky130_fd_sc_hd__o211a_1 _20669_ (.A1(\datamem.data_ram[53][29] ),
    .A2(_06823_),
    .B1(_06733_),
    .C1(_07959_),
    .X(_07960_));
 sky130_fd_sc_hd__o211a_1 _20670_ (.A1(\datamem.data_ram[50][29] ),
    .A2(_06804_),
    .B1(_07957_),
    .C1(_07960_),
    .X(_07961_));
 sky130_fd_sc_hd__o31a_1 _20671_ (.A1(_06752_),
    .A2(_07956_),
    .A3(_07961_),
    .B1(_06594_),
    .X(_07962_));
 sky130_fd_sc_hd__o31a_1 _20672_ (.A1(_06715_),
    .A2(_07946_),
    .A3(_07951_),
    .B1(_07962_),
    .X(_07963_));
 sky130_fd_sc_hd__a211oi_2 _20673_ (.A1(_06596_),
    .A2(_07930_),
    .B1(_07941_),
    .C1(_07963_),
    .Y(_07964_));
 sky130_fd_sc_hd__mux2_1 _20674_ (.A0(_07920_),
    .A1(net36),
    .S(_06911_),
    .X(_07965_));
 sky130_fd_sc_hd__a22o_1 _20675_ (.A1(\datamem.data_ram[46][5] ),
    .A2(_06978_),
    .B1(_06948_),
    .B2(\datamem.data_ram[41][5] ),
    .X(_07966_));
 sky130_fd_sc_hd__a221o_1 _20676_ (.A1(\datamem.data_ram[40][5] ),
    .A2(_07138_),
    .B1(_06977_),
    .B2(\datamem.data_ram[44][5] ),
    .C1(_07966_),
    .X(_07967_));
 sky130_fd_sc_hd__a22o_1 _20677_ (.A1(\datamem.data_ram[42][5] ),
    .A2(_06989_),
    .B1(_06921_),
    .B2(\datamem.data_ram[45][5] ),
    .X(_07968_));
 sky130_fd_sc_hd__a221o_1 _20678_ (.A1(\datamem.data_ram[43][5] ),
    .A2(_07137_),
    .B1(_07125_),
    .B2(\datamem.data_ram[47][5] ),
    .C1(_07968_),
    .X(_07969_));
 sky130_fd_sc_hd__or3_1 _20679_ (.A(_07131_),
    .B(_07967_),
    .C(_07969_),
    .X(_07970_));
 sky130_fd_sc_hd__a22o_1 _20680_ (.A1(\datamem.data_ram[37][5] ),
    .A2(_07132_),
    .B1(_07123_),
    .B2(\datamem.data_ram[36][5] ),
    .X(_07971_));
 sky130_fd_sc_hd__a22o_1 _20681_ (.A1(\datamem.data_ram[38][5] ),
    .A2(_06978_),
    .B1(_06949_),
    .B2(\datamem.data_ram[33][5] ),
    .X(_07972_));
 sky130_fd_sc_hd__a221o_1 _20682_ (.A1(\datamem.data_ram[35][5] ),
    .A2(_06943_),
    .B1(_06993_),
    .B2(\datamem.data_ram[39][5] ),
    .C1(_06602_),
    .X(_07973_));
 sky130_fd_sc_hd__a211o_1 _20683_ (.A1(\datamem.data_ram[32][5] ),
    .A2(_07122_),
    .B1(_07972_),
    .C1(_07973_),
    .X(_07974_));
 sky130_fd_sc_hd__a211o_1 _20684_ (.A1(\datamem.data_ram[34][5] ),
    .A2(_07136_),
    .B1(_07971_),
    .C1(_07974_),
    .X(_07975_));
 sky130_fd_sc_hd__a221o_1 _20685_ (.A1(\datamem.data_ram[53][5] ),
    .A2(_06970_),
    .B1(_07137_),
    .B2(\datamem.data_ram[51][5] ),
    .C1(_06603_),
    .X(_07976_));
 sky130_fd_sc_hd__a22o_1 _20686_ (.A1(\datamem.data_ram[52][5] ),
    .A2(_06955_),
    .B1(_06948_),
    .B2(\datamem.data_ram[49][5] ),
    .X(_07977_));
 sky130_fd_sc_hd__a21o_1 _20687_ (.A1(\datamem.data_ram[55][5] ),
    .A2(_06993_),
    .B1(_07977_),
    .X(_07978_));
 sky130_fd_sc_hd__a22o_1 _20688_ (.A1(\datamem.data_ram[54][5] ),
    .A2(_06978_),
    .B1(_07000_),
    .B2(\datamem.data_ram[50][5] ),
    .X(_07979_));
 sky130_fd_sc_hd__a211o_1 _20689_ (.A1(\datamem.data_ram[48][5] ),
    .A2(_07122_),
    .B1(_07978_),
    .C1(_07979_),
    .X(_07980_));
 sky130_fd_sc_hd__a22o_1 _20690_ (.A1(\datamem.data_ram[58][5] ),
    .A2(_07000_),
    .B1(_07138_),
    .B2(\datamem.data_ram[56][5] ),
    .X(_07981_));
 sky130_fd_sc_hd__a22o_1 _20691_ (.A1(\datamem.data_ram[61][5] ),
    .A2(_06969_),
    .B1(_06955_),
    .B2(\datamem.data_ram[60][5] ),
    .X(_07982_));
 sky130_fd_sc_hd__a221o_1 _20692_ (.A1(\datamem.data_ram[59][5] ),
    .A2(_06961_),
    .B1(_06926_),
    .B2(\datamem.data_ram[63][5] ),
    .C1(_06679_),
    .X(_07983_));
 sky130_fd_sc_hd__a211o_1 _20693_ (.A1(\datamem.data_ram[57][5] ),
    .A2(_06949_),
    .B1(_07982_),
    .C1(_07983_),
    .X(_07984_));
 sky130_fd_sc_hd__a211o_1 _20694_ (.A1(\datamem.data_ram[62][5] ),
    .A2(_07159_),
    .B1(_07981_),
    .C1(_07984_),
    .X(_07985_));
 sky130_fd_sc_hd__o211a_1 _20695_ (.A1(_07976_),
    .A2(_07980_),
    .B1(_07071_),
    .C1(_07985_),
    .X(_07986_));
 sky130_fd_sc_hd__a31o_1 _20696_ (.A1(_06916_),
    .A2(_07970_),
    .A3(_07975_),
    .B1(_07986_),
    .X(_07987_));
 sky130_fd_sc_hd__a22o_1 _20697_ (.A1(\datamem.data_ram[2][5] ),
    .A2(_07000_),
    .B1(_06927_),
    .B2(\datamem.data_ram[7][5] ),
    .X(_07988_));
 sky130_fd_sc_hd__a22o_1 _20698_ (.A1(\datamem.data_ram[5][5] ),
    .A2(_06969_),
    .B1(_06955_),
    .B2(\datamem.data_ram[4][5] ),
    .X(_07989_));
 sky130_fd_sc_hd__a221o_1 _20699_ (.A1(\datamem.data_ram[0][5] ),
    .A2(_06937_),
    .B1(_06961_),
    .B2(\datamem.data_ram[3][5] ),
    .C1(_06742_),
    .X(_07990_));
 sky130_fd_sc_hd__a211o_1 _20700_ (.A1(\datamem.data_ram[6][5] ),
    .A2(_07127_),
    .B1(_07989_),
    .C1(_07990_),
    .X(_07991_));
 sky130_fd_sc_hd__a211o_1 _20701_ (.A1(\datamem.data_ram[1][5] ),
    .A2(_07133_),
    .B1(_07988_),
    .C1(_07991_),
    .X(_07992_));
 sky130_fd_sc_hd__a22o_1 _20702_ (.A1(\datamem.data_ram[14][5] ),
    .A2(_07127_),
    .B1(_07000_),
    .B2(\datamem.data_ram[10][5] ),
    .X(_07993_));
 sky130_fd_sc_hd__a22o_1 _20703_ (.A1(\datamem.data_ram[12][5] ),
    .A2(_06955_),
    .B1(_06958_),
    .B2(\datamem.data_ram[9][5] ),
    .X(_07994_));
 sky130_fd_sc_hd__a221o_1 _20704_ (.A1(\datamem.data_ram[8][5] ),
    .A2(_06937_),
    .B1(_06925_),
    .B2(\datamem.data_ram[15][5] ),
    .C1(_06679_),
    .X(_07995_));
 sky130_fd_sc_hd__a211o_1 _20705_ (.A1(\datamem.data_ram[13][5] ),
    .A2(_06921_),
    .B1(_07994_),
    .C1(_07995_),
    .X(_07996_));
 sky130_fd_sc_hd__a211o_1 _20706_ (.A1(\datamem.data_ram[11][5] ),
    .A2(_07137_),
    .B1(_07993_),
    .C1(_07996_),
    .X(_07997_));
 sky130_fd_sc_hd__a21o_1 _20707_ (.A1(_07992_),
    .A2(_07997_),
    .B1(_07154_),
    .X(_07998_));
 sky130_fd_sc_hd__a22o_1 _20708_ (.A1(\datamem.data_ram[24][5] ),
    .A2(_07138_),
    .B1(_06949_),
    .B2(\datamem.data_ram[25][5] ),
    .X(_07999_));
 sky130_fd_sc_hd__a22o_1 _20709_ (.A1(\datamem.data_ram[26][5] ),
    .A2(_06932_),
    .B1(_06969_),
    .B2(\datamem.data_ram[29][5] ),
    .X(_08000_));
 sky130_fd_sc_hd__a221o_1 _20710_ (.A1(\datamem.data_ram[30][5] ),
    .A2(_06952_),
    .B1(_06925_),
    .B2(\datamem.data_ram[31][5] ),
    .C1(_06679_),
    .X(_08001_));
 sky130_fd_sc_hd__a211o_1 _20711_ (.A1(\datamem.data_ram[27][5] ),
    .A2(_06966_),
    .B1(_08000_),
    .C1(_08001_),
    .X(_08002_));
 sky130_fd_sc_hd__a211o_1 _20712_ (.A1(\datamem.data_ram[28][5] ),
    .A2(_07123_),
    .B1(_07999_),
    .C1(_08002_),
    .X(_08003_));
 sky130_fd_sc_hd__a22o_1 _20713_ (.A1(\datamem.data_ram[16][5] ),
    .A2(_06990_),
    .B1(_06976_),
    .B2(\datamem.data_ram[20][5] ),
    .X(_08004_));
 sky130_fd_sc_hd__a22o_1 _20714_ (.A1(\datamem.data_ram[18][5] ),
    .A2(_06932_),
    .B1(_06958_),
    .B2(\datamem.data_ram[17][5] ),
    .X(_08005_));
 sky130_fd_sc_hd__a221o_1 _20715_ (.A1(\datamem.data_ram[22][5] ),
    .A2(_06952_),
    .B1(_06969_),
    .B2(\datamem.data_ram[21][5] ),
    .C1(_06810_),
    .X(_08006_));
 sky130_fd_sc_hd__a211o_1 _20716_ (.A1(\datamem.data_ram[23][5] ),
    .A2(_06927_),
    .B1(_08005_),
    .C1(_08006_),
    .X(_08007_));
 sky130_fd_sc_hd__a211o_1 _20717_ (.A1(\datamem.data_ram[19][5] ),
    .A2(_07137_),
    .B1(_08004_),
    .C1(_08007_),
    .X(_08008_));
 sky130_fd_sc_hd__a21o_1 _20718_ (.A1(_08003_),
    .A2(_08008_),
    .B1(_07177_),
    .X(_08009_));
 sky130_fd_sc_hd__and3_1 _20719_ (.A(_06988_),
    .B(_07998_),
    .C(_08009_),
    .X(_08010_));
 sky130_fd_sc_hd__o21ai_2 _20720_ (.A1(_06985_),
    .A2(_07987_),
    .B1(_08010_),
    .Y(_08011_));
 sky130_fd_sc_hd__o31a_1 _20721_ (.A1(_06583_),
    .A2(_06588_),
    .A3(_07965_),
    .B1(_08011_),
    .X(_08012_));
 sky130_fd_sc_hd__o21ai_1 _20722_ (.A1(_07227_),
    .A2(_07857_),
    .B1(_08012_),
    .Y(_04442_));
 sky130_fd_sc_hd__mux2_1 _20723_ (.A0(\datamem.data_ram[16][6] ),
    .A1(\datamem.data_ram[17][6] ),
    .S(_07837_),
    .X(_08013_));
 sky130_fd_sc_hd__a221o_1 _20724_ (.A1(_07823_),
    .A2(\datamem.data_ram[18][6] ),
    .B1(\datamem.data_ram[19][6] ),
    .B2(_07837_),
    .C1(_07840_),
    .X(_08014_));
 sky130_fd_sc_hd__o211a_1 _20725_ (.A1(_07822_),
    .A2(_08013_),
    .B1(_08014_),
    .C1(_07845_),
    .X(_08015_));
 sky130_fd_sc_hd__a221o_1 _20726_ (.A1(\datamem.data_ram[22][6] ),
    .A2(_07159_),
    .B1(_06927_),
    .B2(\datamem.data_ram[23][6] ),
    .C1(_07081_),
    .X(_08016_));
 sky130_fd_sc_hd__a221o_1 _20727_ (.A1(\datamem.data_ram[21][6] ),
    .A2(_07132_),
    .B1(_07123_),
    .B2(\datamem.data_ram[20][6] ),
    .C1(_08016_),
    .X(_08017_));
 sky130_fd_sc_hd__mux2_1 _20728_ (.A0(\datamem.data_ram[30][6] ),
    .A1(\datamem.data_ram[31][6] ),
    .S(_07837_),
    .X(_08018_));
 sky130_fd_sc_hd__mux2_1 _20729_ (.A0(\datamem.data_ram[28][6] ),
    .A1(\datamem.data_ram[29][6] ),
    .S(_07829_),
    .X(_08019_));
 sky130_fd_sc_hd__mux4_1 _20730_ (.A0(\datamem.data_ram[24][6] ),
    .A1(\datamem.data_ram[25][6] ),
    .A2(\datamem.data_ram[26][6] ),
    .A3(\datamem.data_ram[27][6] ),
    .S0(_07836_),
    .S1(_07822_),
    .X(_08020_));
 sky130_fd_sc_hd__a22o_1 _20731_ (.A1(_06615_),
    .A2(_08019_),
    .B1(_08020_),
    .B2(_07845_),
    .X(_08021_));
 sky130_fd_sc_hd__a211o_1 _20732_ (.A1(_06623_),
    .A2(_08018_),
    .B1(_08021_),
    .C1(_07131_),
    .X(_08022_));
 sky130_fd_sc_hd__o211a_1 _20733_ (.A1(_08015_),
    .A2(_08017_),
    .B1(_06797_),
    .C1(_08022_),
    .X(_08023_));
 sky130_fd_sc_hd__mux2_1 _20734_ (.A0(\datamem.data_ram[34][6] ),
    .A1(\datamem.data_ram[35][6] ),
    .S(_07837_),
    .X(_08024_));
 sky130_fd_sc_hd__mux2_1 _20735_ (.A0(\datamem.data_ram[38][6] ),
    .A1(\datamem.data_ram[39][6] ),
    .S(_07828_),
    .X(_08025_));
 sky130_fd_sc_hd__mux2_1 _20736_ (.A0(\datamem.data_ram[36][6] ),
    .A1(\datamem.data_ram[37][6] ),
    .S(_07828_),
    .X(_08026_));
 sky130_fd_sc_hd__mux2_1 _20737_ (.A0(_08025_),
    .A1(_08026_),
    .S(_07840_),
    .X(_08027_));
 sky130_fd_sc_hd__a22o_1 _20738_ (.A1(\datamem.data_ram[32][6] ),
    .A2(_07122_),
    .B1(_08027_),
    .B2(_07868_),
    .X(_08028_));
 sky130_fd_sc_hd__a221o_1 _20739_ (.A1(\datamem.data_ram[33][6] ),
    .A2(_06997_),
    .B1(_08024_),
    .B2(_07636_),
    .C1(_08028_),
    .X(_08029_));
 sky130_fd_sc_hd__a221o_1 _20740_ (.A1(\datamem.data_ram[42][6] ),
    .A2(_07000_),
    .B1(_07137_),
    .B2(\datamem.data_ram[43][6] ),
    .C1(_06777_),
    .X(_08030_));
 sky130_fd_sc_hd__a31o_1 _20741_ (.A1(\datamem.data_ram[41][6] ),
    .A2(_07839_),
    .A3(_07845_),
    .B1(_07832_),
    .X(_08031_));
 sky130_fd_sc_hd__a221o_1 _20742_ (.A1(\datamem.data_ram[47][6] ),
    .A2(_06623_),
    .B1(_06615_),
    .B2(\datamem.data_ram[45][6] ),
    .C1(_08031_),
    .X(_08032_));
 sky130_fd_sc_hd__a31o_1 _20743_ (.A1(\rvcpu.dp.plem.ALUResultM[4] ),
    .A2(\datamem.data_ram[46][6] ),
    .A3(_07821_),
    .B1(_07836_),
    .X(_08033_));
 sky130_fd_sc_hd__a221o_1 _20744_ (.A1(\datamem.data_ram[44][6] ),
    .A2(_06615_),
    .B1(_06642_),
    .B2(\datamem.data_ram[40][6] ),
    .C1(_08033_),
    .X(_08034_));
 sky130_fd_sc_hd__and2_1 _20745_ (.A(_08032_),
    .B(_08034_),
    .X(_08035_));
 sky130_fd_sc_hd__or2_1 _20746_ (.A(_08030_),
    .B(_08035_),
    .X(_08036_));
 sky130_fd_sc_hd__o211a_1 _20747_ (.A1(_06604_),
    .A2(_08029_),
    .B1(_08036_),
    .C1(_07858_),
    .X(_08037_));
 sky130_fd_sc_hd__or2_1 _20748_ (.A(\datamem.data_ram[8][6] ),
    .B(_07829_),
    .X(_08038_));
 sky130_fd_sc_hd__or2_1 _20749_ (.A(\datamem.data_ram[9][6] ),
    .B(_07833_),
    .X(_08039_));
 sky130_fd_sc_hd__mux2_1 _20750_ (.A0(\datamem.data_ram[12][6] ),
    .A1(\datamem.data_ram[13][6] ),
    .S(_07836_),
    .X(_08040_));
 sky130_fd_sc_hd__a32o_1 _20751_ (.A1(_06642_),
    .A2(_08038_),
    .A3(_08039_),
    .B1(_08040_),
    .B2(_06615_),
    .X(_08041_));
 sky130_fd_sc_hd__or2_1 _20752_ (.A(\datamem.data_ram[14][6] ),
    .B(_07829_),
    .X(_08042_));
 sky130_fd_sc_hd__o211a_1 _20753_ (.A1(\datamem.data_ram[15][6] ),
    .A2(_07833_),
    .B1(_08042_),
    .C1(_06623_),
    .X(_08043_));
 sky130_fd_sc_hd__o221a_1 _20754_ (.A1(_07635_),
    .A2(\datamem.data_ram[10][6] ),
    .B1(\datamem.data_ram[11][6] ),
    .B2(_07833_),
    .C1(_07636_),
    .X(_08044_));
 sky130_fd_sc_hd__or3_2 _20755_ (.A(_08041_),
    .B(_08043_),
    .C(_08044_),
    .X(_08045_));
 sky130_fd_sc_hd__mux2_1 _20756_ (.A0(\datamem.data_ram[6][6] ),
    .A1(\datamem.data_ram[7][6] ),
    .S(_07828_),
    .X(_08046_));
 sky130_fd_sc_hd__mux2_1 _20757_ (.A0(\datamem.data_ram[4][6] ),
    .A1(\datamem.data_ram[5][6] ),
    .S(_07828_),
    .X(_08047_));
 sky130_fd_sc_hd__mux2_1 _20758_ (.A0(_08046_),
    .A1(_08047_),
    .S(_07840_),
    .X(_08048_));
 sky130_fd_sc_hd__or2_1 _20759_ (.A(\datamem.data_ram[3][6] ),
    .B(_07832_),
    .X(_08049_));
 sky130_fd_sc_hd__o211a_1 _20760_ (.A1(\datamem.data_ram[2][6] ),
    .A2(_07837_),
    .B1(_08049_),
    .C1(_07636_),
    .X(_08050_));
 sky130_fd_sc_hd__a221o_1 _20761_ (.A1(\datamem.data_ram[0][6] ),
    .A2(_07122_),
    .B1(_08048_),
    .B2(_07868_),
    .C1(_08050_),
    .X(_08051_));
 sky130_fd_sc_hd__a211o_1 _20762_ (.A1(\datamem.data_ram[1][6] ),
    .A2(_06997_),
    .B1(_08051_),
    .C1(_06604_),
    .X(_08052_));
 sky130_fd_sc_hd__o211a_1 _20763_ (.A1(_07131_),
    .A2(_08045_),
    .B1(_08052_),
    .C1(_06596_),
    .X(_08053_));
 sky130_fd_sc_hd__a22o_1 _20764_ (.A1(\datamem.data_ram[50][6] ),
    .A2(_07000_),
    .B1(_07133_),
    .B2(\datamem.data_ram[49][6] ),
    .X(_08054_));
 sky130_fd_sc_hd__a22o_1 _20765_ (.A1(\datamem.data_ram[54][6] ),
    .A2(_07159_),
    .B1(_07137_),
    .B2(\datamem.data_ram[51][6] ),
    .X(_08055_));
 sky130_fd_sc_hd__a22o_1 _20766_ (.A1(\datamem.data_ram[48][6] ),
    .A2(_07138_),
    .B1(_07123_),
    .B2(\datamem.data_ram[52][6] ),
    .X(_08056_));
 sky130_fd_sc_hd__a22o_1 _20767_ (.A1(\datamem.data_ram[53][6] ),
    .A2(_06970_),
    .B1(_07125_),
    .B2(\datamem.data_ram[55][6] ),
    .X(_08057_));
 sky130_fd_sc_hd__or4_1 _20768_ (.A(_08054_),
    .B(_08055_),
    .C(_08056_),
    .D(_08057_),
    .X(_08058_));
 sky130_fd_sc_hd__nor2_1 _20769_ (.A(_06604_),
    .B(_07872_),
    .Y(_08059_));
 sky130_fd_sc_hd__mux2_1 _20770_ (.A0(\datamem.data_ram[60][6] ),
    .A1(\datamem.data_ram[61][6] ),
    .S(_07829_),
    .X(_08060_));
 sky130_fd_sc_hd__and2_1 _20771_ (.A(_07635_),
    .B(\datamem.data_ram[63][6] ),
    .X(_08061_));
 sky130_fd_sc_hd__a211o_1 _20772_ (.A1(\datamem.data_ram[62][6] ),
    .A2(_07833_),
    .B1(_08061_),
    .C1(_07840_),
    .X(_08062_));
 sky130_fd_sc_hd__o211a_1 _20773_ (.A1(_07822_),
    .A2(_08060_),
    .B1(_08062_),
    .C1(_07868_),
    .X(_08063_));
 sky130_fd_sc_hd__a22o_1 _20774_ (.A1(\datamem.data_ram[56][6] ),
    .A2(_07122_),
    .B1(_07133_),
    .B2(\datamem.data_ram[57][6] ),
    .X(_08064_));
 sky130_fd_sc_hd__a22o_1 _20775_ (.A1(\datamem.data_ram[58][6] ),
    .A2(_07136_),
    .B1(_07137_),
    .B2(\datamem.data_ram[59][6] ),
    .X(_08065_));
 sky130_fd_sc_hd__nor2_1 _20776_ (.A(_06681_),
    .B(_07872_),
    .Y(_08066_));
 sky130_fd_sc_hd__o31a_1 _20777_ (.A1(_08063_),
    .A2(_08064_),
    .A3(_08065_),
    .B1(_08066_),
    .X(_08067_));
 sky130_fd_sc_hd__a21o_1 _20778_ (.A1(_08058_),
    .A2(_08059_),
    .B1(_08067_),
    .X(_08068_));
 sky130_fd_sc_hd__or4_2 _20779_ (.A(_08023_),
    .B(_08037_),
    .C(_08053_),
    .D(_08068_),
    .X(_08069_));
 sky130_fd_sc_hd__mux2_1 _20780_ (.A0(\datamem.data_ram[4][30] ),
    .A1(\datamem.data_ram[5][30] ),
    .S(_07849_),
    .X(_08070_));
 sky130_fd_sc_hd__mux2_1 _20781_ (.A0(\datamem.data_ram[6][30] ),
    .A1(\datamem.data_ram[7][30] ),
    .S(_07836_),
    .X(_08071_));
 sky130_fd_sc_hd__a221o_1 _20782_ (.A1(_07840_),
    .A2(_08070_),
    .B1(_08071_),
    .B2(\rvcpu.dp.plem.ALUResultM[3] ),
    .C1(_07845_),
    .X(_08072_));
 sky130_fd_sc_hd__o22a_1 _20783_ (.A1(\datamem.data_ram[0][30] ),
    .A2(_06779_),
    .B1(_06783_),
    .B2(\datamem.data_ram[1][30] ),
    .X(_08073_));
 sky130_fd_sc_hd__o221a_1 _20784_ (.A1(\datamem.data_ram[2][30] ),
    .A2(_07023_),
    .B1(_06739_),
    .B2(\datamem.data_ram[3][30] ),
    .C1(_08073_),
    .X(_08074_));
 sky130_fd_sc_hd__or2_1 _20785_ (.A(\datamem.data_ram[17][30] ),
    .B(_07832_),
    .X(_08075_));
 sky130_fd_sc_hd__o21a_1 _20786_ (.A1(\datamem.data_ram[16][30] ),
    .A2(_07828_),
    .B1(_07839_),
    .X(_08076_));
 sky130_fd_sc_hd__mux2_1 _20787_ (.A0(\datamem.data_ram[18][30] ),
    .A1(\datamem.data_ram[19][30] ),
    .S(_07835_),
    .X(_08077_));
 sky130_fd_sc_hd__a221o_1 _20788_ (.A1(_08075_),
    .A2(_08076_),
    .B1(_08077_),
    .B2(_07822_),
    .C1(_07868_),
    .X(_08078_));
 sky130_fd_sc_hd__o221a_1 _20789_ (.A1(\datamem.data_ram[23][30] ),
    .A2(_06761_),
    .B1(_07024_),
    .B2(\datamem.data_ram[20][30] ),
    .C1(_06714_),
    .X(_08079_));
 sky130_fd_sc_hd__o22a_1 _20790_ (.A1(\datamem.data_ram[22][30] ),
    .A2(_06629_),
    .B1(_06703_),
    .B2(\datamem.data_ram[21][30] ),
    .X(_08080_));
 sky130_fd_sc_hd__a31o_1 _20791_ (.A1(_08078_),
    .A2(_08079_),
    .A3(_08080_),
    .B1(_06712_),
    .X(_08081_));
 sky130_fd_sc_hd__a31o_1 _20792_ (.A1(_06753_),
    .A2(_08072_),
    .A3(_08074_),
    .B1(_08081_),
    .X(_08082_));
 sky130_fd_sc_hd__mux2_1 _20793_ (.A0(\datamem.data_ram[34][30] ),
    .A1(\datamem.data_ram[35][30] ),
    .S(_07849_),
    .X(_08083_));
 sky130_fd_sc_hd__a221o_1 _20794_ (.A1(\datamem.data_ram[32][30] ),
    .A2(_06990_),
    .B1(_08083_),
    .B2(_07636_),
    .C1(_07903_),
    .X(_08084_));
 sky130_fd_sc_hd__mux2_1 _20795_ (.A0(\datamem.data_ram[36][30] ),
    .A1(\datamem.data_ram[37][30] ),
    .S(_07835_),
    .X(_08085_));
 sky130_fd_sc_hd__mux2_1 _20796_ (.A0(\datamem.data_ram[38][30] ),
    .A1(\datamem.data_ram[39][30] ),
    .S(_07835_),
    .X(_08086_));
 sky130_fd_sc_hd__mux2_1 _20797_ (.A0(_08085_),
    .A1(_08086_),
    .S(_07822_),
    .X(_08087_));
 sky130_fd_sc_hd__a22o_1 _20798_ (.A1(\datamem.data_ram[33][30] ),
    .A2(_06949_),
    .B1(_08087_),
    .B2(\rvcpu.dp.plem.ALUResultM[4] ),
    .X(_08088_));
 sky130_fd_sc_hd__and2_1 _20799_ (.A(\datamem.data_ram[50][30] ),
    .B(_07831_),
    .X(_08089_));
 sky130_fd_sc_hd__a211o_1 _20800_ (.A1(\datamem.data_ram[51][30] ),
    .A2(_07849_),
    .B1(_08089_),
    .C1(_07851_),
    .X(_08090_));
 sky130_fd_sc_hd__o221a_1 _20801_ (.A1(\datamem.data_ram[54][30] ),
    .A2(_06629_),
    .B1(_06783_),
    .B2(\datamem.data_ram[49][30] ),
    .C1(_08090_),
    .X(_08091_));
 sky130_fd_sc_hd__o22a_1 _20802_ (.A1(\datamem.data_ram[53][30] ),
    .A2(_06663_),
    .B1(_07230_),
    .B2(\datamem.data_ram[52][30] ),
    .X(_08092_));
 sky130_fd_sc_hd__o221a_1 _20803_ (.A1(\datamem.data_ram[48][30] ),
    .A2(_06779_),
    .B1(_06707_),
    .B2(\datamem.data_ram[55][30] ),
    .C1(_08092_),
    .X(_08093_));
 sky130_fd_sc_hd__a21o_1 _20804_ (.A1(_08091_),
    .A2(_08093_),
    .B1(_07872_),
    .X(_08094_));
 sky130_fd_sc_hd__o211a_1 _20805_ (.A1(_08084_),
    .A2(_08088_),
    .B1(_06681_),
    .C1(_08094_),
    .X(_08095_));
 sky130_fd_sc_hd__mux2_1 _20806_ (.A0(\datamem.data_ram[42][30] ),
    .A1(\datamem.data_ram[43][30] ),
    .S(_07835_),
    .X(_08096_));
 sky130_fd_sc_hd__mux2_1 _20807_ (.A0(\datamem.data_ram[44][30] ),
    .A1(\datamem.data_ram[45][30] ),
    .S(_07826_),
    .X(_08097_));
 sky130_fd_sc_hd__mux2_1 _20808_ (.A0(\datamem.data_ram[46][30] ),
    .A1(\datamem.data_ram[47][30] ),
    .S(_07826_),
    .X(_08098_));
 sky130_fd_sc_hd__mux2_1 _20809_ (.A0(_08097_),
    .A1(_08098_),
    .S(_07820_),
    .X(_08099_));
 sky130_fd_sc_hd__a22o_1 _20810_ (.A1(\datamem.data_ram[41][30] ),
    .A2(_06947_),
    .B1(_08099_),
    .B2(_07867_),
    .X(_08100_));
 sky130_fd_sc_hd__a221o_1 _20811_ (.A1(\datamem.data_ram[40][30] ),
    .A2(_06973_),
    .B1(_08096_),
    .B2(_07636_),
    .C1(_08100_),
    .X(_08101_));
 sky130_fd_sc_hd__o22a_1 _20812_ (.A1(\datamem.data_ram[59][30] ),
    .A2(_06940_),
    .B1(_06934_),
    .B2(\datamem.data_ram[57][30] ),
    .X(_08102_));
 sky130_fd_sc_hd__o221a_1 _20813_ (.A1(\datamem.data_ram[63][30] ),
    .A2(_07860_),
    .B1(_07862_),
    .B2(\datamem.data_ram[61][30] ),
    .C1(_08102_),
    .X(_08103_));
 sky130_fd_sc_hd__or2_1 _20814_ (.A(\datamem.data_ram[56][30] ),
    .B(_06934_),
    .X(_08104_));
 sky130_fd_sc_hd__o221a_1 _20815_ (.A1(\datamem.data_ram[62][30] ),
    .A2(_07859_),
    .B1(_07862_),
    .B2(\datamem.data_ram[60][30] ),
    .C1(_08104_),
    .X(_08105_));
 sky130_fd_sc_hd__o211a_1 _20816_ (.A1(\datamem.data_ram[58][30] ),
    .A2(_06940_),
    .B1(_07832_),
    .C1(_08105_),
    .X(_08106_));
 sky130_fd_sc_hd__a211o_1 _20817_ (.A1(_07829_),
    .A2(_08103_),
    .B1(_08106_),
    .C1(_06751_),
    .X(_08107_));
 sky130_fd_sc_hd__o211a_1 _20818_ (.A1(_06715_),
    .A2(_08101_),
    .B1(_08107_),
    .C1(_06712_),
    .X(_08108_));
 sky130_fd_sc_hd__o22a_1 _20819_ (.A1(\datamem.data_ram[31][30] ),
    .A2(_07860_),
    .B1(_06934_),
    .B2(\datamem.data_ram[25][30] ),
    .X(_08109_));
 sky130_fd_sc_hd__o22a_1 _20820_ (.A1(\datamem.data_ram[27][30] ),
    .A2(_06940_),
    .B1(_07863_),
    .B2(\datamem.data_ram[29][30] ),
    .X(_08110_));
 sky130_fd_sc_hd__a21o_1 _20821_ (.A1(_08109_),
    .A2(_08110_),
    .B1(_07833_),
    .X(_08111_));
 sky130_fd_sc_hd__o22a_1 _20822_ (.A1(\datamem.data_ram[30][30] ),
    .A2(_07860_),
    .B1(_07863_),
    .B2(\datamem.data_ram[28][30] ),
    .X(_08112_));
 sky130_fd_sc_hd__o22a_1 _20823_ (.A1(\datamem.data_ram[26][30] ),
    .A2(_06940_),
    .B1(_06934_),
    .B2(\datamem.data_ram[24][30] ),
    .X(_08113_));
 sky130_fd_sc_hd__a21o_1 _20824_ (.A1(_08112_),
    .A2(_08113_),
    .B1(_07837_),
    .X(_08114_));
 sky130_fd_sc_hd__mux2_1 _20825_ (.A0(\datamem.data_ram[10][30] ),
    .A1(\datamem.data_ram[11][30] ),
    .S(_07827_),
    .X(_08115_));
 sky130_fd_sc_hd__o22a_1 _20826_ (.A1(\datamem.data_ram[13][30] ),
    .A2(_06663_),
    .B1(_08115_),
    .B2(_07851_),
    .X(_08116_));
 sky130_fd_sc_hd__o22a_1 _20827_ (.A1(\datamem.data_ram[14][30] ),
    .A2(_07085_),
    .B1(_06618_),
    .B2(\datamem.data_ram[12][30] ),
    .X(_08117_));
 sky130_fd_sc_hd__o211a_1 _20828_ (.A1(\datamem.data_ram[15][30] ),
    .A2(_06706_),
    .B1(_06595_),
    .C1(_08117_),
    .X(_08118_));
 sky130_fd_sc_hd__o22a_1 _20829_ (.A1(\datamem.data_ram[8][30] ),
    .A2(_06647_),
    .B1(_06782_),
    .B2(\datamem.data_ram[9][30] ),
    .X(_08119_));
 sky130_fd_sc_hd__and3_1 _20830_ (.A(_08116_),
    .B(_08118_),
    .C(_08119_),
    .X(_08120_));
 sky130_fd_sc_hd__a31o_1 _20831_ (.A1(_06796_),
    .A2(_08111_),
    .A3(_08114_),
    .B1(_08120_),
    .X(_08121_));
 sky130_fd_sc_hd__o21a_1 _20832_ (.A1(_08108_),
    .A2(_08121_),
    .B1(_06604_),
    .X(_08122_));
 sky130_fd_sc_hd__a21oi_4 _20833_ (.A1(_08082_),
    .A2(_08095_),
    .B1(_08122_),
    .Y(_08123_));
 sky130_fd_sc_hd__clkbuf_8 _20834_ (.A(\rvcpu.dp.plem.ALUResultM[5] ),
    .X(_08124_));
 sky130_fd_sc_hd__nand2_8 _20835_ (.A(_08124_),
    .B(_06797_),
    .Y(_08125_));
 sky130_fd_sc_hd__mux2_1 _20836_ (.A0(\datamem.data_ram[28][14] ),
    .A1(\datamem.data_ram[29][14] ),
    .S(_07828_),
    .X(_08126_));
 sky130_fd_sc_hd__or2_1 _20837_ (.A(_07635_),
    .B(\datamem.data_ram[30][14] ),
    .X(_08127_));
 sky130_fd_sc_hd__o211a_1 _20838_ (.A1(\datamem.data_ram[31][14] ),
    .A2(_07832_),
    .B1(_08127_),
    .C1(_07821_),
    .X(_08128_));
 sky130_fd_sc_hd__a211o_1 _20839_ (.A1(_07840_),
    .A2(_08126_),
    .B1(_08128_),
    .C1(_07845_),
    .X(_08129_));
 sky130_fd_sc_hd__o221a_1 _20840_ (.A1(\datamem.data_ram[24][14] ),
    .A2(_06649_),
    .B1(_06701_),
    .B2(\datamem.data_ram[25][14] ),
    .C1(_08129_),
    .X(_08130_));
 sky130_fd_sc_hd__o221a_1 _20841_ (.A1(\datamem.data_ram[26][14] ),
    .A2(_07203_),
    .B1(_07077_),
    .B2(\datamem.data_ram[27][14] ),
    .C1(_08130_),
    .X(_08131_));
 sky130_fd_sc_hd__or2_1 _20842_ (.A(_08124_),
    .B(_07177_),
    .X(_08132_));
 sky130_fd_sc_hd__buf_6 _20843_ (.A(_08132_),
    .X(_08133_));
 sky130_fd_sc_hd__mux4_1 _20844_ (.A0(\datamem.data_ram[16][14] ),
    .A1(\datamem.data_ram[17][14] ),
    .A2(\datamem.data_ram[18][14] ),
    .A3(\datamem.data_ram[19][14] ),
    .S0(_07826_),
    .S1(_07821_),
    .X(_08134_));
 sky130_fd_sc_hd__or2_1 _20845_ (.A(_07867_),
    .B(_08134_),
    .X(_08135_));
 sky130_fd_sc_hd__o221a_1 _20846_ (.A1(\datamem.data_ram[22][14] ),
    .A2(_06629_),
    .B1(_06664_),
    .B2(\datamem.data_ram[21][14] ),
    .C1(_08135_),
    .X(_08136_));
 sky130_fd_sc_hd__o221a_1 _20847_ (.A1(\datamem.data_ram[23][14] ),
    .A2(_07021_),
    .B1(_06621_),
    .B2(\datamem.data_ram[20][14] ),
    .C1(_08136_),
    .X(_08137_));
 sky130_fd_sc_hd__mux2_1 _20848_ (.A0(\datamem.data_ram[4][14] ),
    .A1(\datamem.data_ram[5][14] ),
    .S(_07849_),
    .X(_08138_));
 sky130_fd_sc_hd__o22a_1 _20849_ (.A1(\datamem.data_ram[0][14] ),
    .A2(_06648_),
    .B1(_08138_),
    .B2(_07863_),
    .X(_08139_));
 sky130_fd_sc_hd__a221o_1 _20850_ (.A1(_07823_),
    .A2(\datamem.data_ram[6][14] ),
    .B1(\datamem.data_ram[7][14] ),
    .B2(_07849_),
    .C1(_07860_),
    .X(_08140_));
 sky130_fd_sc_hd__mux2_1 _20851_ (.A0(\datamem.data_ram[2][14] ),
    .A1(\datamem.data_ram[3][14] ),
    .S(_07835_),
    .X(_08141_));
 sky130_fd_sc_hd__or2_1 _20852_ (.A(_07851_),
    .B(_08141_),
    .X(_08142_));
 sky130_fd_sc_hd__o211a_1 _20853_ (.A1(\datamem.data_ram[1][14] ),
    .A2(_06658_),
    .B1(_08140_),
    .C1(_08142_),
    .X(_08143_));
 sky130_fd_sc_hd__nand2_8 _20854_ (.A(_06680_),
    .B(_06595_),
    .Y(_08144_));
 sky130_fd_sc_hd__a21o_1 _20855_ (.A1(_08139_),
    .A2(_08143_),
    .B1(_08144_),
    .X(_08145_));
 sky130_fd_sc_hd__a221o_1 _20856_ (.A1(_07635_),
    .A2(\datamem.data_ram[15][14] ),
    .B1(_07832_),
    .B2(\datamem.data_ram[14][14] ),
    .C1(_07845_),
    .X(_08146_));
 sky130_fd_sc_hd__a221o_1 _20857_ (.A1(_07823_),
    .A2(\datamem.data_ram[10][14] ),
    .B1(\datamem.data_ram[11][14] ),
    .B2(_07849_),
    .C1(_07867_),
    .X(_08147_));
 sky130_fd_sc_hd__a21o_1 _20858_ (.A1(_08146_),
    .A2(_08147_),
    .B1(_07840_),
    .X(_08148_));
 sky130_fd_sc_hd__a221o_1 _20859_ (.A1(_07635_),
    .A2(\datamem.data_ram[13][14] ),
    .B1(_07833_),
    .B2(\datamem.data_ram[12][14] ),
    .C1(_07863_),
    .X(_08149_));
 sky130_fd_sc_hd__o22a_1 _20860_ (.A1(\datamem.data_ram[8][14] ),
    .A2(_06648_),
    .B1(_06658_),
    .B2(\datamem.data_ram[9][14] ),
    .X(_08150_));
 sky130_fd_sc_hd__nand2_4 _20861_ (.A(_06967_),
    .B(_06595_),
    .Y(_08151_));
 sky130_fd_sc_hd__a31o_1 _20862_ (.A1(_08148_),
    .A2(_08149_),
    .A3(_08150_),
    .B1(_08151_),
    .X(_08152_));
 sky130_fd_sc_hd__o211a_1 _20863_ (.A1(_08133_),
    .A2(_08137_),
    .B1(_08145_),
    .C1(_08152_),
    .X(_08153_));
 sky130_fd_sc_hd__o22a_1 _20864_ (.A1(\datamem.data_ram[36][14] ),
    .A2(_07862_),
    .B1(_06934_),
    .B2(\datamem.data_ram[32][14] ),
    .X(_08154_));
 sky130_fd_sc_hd__o221a_1 _20865_ (.A1(\datamem.data_ram[38][14] ),
    .A2(_07860_),
    .B1(_07851_),
    .B2(\datamem.data_ram[34][14] ),
    .C1(_08154_),
    .X(_08155_));
 sky130_fd_sc_hd__or2_1 _20866_ (.A(\datamem.data_ram[33][14] ),
    .B(_06934_),
    .X(_08156_));
 sky130_fd_sc_hd__o221a_1 _20867_ (.A1(\datamem.data_ram[39][14] ),
    .A2(_07859_),
    .B1(_07862_),
    .B2(\datamem.data_ram[37][14] ),
    .C1(_08156_),
    .X(_08157_));
 sky130_fd_sc_hd__o211a_1 _20868_ (.A1(\datamem.data_ram[35][14] ),
    .A2(_07851_),
    .B1(_07836_),
    .C1(_08157_),
    .X(_08158_));
 sky130_fd_sc_hd__a21o_1 _20869_ (.A1(_07833_),
    .A2(_08155_),
    .B1(_08158_),
    .X(_08159_));
 sky130_fd_sc_hd__o22a_1 _20870_ (.A1(\datamem.data_ram[53][14] ),
    .A2(_07037_),
    .B1(_06806_),
    .B2(\datamem.data_ram[52][14] ),
    .X(_08160_));
 sky130_fd_sc_hd__and2_1 _20871_ (.A(\datamem.data_ram[50][14] ),
    .B(_07832_),
    .X(_08161_));
 sky130_fd_sc_hd__a211o_1 _20872_ (.A1(\datamem.data_ram[51][14] ),
    .A2(_07849_),
    .B1(_08161_),
    .C1(_07851_),
    .X(_08162_));
 sky130_fd_sc_hd__o211a_1 _20873_ (.A1(\datamem.data_ram[54][14] ),
    .A2(_06683_),
    .B1(_08160_),
    .C1(_08162_),
    .X(_08163_));
 sky130_fd_sc_hd__o22a_1 _20874_ (.A1(\datamem.data_ram[48][14] ),
    .A2(_06647_),
    .B1(_06790_),
    .B2(\datamem.data_ram[49][14] ),
    .X(_08164_));
 sky130_fd_sc_hd__o211a_1 _20875_ (.A1(\datamem.data_ram[55][14] ),
    .A2(_07020_),
    .B1(_08164_),
    .C1(\rvcpu.dp.plem.ALUResultM[6] ),
    .X(_08165_));
 sky130_fd_sc_hd__a221o_1 _20876_ (.A1(_05347_),
    .A2(_08159_),
    .B1(_08163_),
    .B2(_08165_),
    .C1(_08124_),
    .X(_08166_));
 sky130_fd_sc_hd__mux2_1 _20877_ (.A0(\datamem.data_ram[42][14] ),
    .A1(\datamem.data_ram[43][14] ),
    .S(_07828_),
    .X(_08167_));
 sky130_fd_sc_hd__o22a_1 _20878_ (.A1(\datamem.data_ram[40][14] ),
    .A2(_06648_),
    .B1(_08167_),
    .B2(_07851_),
    .X(_08168_));
 sky130_fd_sc_hd__mux2_1 _20879_ (.A0(\datamem.data_ram[44][14] ),
    .A1(\datamem.data_ram[45][14] ),
    .S(_07827_),
    .X(_08169_));
 sky130_fd_sc_hd__mux2_1 _20880_ (.A0(\datamem.data_ram[46][14] ),
    .A1(\datamem.data_ram[47][14] ),
    .S(_07827_),
    .X(_08170_));
 sky130_fd_sc_hd__mux2_1 _20881_ (.A0(_08169_),
    .A1(_08170_),
    .S(_07821_),
    .X(_08171_));
 sky130_fd_sc_hd__o22a_1 _20882_ (.A1(\datamem.data_ram[41][14] ),
    .A2(_06658_),
    .B1(_08171_),
    .B2(_07845_),
    .X(_08172_));
 sky130_fd_sc_hd__o221a_1 _20883_ (.A1(\datamem.data_ram[56][14] ),
    .A2(_06837_),
    .B1(_06829_),
    .B2(\datamem.data_ram[59][14] ),
    .C1(_06714_),
    .X(_08173_));
 sky130_fd_sc_hd__mux2_1 _20884_ (.A0(\datamem.data_ram[60][14] ),
    .A1(\datamem.data_ram[61][14] ),
    .S(_07826_),
    .X(_08174_));
 sky130_fd_sc_hd__or2_1 _20885_ (.A(_07635_),
    .B(\datamem.data_ram[62][14] ),
    .X(_08175_));
 sky130_fd_sc_hd__o211a_1 _20886_ (.A1(\datamem.data_ram[63][14] ),
    .A2(_07831_),
    .B1(_08175_),
    .C1(_07821_),
    .X(_08176_));
 sky130_fd_sc_hd__a211o_1 _20887_ (.A1(_07839_),
    .A2(_08174_),
    .B1(_08176_),
    .C1(_07844_),
    .X(_08177_));
 sky130_fd_sc_hd__o221a_1 _20888_ (.A1(\datamem.data_ram[58][14] ),
    .A2(_06804_),
    .B1(_06790_),
    .B2(\datamem.data_ram[57][14] ),
    .C1(_08177_),
    .X(_08178_));
 sky130_fd_sc_hd__a21bo_1 _20889_ (.A1(_08173_),
    .A2(_08178_),
    .B1_N(_08124_),
    .X(_08179_));
 sky130_fd_sc_hd__a31o_1 _20890_ (.A1(_06753_),
    .A2(_08168_),
    .A3(_08172_),
    .B1(_08179_),
    .X(_08180_));
 sky130_fd_sc_hd__a21o_1 _20891_ (.A1(_08166_),
    .A2(_08180_),
    .B1(_06985_),
    .X(_08181_));
 sky130_fd_sc_hd__o211ai_4 _20892_ (.A1(_08125_),
    .A2(_08131_),
    .B1(_08153_),
    .C1(_08181_),
    .Y(_08182_));
 sky130_fd_sc_hd__o32a_1 _20893_ (.A1(_05391_),
    .A2(_06586_),
    .A3(_08123_),
    .B1(_08182_),
    .B2(_07120_),
    .X(_08183_));
 sky130_fd_sc_hd__mux2_1 _20894_ (.A0(\datamem.data_ram[2][22] ),
    .A1(\datamem.data_ram[3][22] ),
    .S(_07837_),
    .X(_08184_));
 sky130_fd_sc_hd__o221a_1 _20895_ (.A1(\datamem.data_ram[0][22] ),
    .A2(_06649_),
    .B1(_08184_),
    .B2(_07851_),
    .C1(_06681_),
    .X(_08185_));
 sky130_fd_sc_hd__mux2_1 _20896_ (.A0(\datamem.data_ram[4][22] ),
    .A1(\datamem.data_ram[5][22] ),
    .S(_07836_),
    .X(_08186_));
 sky130_fd_sc_hd__mux2_1 _20897_ (.A0(\datamem.data_ram[6][22] ),
    .A1(\datamem.data_ram[7][22] ),
    .S(_07836_),
    .X(_08187_));
 sky130_fd_sc_hd__mux2_1 _20898_ (.A0(_08186_),
    .A1(_08187_),
    .S(_07822_),
    .X(_08188_));
 sky130_fd_sc_hd__o22a_1 _20899_ (.A1(\datamem.data_ram[1][22] ),
    .A2(_06659_),
    .B1(_08188_),
    .B2(_07845_),
    .X(_08189_));
 sky130_fd_sc_hd__and2_1 _20900_ (.A(\datamem.data_ram[12][22] ),
    .B(_07833_),
    .X(_08190_));
 sky130_fd_sc_hd__a211o_1 _20901_ (.A1(\datamem.data_ram[13][22] ),
    .A2(_07837_),
    .B1(_08190_),
    .C1(_07863_),
    .X(_08191_));
 sky130_fd_sc_hd__o221a_1 _20902_ (.A1(_07823_),
    .A2(\datamem.data_ram[11][22] ),
    .B1(_07835_),
    .B2(\datamem.data_ram[10][22] ),
    .C1(_07845_),
    .X(_08192_));
 sky130_fd_sc_hd__o221a_1 _20903_ (.A1(_07635_),
    .A2(\datamem.data_ram[14][22] ),
    .B1(\datamem.data_ram[15][22] ),
    .B2(_07832_),
    .C1(_07867_),
    .X(_08193_));
 sky130_fd_sc_hd__or3_1 _20904_ (.A(_07840_),
    .B(_08192_),
    .C(_08193_),
    .X(_08194_));
 sky130_fd_sc_hd__o211a_1 _20905_ (.A1(\datamem.data_ram[9][22] ),
    .A2(_06701_),
    .B1(_08194_),
    .C1(_07081_),
    .X(_08195_));
 sky130_fd_sc_hd__o211a_1 _20906_ (.A1(\datamem.data_ram[8][22] ),
    .A2(_07191_),
    .B1(_08191_),
    .C1(_08195_),
    .X(_08196_));
 sky130_fd_sc_hd__a211o_1 _20907_ (.A1(_08185_),
    .A2(_08189_),
    .B1(_07071_),
    .C1(_08196_),
    .X(_08197_));
 sky130_fd_sc_hd__o221a_1 _20908_ (.A1(\datamem.data_ram[23][22] ),
    .A2(_07021_),
    .B1(_07182_),
    .B2(\datamem.data_ram[20][22] ),
    .C1(_06681_),
    .X(_08198_));
 sky130_fd_sc_hd__or2_1 _20909_ (.A(\datamem.data_ram[16][22] ),
    .B(_07829_),
    .X(_08199_));
 sky130_fd_sc_hd__o21a_1 _20910_ (.A1(\datamem.data_ram[17][22] ),
    .A2(_07833_),
    .B1(_07840_),
    .X(_08200_));
 sky130_fd_sc_hd__mux2_1 _20911_ (.A0(\datamem.data_ram[18][22] ),
    .A1(\datamem.data_ram[19][22] ),
    .S(_07836_),
    .X(_08201_));
 sky130_fd_sc_hd__a221o_1 _20912_ (.A1(_08199_),
    .A2(_08200_),
    .B1(_08201_),
    .B2(_07822_),
    .C1(_07868_),
    .X(_08202_));
 sky130_fd_sc_hd__o221a_1 _20913_ (.A1(\datamem.data_ram[22][22] ),
    .A2(_07028_),
    .B1(_07019_),
    .B2(\datamem.data_ram[21][22] ),
    .C1(_08202_),
    .X(_08203_));
 sky130_fd_sc_hd__mux2_1 _20914_ (.A0(\datamem.data_ram[30][22] ),
    .A1(\datamem.data_ram[31][22] ),
    .S(_07836_),
    .X(_08204_));
 sky130_fd_sc_hd__mux2_1 _20915_ (.A0(\datamem.data_ram[28][22] ),
    .A1(\datamem.data_ram[29][22] ),
    .S(_07827_),
    .X(_08205_));
 sky130_fd_sc_hd__or2_1 _20916_ (.A(_07863_),
    .B(_08205_),
    .X(_08206_));
 sky130_fd_sc_hd__o221a_1 _20917_ (.A1(\datamem.data_ram[26][22] ),
    .A2(_06692_),
    .B1(_06635_),
    .B2(\datamem.data_ram[27][22] ),
    .C1(_08206_),
    .X(_08207_));
 sky130_fd_sc_hd__o211a_1 _20918_ (.A1(_07860_),
    .A2(_08204_),
    .B1(_08207_),
    .C1(_07081_),
    .X(_08208_));
 sky130_fd_sc_hd__o221a_1 _20919_ (.A1(\datamem.data_ram[24][22] ),
    .A2(_07191_),
    .B1(_06659_),
    .B2(\datamem.data_ram[25][22] ),
    .C1(_08208_),
    .X(_08209_));
 sky130_fd_sc_hd__a211o_1 _20920_ (.A1(_08198_),
    .A2(_08203_),
    .B1(_08209_),
    .C1(_06916_),
    .X(_08210_));
 sky130_fd_sc_hd__mux2_1 _20921_ (.A0(\datamem.data_ram[46][22] ),
    .A1(\datamem.data_ram[47][22] ),
    .S(_07829_),
    .X(_08211_));
 sky130_fd_sc_hd__mux2_1 _20922_ (.A0(\datamem.data_ram[40][22] ),
    .A1(\datamem.data_ram[41][22] ),
    .S(_07827_),
    .X(_08212_));
 sky130_fd_sc_hd__mux2_1 _20923_ (.A0(\datamem.data_ram[42][22] ),
    .A1(\datamem.data_ram[43][22] ),
    .S(_07827_),
    .X(_08213_));
 sky130_fd_sc_hd__mux2_1 _20924_ (.A0(_08212_),
    .A1(_08213_),
    .S(_07821_),
    .X(_08214_));
 sky130_fd_sc_hd__mux2_1 _20925_ (.A0(\datamem.data_ram[44][22] ),
    .A1(\datamem.data_ram[45][22] ),
    .S(_07849_),
    .X(_08215_));
 sky130_fd_sc_hd__o22a_1 _20926_ (.A1(_07868_),
    .A2(_08214_),
    .B1(_08215_),
    .B2(_07863_),
    .X(_08216_));
 sky130_fd_sc_hd__o21a_1 _20927_ (.A1(_07860_),
    .A2(_08211_),
    .B1(_08216_),
    .X(_08217_));
 sky130_fd_sc_hd__mux2_1 _20928_ (.A0(\datamem.data_ram[38][22] ),
    .A1(\datamem.data_ram[39][22] ),
    .S(_07827_),
    .X(_08218_));
 sky130_fd_sc_hd__mux2_1 _20929_ (.A0(\datamem.data_ram[36][22] ),
    .A1(\datamem.data_ram[37][22] ),
    .S(_07827_),
    .X(_08219_));
 sky130_fd_sc_hd__mux2_1 _20930_ (.A0(_08218_),
    .A1(_08219_),
    .S(_07839_),
    .X(_08220_));
 sky130_fd_sc_hd__or2_1 _20931_ (.A(\datamem.data_ram[35][22] ),
    .B(_07831_),
    .X(_08221_));
 sky130_fd_sc_hd__o211a_1 _20932_ (.A1(\datamem.data_ram[34][22] ),
    .A2(_07849_),
    .B1(_08221_),
    .C1(_07636_),
    .X(_08222_));
 sky130_fd_sc_hd__a221o_1 _20933_ (.A1(\datamem.data_ram[32][22] ),
    .A2(_06973_),
    .B1(_08220_),
    .B2(_07868_),
    .C1(_08222_),
    .X(_08223_));
 sky130_fd_sc_hd__a211o_1 _20934_ (.A1(\datamem.data_ram[33][22] ),
    .A2(_07133_),
    .B1(_08223_),
    .C1(_06603_),
    .X(_08224_));
 sky130_fd_sc_hd__o21a_1 _20935_ (.A1(_06681_),
    .A2(_08217_),
    .B1(_08224_),
    .X(_08225_));
 sky130_fd_sc_hd__o221a_1 _20936_ (.A1(\datamem.data_ram[54][22] ),
    .A2(_06630_),
    .B1(_06665_),
    .B2(\datamem.data_ram[53][22] ),
    .C1(_06777_),
    .X(_08226_));
 sky130_fd_sc_hd__or2_1 _20937_ (.A(\datamem.data_ram[49][22] ),
    .B(_07832_),
    .X(_08227_));
 sky130_fd_sc_hd__o21a_1 _20938_ (.A1(\datamem.data_ram[48][22] ),
    .A2(_07828_),
    .B1(_07839_),
    .X(_08228_));
 sky130_fd_sc_hd__mux2_1 _20939_ (.A0(\datamem.data_ram[50][22] ),
    .A1(\datamem.data_ram[51][22] ),
    .S(_07835_),
    .X(_08229_));
 sky130_fd_sc_hd__a221o_1 _20940_ (.A1(_08227_),
    .A2(_08228_),
    .B1(_08229_),
    .B2(_07822_),
    .C1(_07868_),
    .X(_08230_));
 sky130_fd_sc_hd__o221a_1 _20941_ (.A1(\datamem.data_ram[55][22] ),
    .A2(_07021_),
    .B1(_06621_),
    .B2(\datamem.data_ram[52][22] ),
    .C1(_08230_),
    .X(_08231_));
 sky130_fd_sc_hd__o22a_1 _20942_ (.A1(\datamem.data_ram[59][22] ),
    .A2(_07851_),
    .B1(_06934_),
    .B2(\datamem.data_ram[57][22] ),
    .X(_08232_));
 sky130_fd_sc_hd__o221a_1 _20943_ (.A1(\datamem.data_ram[63][22] ),
    .A2(_07860_),
    .B1(_07863_),
    .B2(\datamem.data_ram[61][22] ),
    .C1(_08232_),
    .X(_08233_));
 sky130_fd_sc_hd__o22a_1 _20944_ (.A1(\datamem.data_ram[58][22] ),
    .A2(_06940_),
    .B1(_06934_),
    .B2(\datamem.data_ram[56][22] ),
    .X(_08234_));
 sky130_fd_sc_hd__o221a_1 _20945_ (.A1(\datamem.data_ram[62][22] ),
    .A2(_07860_),
    .B1(_07863_),
    .B2(\datamem.data_ram[60][22] ),
    .C1(_08234_),
    .X(_08235_));
 sky130_fd_sc_hd__or2_1 _20946_ (.A(_07829_),
    .B(_08235_),
    .X(_08236_));
 sky130_fd_sc_hd__o211a_1 _20947_ (.A1(_07823_),
    .A2(_08233_),
    .B1(_08236_),
    .C1(_07081_),
    .X(_08237_));
 sky130_fd_sc_hd__a211o_1 _20948_ (.A1(_08226_),
    .A2(_08231_),
    .B1(_08237_),
    .C1(_06753_),
    .X(_08238_));
 sky130_fd_sc_hd__o211a_1 _20949_ (.A1(_07071_),
    .A2(_08225_),
    .B1(_08238_),
    .C1(_06713_),
    .X(_08239_));
 sky130_fd_sc_hd__a31oi_4 _20950_ (.A1(_06985_),
    .A2(_08197_),
    .A3(_08210_),
    .B1(_08239_),
    .Y(_08240_));
 sky130_fd_sc_hd__o22a_1 _20951_ (.A1(_06590_),
    .A2(_08183_),
    .B1(_08240_),
    .B2(_07227_),
    .X(_08241_));
 sky130_fd_sc_hd__a21bo_1 _20952_ (.A1(_06988_),
    .A2(_08069_),
    .B1_N(_08241_),
    .X(_04443_));
 sky130_fd_sc_hd__o221a_1 _20953_ (.A1(\datamem.data_ram[54][15] ),
    .A2(_06625_),
    .B1(_06667_),
    .B2(\datamem.data_ram[55][15] ),
    .C1(_06676_),
    .X(_08242_));
 sky130_fd_sc_hd__or2_1 _20954_ (.A(\datamem.data_ram[49][15] ),
    .B(_06639_),
    .X(_08243_));
 sky130_fd_sc_hd__o21a_1 _20955_ (.A1(\datamem.data_ram[48][15] ),
    .A2(_06933_),
    .B1(_06606_),
    .X(_08244_));
 sky130_fd_sc_hd__mux2_1 _20956_ (.A0(\datamem.data_ram[50][15] ),
    .A1(\datamem.data_ram[51][15] ),
    .S(_06652_),
    .X(_08245_));
 sky130_fd_sc_hd__a221o_1 _20957_ (.A1(_08243_),
    .A2(_08244_),
    .B1(_08245_),
    .B2(_07819_),
    .C1(_06641_),
    .X(_08246_));
 sky130_fd_sc_hd__o221a_1 _20958_ (.A1(\datamem.data_ram[53][15] ),
    .A2(_06660_),
    .B1(_06616_),
    .B2(\datamem.data_ram[52][15] ),
    .C1(_08246_),
    .X(_08247_));
 sky130_fd_sc_hd__mux2_1 _20959_ (.A0(\datamem.data_ram[60][15] ),
    .A1(\datamem.data_ram[61][15] ),
    .S(_06933_),
    .X(_08248_));
 sky130_fd_sc_hd__o22a_1 _20960_ (.A1(\datamem.data_ram[58][15] ),
    .A2(_06608_),
    .B1(_06917_),
    .B2(_08248_),
    .X(_08249_));
 sky130_fd_sc_hd__mux2_1 _20961_ (.A0(\datamem.data_ram[62][15] ),
    .A1(\datamem.data_ram[63][15] ),
    .S(_06651_),
    .X(_08250_));
 sky130_fd_sc_hd__o22a_1 _20962_ (.A1(\datamem.data_ram[59][15] ),
    .A2(_06631_),
    .B1(_08250_),
    .B2(_06922_),
    .X(_08251_));
 sky130_fd_sc_hd__o211a_1 _20963_ (.A1(\datamem.data_ram[57][15] ),
    .A2(_06653_),
    .B1(_08251_),
    .C1(_06598_),
    .X(_08252_));
 sky130_fd_sc_hd__o211a_1 _20964_ (.A1(\datamem.data_ram[56][15] ),
    .A2(_06644_),
    .B1(_08249_),
    .C1(_08252_),
    .X(_08253_));
 sky130_fd_sc_hd__a21o_1 _20965_ (.A1(_08242_),
    .A2(_08247_),
    .B1(_08253_),
    .X(_08254_));
 sky130_fd_sc_hd__mux2_1 _20966_ (.A0(\datamem.data_ram[38][15] ),
    .A1(\datamem.data_ram[39][15] ),
    .S(_06651_),
    .X(_08255_));
 sky130_fd_sc_hd__mux2_1 _20967_ (.A0(\datamem.data_ram[36][15] ),
    .A1(\datamem.data_ram[37][15] ),
    .S(_06651_),
    .X(_08256_));
 sky130_fd_sc_hd__mux2_1 _20968_ (.A0(_08255_),
    .A1(_08256_),
    .S(_06606_),
    .X(_08257_));
 sky130_fd_sc_hd__or2_1 _20969_ (.A(\datamem.data_ram[35][15] ),
    .B(_06639_),
    .X(_08258_));
 sky130_fd_sc_hd__o211a_1 _20970_ (.A1(\datamem.data_ram[34][15] ),
    .A2(_07911_),
    .B1(_08258_),
    .C1(_06607_),
    .X(_08259_));
 sky130_fd_sc_hd__a221o_1 _20971_ (.A1(\datamem.data_ram[32][15] ),
    .A2(_06935_),
    .B1(_08257_),
    .B2(_06641_),
    .C1(_08259_),
    .X(_08260_));
 sky130_fd_sc_hd__a211o_1 _20972_ (.A1(\datamem.data_ram[33][15] ),
    .A2(_06945_),
    .B1(_08260_),
    .C1(_06598_),
    .X(_08261_));
 sky130_fd_sc_hd__mux2_1 _20973_ (.A0(\datamem.data_ram[40][15] ),
    .A1(\datamem.data_ram[41][15] ),
    .S(_06652_),
    .X(_08262_));
 sky130_fd_sc_hd__mux2_1 _20974_ (.A0(\datamem.data_ram[42][15] ),
    .A1(\datamem.data_ram[43][15] ),
    .S(_06652_),
    .X(_08263_));
 sky130_fd_sc_hd__mux2_1 _20975_ (.A0(_08262_),
    .A1(_08263_),
    .S(_07819_),
    .X(_08264_));
 sky130_fd_sc_hd__mux2_1 _20976_ (.A0(\datamem.data_ram[44][15] ),
    .A1(\datamem.data_ram[45][15] ),
    .S(_06933_),
    .X(_08265_));
 sky130_fd_sc_hd__a221o_1 _20977_ (.A1(net122),
    .A2(\datamem.data_ram[47][15] ),
    .B1(_06639_),
    .B2(\datamem.data_ram[46][15] ),
    .C1(_07838_),
    .X(_08266_));
 sky130_fd_sc_hd__o211a_1 _20978_ (.A1(_07819_),
    .A2(_08265_),
    .B1(_08266_),
    .C1(_06641_),
    .X(_08267_));
 sky130_fd_sc_hd__a211o_1 _20979_ (.A1(_07844_),
    .A2(_08264_),
    .B1(_08267_),
    .C1(_06676_),
    .X(_08268_));
 sky130_fd_sc_hd__a21o_1 _20980_ (.A1(_08261_),
    .A2(_08268_),
    .B1(_07903_),
    .X(_08269_));
 sky130_fd_sc_hd__mux2_1 _20981_ (.A0(\datamem.data_ram[12][15] ),
    .A1(\datamem.data_ram[13][15] ),
    .S(_06650_),
    .X(_08270_));
 sky130_fd_sc_hd__mux2_1 _20982_ (.A0(\datamem.data_ram[14][15] ),
    .A1(\datamem.data_ram[15][15] ),
    .S(_06650_),
    .X(_08271_));
 sky130_fd_sc_hd__mux2_1 _20983_ (.A0(_08270_),
    .A1(_08271_),
    .S(_06640_),
    .X(_08272_));
 sky130_fd_sc_hd__mux2_1 _20984_ (.A0(\datamem.data_ram[10][15] ),
    .A1(\datamem.data_ram[11][15] ),
    .S(_06651_),
    .X(_08273_));
 sky130_fd_sc_hd__or2_1 _20985_ (.A(_06928_),
    .B(_08273_),
    .X(_08274_));
 sky130_fd_sc_hd__o221a_1 _20986_ (.A1(\datamem.data_ram[8][15] ),
    .A2(_06643_),
    .B1(_08272_),
    .B2(_06614_),
    .C1(_08274_),
    .X(_08275_));
 sky130_fd_sc_hd__o211a_1 _20987_ (.A1(\datamem.data_ram[9][15] ),
    .A2(_06653_),
    .B1(_08275_),
    .C1(_06597_),
    .X(_08276_));
 sky130_fd_sc_hd__mux2_1 _20988_ (.A0(\datamem.data_ram[4][15] ),
    .A1(\datamem.data_ram[5][15] ),
    .S(_06652_),
    .X(_08277_));
 sky130_fd_sc_hd__mux2_1 _20989_ (.A0(\datamem.data_ram[0][15] ),
    .A1(\datamem.data_ram[1][15] ),
    .S(_06650_),
    .X(_08278_));
 sky130_fd_sc_hd__mux2_1 _20990_ (.A0(\datamem.data_ram[2][15] ),
    .A1(\datamem.data_ram[3][15] ),
    .S(_06650_),
    .X(_08279_));
 sky130_fd_sc_hd__mux2_1 _20991_ (.A0(_08278_),
    .A1(_08279_),
    .S(_06640_),
    .X(_08280_));
 sky130_fd_sc_hd__mux2_1 _20992_ (.A0(\datamem.data_ram[6][15] ),
    .A1(\datamem.data_ram[7][15] ),
    .S(_06651_),
    .X(_08281_));
 sky130_fd_sc_hd__o22a_1 _20993_ (.A1(_06641_),
    .A2(_08280_),
    .B1(_08281_),
    .B2(_06922_),
    .X(_08282_));
 sky130_fd_sc_hd__o211a_1 _20994_ (.A1(_06917_),
    .A2(_08277_),
    .B1(_08282_),
    .C1(_06675_),
    .X(_08283_));
 sky130_fd_sc_hd__or3_1 _20995_ (.A(_06594_),
    .B(_08276_),
    .C(_08283_),
    .X(_08284_));
 sky130_fd_sc_hd__mux2_1 _20996_ (.A0(\datamem.data_ram[30][15] ),
    .A1(\datamem.data_ram[31][15] ),
    .S(_06651_),
    .X(_08285_));
 sky130_fd_sc_hd__o22a_1 _20997_ (.A1(\datamem.data_ram[25][15] ),
    .A2(_06653_),
    .B1(_08285_),
    .B2(_06922_),
    .X(_08286_));
 sky130_fd_sc_hd__o221a_1 _20998_ (.A1(\datamem.data_ram[24][15] ),
    .A2(_06643_),
    .B1(_06616_),
    .B2(\datamem.data_ram[28][15] ),
    .C1(_08286_),
    .X(_08287_));
 sky130_fd_sc_hd__o22a_1 _20999_ (.A1(\datamem.data_ram[26][15] ),
    .A2(_06608_),
    .B1(_06631_),
    .B2(\datamem.data_ram[27][15] ),
    .X(_08288_));
 sky130_fd_sc_hd__o211a_1 _21000_ (.A1(\datamem.data_ram[29][15] ),
    .A2(_06660_),
    .B1(_08288_),
    .C1(_08124_),
    .X(_08289_));
 sky130_fd_sc_hd__o22a_1 _21001_ (.A1(\datamem.data_ram[21][15] ),
    .A2(_06660_),
    .B1(_06643_),
    .B2(\datamem.data_ram[16][15] ),
    .X(_08290_));
 sky130_fd_sc_hd__o221a_1 _21002_ (.A1(\datamem.data_ram[23][15] ),
    .A2(_06667_),
    .B1(_06616_),
    .B2(\datamem.data_ram[20][15] ),
    .C1(_08290_),
    .X(_08291_));
 sky130_fd_sc_hd__and2_1 _21003_ (.A(\datamem.data_ram[18][15] ),
    .B(_06639_),
    .X(_08292_));
 sky130_fd_sc_hd__a211o_1 _21004_ (.A1(\datamem.data_ram[19][15] ),
    .A2(_07911_),
    .B1(_08292_),
    .C1(_06928_),
    .X(_08293_));
 sky130_fd_sc_hd__o21ba_1 _21005_ (.A1(\datamem.data_ram[22][15] ),
    .A2(_06624_),
    .B1_N(\rvcpu.dp.plem.ALUResultM[5] ),
    .X(_08294_));
 sky130_fd_sc_hd__o211a_1 _21006_ (.A1(\datamem.data_ram[17][15] ),
    .A2(_06653_),
    .B1(_08293_),
    .C1(_08294_),
    .X(_08295_));
 sky130_fd_sc_hd__a22o_1 _21007_ (.A1(_08287_),
    .A2(_08289_),
    .B1(_08291_),
    .B2(_08295_),
    .X(_08296_));
 sky130_fd_sc_hd__a22o_1 _21008_ (.A1(_07176_),
    .A2(_08284_),
    .B1(_08296_),
    .B2(_06592_),
    .X(_08297_));
 sky130_fd_sc_hd__o211a_2 _21009_ (.A1(_07872_),
    .A2(_08254_),
    .B1(_08269_),
    .C1(_08297_),
    .X(_08298_));
 sky130_fd_sc_hd__inv_2 _21010_ (.A(_08298_),
    .Y(_08299_));
 sky130_fd_sc_hd__mux2_1 _21011_ (.A0(\datamem.data_ram[62][31] ),
    .A1(\datamem.data_ram[63][31] ),
    .S(_07912_),
    .X(_08300_));
 sky130_fd_sc_hd__or2_1 _21012_ (.A(_07859_),
    .B(_08300_),
    .X(_08301_));
 sky130_fd_sc_hd__o221a_1 _21013_ (.A1(\datamem.data_ram[56][31] ),
    .A2(_06811_),
    .B1(_06812_),
    .B2(\datamem.data_ram[59][31] ),
    .C1(_08301_),
    .X(_08302_));
 sky130_fd_sc_hd__mux2_1 _21014_ (.A0(\datamem.data_ram[60][31] ),
    .A1(\datamem.data_ram[61][31] ),
    .S(_07912_),
    .X(_08303_));
 sky130_fd_sc_hd__or2_1 _21015_ (.A(_07862_),
    .B(_08303_),
    .X(_08304_));
 sky130_fd_sc_hd__o221a_1 _21016_ (.A1(\datamem.data_ram[58][31] ),
    .A2(_06802_),
    .B1(_06780_),
    .B2(\datamem.data_ram[57][31] ),
    .C1(_08304_),
    .X(_08305_));
 sky130_fd_sc_hd__mux2_1 _21017_ (.A0(\datamem.data_ram[50][31] ),
    .A1(\datamem.data_ram[51][31] ),
    .S(_06652_),
    .X(_08306_));
 sky130_fd_sc_hd__o22a_1 _21018_ (.A1(\datamem.data_ram[48][31] ),
    .A2(_06643_),
    .B1(_08306_),
    .B2(_06940_),
    .X(_08307_));
 sky130_fd_sc_hd__o211a_1 _21019_ (.A1(\datamem.data_ram[55][31] ),
    .A2(_06667_),
    .B1(_08307_),
    .C1(_06676_),
    .X(_08308_));
 sky130_fd_sc_hd__o221a_1 _21020_ (.A1(\datamem.data_ram[53][31] ),
    .A2(_06721_),
    .B1(_06654_),
    .B2(\datamem.data_ram[49][31] ),
    .C1(_08308_),
    .X(_08309_));
 sky130_fd_sc_hd__o221a_1 _21021_ (.A1(\datamem.data_ram[54][31] ),
    .A2(_06626_),
    .B1(_06685_),
    .B2(\datamem.data_ram[52][31] ),
    .C1(_08309_),
    .X(_08310_));
 sky130_fd_sc_hd__a31o_1 _21022_ (.A1(_06851_),
    .A2(_08302_),
    .A3(_08305_),
    .B1(_08310_),
    .X(_08311_));
 sky130_fd_sc_hd__o22a_1 _21023_ (.A1(\datamem.data_ram[27][31] ),
    .A2(_06729_),
    .B1(_06654_),
    .B2(\datamem.data_ram[25][31] ),
    .X(_08312_));
 sky130_fd_sc_hd__mux2_1 _21024_ (.A0(\datamem.data_ram[30][31] ),
    .A1(\datamem.data_ram[31][31] ),
    .S(_07912_),
    .X(_08313_));
 sky130_fd_sc_hd__mux2_1 _21025_ (.A0(\datamem.data_ram[28][31] ),
    .A1(\datamem.data_ram[29][31] ),
    .S(_07911_),
    .X(_08314_));
 sky130_fd_sc_hd__or2_1 _21026_ (.A(_06917_),
    .B(_08314_),
    .X(_08315_));
 sky130_fd_sc_hd__o221a_1 _21027_ (.A1(\datamem.data_ram[24][31] ),
    .A2(_06644_),
    .B1(_08313_),
    .B2(_07859_),
    .C1(_08315_),
    .X(_08316_));
 sky130_fd_sc_hd__o211a_1 _21028_ (.A1(\datamem.data_ram[26][31] ),
    .A2(_06802_),
    .B1(_08312_),
    .C1(_08316_),
    .X(_08317_));
 sky130_fd_sc_hd__or2_1 _21029_ (.A(\datamem.data_ram[16][31] ),
    .B(_07912_),
    .X(_08318_));
 sky130_fd_sc_hd__o21a_1 _21030_ (.A1(\datamem.data_ram[17][31] ),
    .A2(_06944_),
    .B1(_07838_),
    .X(_08319_));
 sky130_fd_sc_hd__mux2_1 _21031_ (.A0(\datamem.data_ram[18][31] ),
    .A1(\datamem.data_ram[19][31] ),
    .S(_07824_),
    .X(_08320_));
 sky130_fd_sc_hd__a221o_1 _21032_ (.A1(_08318_),
    .A2(_08319_),
    .B1(_08320_),
    .B2(_07820_),
    .C1(_07866_),
    .X(_08321_));
 sky130_fd_sc_hd__o221a_1 _21033_ (.A1(\datamem.data_ram[21][31] ),
    .A2(_06721_),
    .B1(_06667_),
    .B2(\datamem.data_ram[23][31] ),
    .C1(_06676_),
    .X(_08322_));
 sky130_fd_sc_hd__o22a_1 _21034_ (.A1(\datamem.data_ram[22][31] ),
    .A2(_06625_),
    .B1(_06684_),
    .B2(\datamem.data_ram[20][31] ),
    .X(_08323_));
 sky130_fd_sc_hd__and3_1 _21035_ (.A(_08321_),
    .B(_08322_),
    .C(_08323_),
    .X(_08324_));
 sky130_fd_sc_hd__a211o_1 _21036_ (.A1(_06851_),
    .A2(_08317_),
    .B1(_08324_),
    .C1(_07176_),
    .X(_08325_));
 sky130_fd_sc_hd__mux2_1 _21037_ (.A0(\datamem.data_ram[12][31] ),
    .A1(\datamem.data_ram[13][31] ),
    .S(_07824_),
    .X(_08326_));
 sky130_fd_sc_hd__o221a_1 _21038_ (.A1(_06605_),
    .A2(\datamem.data_ram[11][31] ),
    .B1(_06933_),
    .B2(\datamem.data_ram[10][31] ),
    .C1(_07844_),
    .X(_08327_));
 sky130_fd_sc_hd__o221a_1 _21039_ (.A1(net122),
    .A2(\datamem.data_ram[14][31] ),
    .B1(\datamem.data_ram[15][31] ),
    .B2(_06639_),
    .C1(_06641_),
    .X(_08328_));
 sky130_fd_sc_hd__or3_1 _21040_ (.A(_07838_),
    .B(_08327_),
    .C(_08328_),
    .X(_08329_));
 sky130_fd_sc_hd__o221a_1 _21041_ (.A1(\datamem.data_ram[8][31] ),
    .A2(_06644_),
    .B1(_08326_),
    .B2(_06917_),
    .C1(_08329_),
    .X(_08330_));
 sky130_fd_sc_hd__o211a_1 _21042_ (.A1(\datamem.data_ram[9][31] ),
    .A2(_06655_),
    .B1(_08330_),
    .C1(_06599_),
    .X(_08331_));
 sky130_fd_sc_hd__mux2_1 _21043_ (.A0(\datamem.data_ram[6][31] ),
    .A1(\datamem.data_ram[7][31] ),
    .S(_07874_),
    .X(_08332_));
 sky130_fd_sc_hd__mux2_1 _21044_ (.A0(\datamem.data_ram[0][31] ),
    .A1(\datamem.data_ram[1][31] ),
    .S(_06933_),
    .X(_08333_));
 sky130_fd_sc_hd__mux2_1 _21045_ (.A0(\datamem.data_ram[2][31] ),
    .A1(\datamem.data_ram[3][31] ),
    .S(_06933_),
    .X(_08334_));
 sky130_fd_sc_hd__mux2_1 _21046_ (.A0(_08333_),
    .A1(_08334_),
    .S(_07819_),
    .X(_08335_));
 sky130_fd_sc_hd__mux2_1 _21047_ (.A0(\datamem.data_ram[4][31] ),
    .A1(\datamem.data_ram[5][31] ),
    .S(_07912_),
    .X(_08336_));
 sky130_fd_sc_hd__o22a_1 _21048_ (.A1(_07866_),
    .A2(_08335_),
    .B1(_08336_),
    .B2(_07862_),
    .X(_08337_));
 sky130_fd_sc_hd__o211a_1 _21049_ (.A1(_07859_),
    .A2(_08332_),
    .B1(_08337_),
    .C1(_06732_),
    .X(_08338_));
 sky130_fd_sc_hd__mux2_1 _21050_ (.A0(\datamem.data_ram[38][31] ),
    .A1(\datamem.data_ram[39][31] ),
    .S(_07826_),
    .X(_08339_));
 sky130_fd_sc_hd__mux2_1 _21051_ (.A0(\datamem.data_ram[32][31] ),
    .A1(\datamem.data_ram[33][31] ),
    .S(_07911_),
    .X(_08340_));
 sky130_fd_sc_hd__mux2_1 _21052_ (.A0(\datamem.data_ram[34][31] ),
    .A1(\datamem.data_ram[35][31] ),
    .S(_07911_),
    .X(_08341_));
 sky130_fd_sc_hd__mux2_1 _21053_ (.A0(_08340_),
    .A1(_08341_),
    .S(_07819_),
    .X(_08342_));
 sky130_fd_sc_hd__mux2_1 _21054_ (.A0(\datamem.data_ram[36][31] ),
    .A1(\datamem.data_ram[37][31] ),
    .S(_07825_),
    .X(_08343_));
 sky130_fd_sc_hd__o22a_1 _21055_ (.A1(_07866_),
    .A2(_08342_),
    .B1(_08343_),
    .B2(_07862_),
    .X(_08344_));
 sky130_fd_sc_hd__o211a_1 _21056_ (.A1(_07859_),
    .A2(_08339_),
    .B1(_08344_),
    .C1(_06732_),
    .X(_08345_));
 sky130_fd_sc_hd__mux2_1 _21057_ (.A0(\datamem.data_ram[44][31] ),
    .A1(\datamem.data_ram[45][31] ),
    .S(_07825_),
    .X(_08346_));
 sky130_fd_sc_hd__or2_1 _21058_ (.A(_07862_),
    .B(_08346_),
    .X(_08347_));
 sky130_fd_sc_hd__mux2_1 _21059_ (.A0(\datamem.data_ram[46][31] ),
    .A1(\datamem.data_ram[47][31] ),
    .S(_07825_),
    .X(_08348_));
 sky130_fd_sc_hd__mux4_1 _21060_ (.A0(\datamem.data_ram[40][31] ),
    .A1(\datamem.data_ram[41][31] ),
    .A2(\datamem.data_ram[42][31] ),
    .A3(\datamem.data_ram[43][31] ),
    .S0(_07824_),
    .S1(_07819_),
    .X(_08349_));
 sky130_fd_sc_hd__o22a_1 _21061_ (.A1(_07859_),
    .A2(_08348_),
    .B1(_08349_),
    .B2(_07866_),
    .X(_08350_));
 sky130_fd_sc_hd__a31o_1 _21062_ (.A1(_06599_),
    .A2(_08347_),
    .A3(_08350_),
    .B1(_07903_),
    .X(_08351_));
 sky130_fd_sc_hd__o32a_1 _21063_ (.A1(_07154_),
    .A2(_08331_),
    .A3(_08338_),
    .B1(_08345_),
    .B2(_08351_),
    .X(_08352_));
 sky130_fd_sc_hd__o211ai_4 _21064_ (.A1(_07872_),
    .A2(_08311_),
    .B1(_08325_),
    .C1(_08352_),
    .Y(_08353_));
 sky130_fd_sc_hd__mux2_1 _21065_ (.A0(_08299_),
    .A1(_08353_),
    .S(_06911_),
    .X(_08354_));
 sky130_fd_sc_hd__nor2_4 _21066_ (.A(_05347_),
    .B(_06860_),
    .Y(_08355_));
 sky130_fd_sc_hd__and2_1 _21067_ (.A(_06585_),
    .B(\datamem.data_ram[61][7] ),
    .X(_08356_));
 sky130_fd_sc_hd__a221o_1 _21068_ (.A1(\datamem.data_ram[60][7] ),
    .A2(_06944_),
    .B1(_08356_),
    .B2(_06666_),
    .C1(_06640_),
    .X(_08357_));
 sky130_fd_sc_hd__a221o_1 _21069_ (.A1(_06666_),
    .A2(\datamem.data_ram[63][7] ),
    .B1(_06944_),
    .B2(\datamem.data_ram[62][7] ),
    .C1(_07838_),
    .X(_08358_));
 sky130_fd_sc_hd__and3_1 _21070_ (.A(_07866_),
    .B(_08357_),
    .C(_08358_),
    .X(_08359_));
 sky130_fd_sc_hd__a221o_1 _21071_ (.A1(\datamem.data_ram[58][7] ),
    .A2(_06930_),
    .B1(_06946_),
    .B2(\datamem.data_ram[57][7] ),
    .C1(_08359_),
    .X(_08360_));
 sky130_fd_sc_hd__a221o_1 _21072_ (.A1(\datamem.data_ram[56][7] ),
    .A2(_06935_),
    .B1(_06941_),
    .B2(\datamem.data_ram[59][7] ),
    .C1(_08360_),
    .X(_08361_));
 sky130_fd_sc_hd__o221a_1 _21073_ (.A1(_07635_),
    .A2(\datamem.data_ram[46][7] ),
    .B1(\datamem.data_ram[47][7] ),
    .B2(_07831_),
    .C1(\rvcpu.dp.plem.ALUResultM[3] ),
    .X(_08362_));
 sky130_fd_sc_hd__or2_1 _21074_ (.A(\datamem.data_ram[44][7] ),
    .B(_07825_),
    .X(_08363_));
 sky130_fd_sc_hd__o211a_1 _21075_ (.A1(\datamem.data_ram[45][7] ),
    .A2(_07831_),
    .B1(_08363_),
    .C1(_05371_),
    .X(_08364_));
 sky130_fd_sc_hd__mux2_1 _21076_ (.A0(\datamem.data_ram[40][7] ),
    .A1(\datamem.data_ram[41][7] ),
    .S(_07825_),
    .X(_08365_));
 sky130_fd_sc_hd__o221a_1 _21077_ (.A1(_07823_),
    .A2(\datamem.data_ram[43][7] ),
    .B1(_07874_),
    .B2(\datamem.data_ram[42][7] ),
    .C1(\rvcpu.dp.plem.ALUResultM[3] ),
    .X(_08366_));
 sky130_fd_sc_hd__a211o_1 _21078_ (.A1(_05371_),
    .A2(_08365_),
    .B1(_08366_),
    .C1(\rvcpu.dp.plem.ALUResultM[4] ),
    .X(_08367_));
 sky130_fd_sc_hd__o311a_1 _21079_ (.A1(_06622_),
    .A2(_08362_),
    .A3(_08364_),
    .B1(_08367_),
    .C1(_07858_),
    .X(_08368_));
 sky130_fd_sc_hd__a211o_1 _21080_ (.A1(_08355_),
    .A2(_08361_),
    .B1(_08368_),
    .C1(_06733_),
    .X(_08369_));
 sky130_fd_sc_hd__o221a_1 _21081_ (.A1(_06605_),
    .A2(\datamem.data_ram[35][7] ),
    .B1(_07825_),
    .B2(\datamem.data_ram[34][7] ),
    .C1(_07844_),
    .X(_08370_));
 sky130_fd_sc_hd__o221a_1 _21082_ (.A1(_07823_),
    .A2(\datamem.data_ram[39][7] ),
    .B1(_07825_),
    .B2(\datamem.data_ram[38][7] ),
    .C1(_07866_),
    .X(_08371_));
 sky130_fd_sc_hd__o21a_1 _21083_ (.A1(_08370_),
    .A2(_08371_),
    .B1(_07820_),
    .X(_08372_));
 sky130_fd_sc_hd__mux2_1 _21084_ (.A0(\datamem.data_ram[36][7] ),
    .A1(\datamem.data_ram[37][7] ),
    .S(_07912_),
    .X(_08373_));
 sky130_fd_sc_hd__a22o_1 _21085_ (.A1(\datamem.data_ram[33][7] ),
    .A2(_06946_),
    .B1(_08373_),
    .B2(_06615_),
    .X(_08374_));
 sky130_fd_sc_hd__a211o_1 _21086_ (.A1(\datamem.data_ram[32][7] ),
    .A2(_06935_),
    .B1(_08372_),
    .C1(_08374_),
    .X(_08375_));
 sky130_fd_sc_hd__o221a_1 _21087_ (.A1(_06605_),
    .A2(\datamem.data_ram[51][7] ),
    .B1(_07911_),
    .B2(\datamem.data_ram[50][7] ),
    .C1(_07636_),
    .X(_08376_));
 sky130_fd_sc_hd__a221o_1 _21088_ (.A1(\datamem.data_ram[53][7] ),
    .A2(_06918_),
    .B1(_06923_),
    .B2(\datamem.data_ram[55][7] ),
    .C1(_08376_),
    .X(_08377_));
 sky130_fd_sc_hd__a221o_1 _21089_ (.A1(\datamem.data_ram[48][7] ),
    .A2(_06935_),
    .B1(_06953_),
    .B2(\datamem.data_ram[52][7] ),
    .C1(_08377_),
    .X(_08378_));
 sky130_fd_sc_hd__a221o_1 _21090_ (.A1(\datamem.data_ram[54][7] ),
    .A2(_06950_),
    .B1(_06946_),
    .B2(\datamem.data_ram[49][7] ),
    .C1(_08378_),
    .X(_08379_));
 sky130_fd_sc_hd__a221o_1 _21091_ (.A1(_07858_),
    .A2(_08375_),
    .B1(_08379_),
    .B2(_08355_),
    .C1(_06741_),
    .X(_08380_));
 sky130_fd_sc_hd__mux2_1 _21092_ (.A0(\datamem.data_ram[2][7] ),
    .A1(\datamem.data_ram[3][7] ),
    .S(_07912_),
    .X(_08381_));
 sky130_fd_sc_hd__a221o_1 _21093_ (.A1(\datamem.data_ram[0][7] ),
    .A2(_06935_),
    .B1(_08381_),
    .B2(_07636_),
    .C1(_06598_),
    .X(_08382_));
 sky130_fd_sc_hd__mux2_1 _21094_ (.A0(\datamem.data_ram[6][7] ),
    .A1(\datamem.data_ram[7][7] ),
    .S(_07824_),
    .X(_08383_));
 sky130_fd_sc_hd__mux2_1 _21095_ (.A0(\datamem.data_ram[4][7] ),
    .A1(\datamem.data_ram[5][7] ),
    .S(_07911_),
    .X(_08384_));
 sky130_fd_sc_hd__mux2_1 _21096_ (.A0(_08383_),
    .A1(_08384_),
    .S(_07838_),
    .X(_08385_));
 sky130_fd_sc_hd__a22o_1 _21097_ (.A1(\datamem.data_ram[1][7] ),
    .A2(_06946_),
    .B1(_08385_),
    .B2(_07867_),
    .X(_08386_));
 sky130_fd_sc_hd__mux2_1 _21098_ (.A0(\datamem.data_ram[12][7] ),
    .A1(\datamem.data_ram[13][7] ),
    .S(_07874_),
    .X(_08387_));
 sky130_fd_sc_hd__mux2_1 _21099_ (.A0(\datamem.data_ram[14][7] ),
    .A1(\datamem.data_ram[15][7] ),
    .S(_07824_),
    .X(_08388_));
 sky130_fd_sc_hd__or2_1 _21100_ (.A(\datamem.data_ram[8][7] ),
    .B(_06652_),
    .X(_08389_));
 sky130_fd_sc_hd__o211a_1 _21101_ (.A1(\datamem.data_ram[9][7] ),
    .A2(_06944_),
    .B1(_06642_),
    .C1(_08389_),
    .X(_08390_));
 sky130_fd_sc_hd__o221a_1 _21102_ (.A1(_06666_),
    .A2(\datamem.data_ram[10][7] ),
    .B1(\datamem.data_ram[11][7] ),
    .B2(_06944_),
    .C1(_07636_),
    .X(_08391_));
 sky130_fd_sc_hd__a211o_1 _21103_ (.A1(_06623_),
    .A2(_08388_),
    .B1(_08390_),
    .C1(_08391_),
    .X(_08392_));
 sky130_fd_sc_hd__a211o_1 _21104_ (.A1(_06615_),
    .A2(_08387_),
    .B1(_08392_),
    .C1(_06677_),
    .X(_08393_));
 sky130_fd_sc_hd__o211a_1 _21105_ (.A1(_08382_),
    .A2(_08386_),
    .B1(_06860_),
    .C1(_08393_),
    .X(_08394_));
 sky130_fd_sc_hd__mux2_1 _21106_ (.A0(\datamem.data_ram[18][7] ),
    .A1(\datamem.data_ram[19][7] ),
    .S(_06651_),
    .X(_08395_));
 sky130_fd_sc_hd__mux2_1 _21107_ (.A0(\datamem.data_ram[16][7] ),
    .A1(\datamem.data_ram[17][7] ),
    .S(_06651_),
    .X(_08396_));
 sky130_fd_sc_hd__or2_1 _21108_ (.A(_06640_),
    .B(_08396_),
    .X(_08397_));
 sky130_fd_sc_hd__o211a_1 _21109_ (.A1(_07838_),
    .A2(_08395_),
    .B1(_08397_),
    .C1(_07844_),
    .X(_08398_));
 sky130_fd_sc_hd__a221o_1 _21110_ (.A1(\datamem.data_ram[22][7] ),
    .A2(_06950_),
    .B1(_06919_),
    .B2(\datamem.data_ram[21][7] ),
    .C1(_08398_),
    .X(_08399_));
 sky130_fd_sc_hd__a221o_1 _21111_ (.A1(\datamem.data_ram[23][7] ),
    .A2(_06924_),
    .B1(_06953_),
    .B2(\datamem.data_ram[20][7] ),
    .C1(_08399_),
    .X(_08400_));
 sky130_fd_sc_hd__or2_1 _21112_ (.A(\datamem.data_ram[29][7] ),
    .B(_06639_),
    .X(_08401_));
 sky130_fd_sc_hd__o211a_1 _21113_ (.A1(\datamem.data_ram[28][7] ),
    .A2(_06652_),
    .B1(_08401_),
    .C1(_06615_),
    .X(_08402_));
 sky130_fd_sc_hd__a221o_1 _21114_ (.A1(\datamem.data_ram[30][7] ),
    .A2(_06950_),
    .B1(_06923_),
    .B2(\datamem.data_ram[31][7] ),
    .C1(_08402_),
    .X(_08403_));
 sky130_fd_sc_hd__a221o_1 _21115_ (.A1(\datamem.data_ram[26][7] ),
    .A2(_06929_),
    .B1(_06935_),
    .B2(\datamem.data_ram[24][7] ),
    .C1(_08403_),
    .X(_08404_));
 sky130_fd_sc_hd__a221o_2 _21116_ (.A1(\datamem.data_ram[27][7] ),
    .A2(_06941_),
    .B1(_06946_),
    .B2(\datamem.data_ram[25][7] ),
    .C1(_08404_),
    .X(_08405_));
 sky130_fd_sc_hd__a22o_1 _21117_ (.A1(_06732_),
    .A2(_08400_),
    .B1(_08405_),
    .B2(_08124_),
    .X(_08406_));
 sky130_fd_sc_hd__o22a_1 _21118_ (.A1(_06796_),
    .A2(_08394_),
    .B1(_08406_),
    .B2(_06751_),
    .X(_08407_));
 sky130_fd_sc_hd__a21oi_2 _21119_ (.A1(_08369_),
    .A2(_08380_),
    .B1(_08407_),
    .Y(_08408_));
 sky130_fd_sc_hd__mux2_1 _21120_ (.A0(\datamem.data_ram[44][23] ),
    .A1(\datamem.data_ram[45][23] ),
    .S(_07874_),
    .X(_08409_));
 sky130_fd_sc_hd__and2_1 _21121_ (.A(_06666_),
    .B(\datamem.data_ram[47][23] ),
    .X(_08410_));
 sky130_fd_sc_hd__a211o_1 _21122_ (.A1(\datamem.data_ram[46][23] ),
    .A2(_07831_),
    .B1(_08410_),
    .C1(_07838_),
    .X(_08411_));
 sky130_fd_sc_hd__o211a_1 _21123_ (.A1(_07820_),
    .A2(_08409_),
    .B1(_08411_),
    .C1(_07867_),
    .X(_08412_));
 sky130_fd_sc_hd__mux2_1 _21124_ (.A0(\datamem.data_ram[40][23] ),
    .A1(\datamem.data_ram[41][23] ),
    .S(_07874_),
    .X(_08413_));
 sky130_fd_sc_hd__a221o_1 _21125_ (.A1(_06666_),
    .A2(\datamem.data_ram[43][23] ),
    .B1(_06944_),
    .B2(\datamem.data_ram[42][23] ),
    .C1(_07838_),
    .X(_08414_));
 sky130_fd_sc_hd__o211a_1 _21126_ (.A1(_07820_),
    .A2(_08413_),
    .B1(_08414_),
    .C1(_07844_),
    .X(_08415_));
 sky130_fd_sc_hd__mux2_1 _21127_ (.A0(\datamem.data_ram[36][23] ),
    .A1(\datamem.data_ram[37][23] ),
    .S(_07826_),
    .X(_08416_));
 sky130_fd_sc_hd__mux2_1 _21128_ (.A0(\datamem.data_ram[38][23] ),
    .A1(\datamem.data_ram[39][23] ),
    .S(_07912_),
    .X(_08417_));
 sky130_fd_sc_hd__or2_1 _21129_ (.A(_07839_),
    .B(_08417_),
    .X(_08418_));
 sky130_fd_sc_hd__o211a_1 _21130_ (.A1(_07820_),
    .A2(_08416_),
    .B1(_08418_),
    .C1(_07867_),
    .X(_08419_));
 sky130_fd_sc_hd__mux4_1 _21131_ (.A0(\datamem.data_ram[32][23] ),
    .A1(\datamem.data_ram[33][23] ),
    .A2(\datamem.data_ram[34][23] ),
    .A3(\datamem.data_ram[35][23] ),
    .S0(_07874_),
    .S1(_07820_),
    .X(_08420_));
 sky130_fd_sc_hd__a21o_1 _21132_ (.A1(_07844_),
    .A2(_08420_),
    .B1(_06599_),
    .X(_08421_));
 sky130_fd_sc_hd__o32a_1 _21133_ (.A1(_06678_),
    .A2(_08412_),
    .A3(_08415_),
    .B1(_08419_),
    .B2(_08421_),
    .X(_08422_));
 sky130_fd_sc_hd__o221a_1 _21134_ (.A1(\datamem.data_ram[54][23] ),
    .A2(_06717_),
    .B1(_06725_),
    .B2(\datamem.data_ram[55][23] ),
    .C1(_06732_),
    .X(_08423_));
 sky130_fd_sc_hd__or2_1 _21135_ (.A(\datamem.data_ram[49][23] ),
    .B(_06944_),
    .X(_08424_));
 sky130_fd_sc_hd__o21a_1 _21136_ (.A1(\datamem.data_ram[48][23] ),
    .A2(_07874_),
    .B1(_07838_),
    .X(_08425_));
 sky130_fd_sc_hd__mux2_1 _21137_ (.A0(\datamem.data_ram[50][23] ),
    .A1(\datamem.data_ram[51][23] ),
    .S(_07825_),
    .X(_08426_));
 sky130_fd_sc_hd__a221o_1 _21138_ (.A1(_08424_),
    .A2(_08425_),
    .B1(_08426_),
    .B2(_07820_),
    .C1(_07866_),
    .X(_08427_));
 sky130_fd_sc_hd__o221a_1 _21139_ (.A1(\datamem.data_ram[53][23] ),
    .A2(_06722_),
    .B1(_06765_),
    .B2(\datamem.data_ram[52][23] ),
    .C1(_08427_),
    .X(_08428_));
 sky130_fd_sc_hd__or2_1 _21140_ (.A(\datamem.data_ram[56][23] ),
    .B(_06644_),
    .X(_08429_));
 sky130_fd_sc_hd__o221a_1 _21141_ (.A1(\datamem.data_ram[58][23] ),
    .A2(_06689_),
    .B1(_06729_),
    .B2(\datamem.data_ram[59][23] ),
    .C1(_08429_),
    .X(_08430_));
 sky130_fd_sc_hd__o22a_1 _21142_ (.A1(\datamem.data_ram[63][23] ),
    .A2(_07859_),
    .B1(_06917_),
    .B2(\datamem.data_ram[61][23] ),
    .X(_08431_));
 sky130_fd_sc_hd__o22a_1 _21143_ (.A1(\datamem.data_ram[62][23] ),
    .A2(_06922_),
    .B1(_06917_),
    .B2(\datamem.data_ram[60][23] ),
    .X(_08432_));
 sky130_fd_sc_hd__o221a_1 _21144_ (.A1(\datamem.data_ram[57][23] ),
    .A2(_06654_),
    .B1(_08432_),
    .B2(_07874_),
    .C1(_06598_),
    .X(_08433_));
 sky130_fd_sc_hd__o21a_1 _21145_ (.A1(_07831_),
    .A2(_08431_),
    .B1(_08433_),
    .X(_08434_));
 sky130_fd_sc_hd__a21o_1 _21146_ (.A1(_08430_),
    .A2(_08434_),
    .B1(_07872_),
    .X(_08435_));
 sky130_fd_sc_hd__a21o_1 _21147_ (.A1(_08423_),
    .A2(_08428_),
    .B1(_08435_),
    .X(_08436_));
 sky130_fd_sc_hd__or2_1 _21148_ (.A(\datamem.data_ram[20][23] ),
    .B(_06684_),
    .X(_08437_));
 sky130_fd_sc_hd__o22a_1 _21149_ (.A1(\datamem.data_ram[22][23] ),
    .A2(_06625_),
    .B1(_06645_),
    .B2(\datamem.data_ram[16][23] ),
    .X(_08438_));
 sky130_fd_sc_hd__o22a_1 _21150_ (.A1(\datamem.data_ram[23][23] ),
    .A2(_06667_),
    .B1(_06653_),
    .B2(\datamem.data_ram[17][23] ),
    .X(_08439_));
 sky130_fd_sc_hd__o221a_1 _21151_ (.A1(\datamem.data_ram[18][23] ),
    .A2(_06608_),
    .B1(_06631_),
    .B2(\datamem.data_ram[19][23] ),
    .C1(_06676_),
    .X(_08440_));
 sky130_fd_sc_hd__o211a_1 _21152_ (.A1(\datamem.data_ram[21][23] ),
    .A2(_06721_),
    .B1(_08439_),
    .C1(_08440_),
    .X(_08441_));
 sky130_fd_sc_hd__mux2_1 _21153_ (.A0(\datamem.data_ram[28][23] ),
    .A1(\datamem.data_ram[29][23] ),
    .S(_07825_),
    .X(_08442_));
 sky130_fd_sc_hd__mux2_1 _21154_ (.A0(\datamem.data_ram[30][23] ),
    .A1(\datamem.data_ram[31][23] ),
    .S(_07824_),
    .X(_08443_));
 sky130_fd_sc_hd__mux4_1 _21155_ (.A0(\datamem.data_ram[24][23] ),
    .A1(\datamem.data_ram[25][23] ),
    .A2(\datamem.data_ram[26][23] ),
    .A3(\datamem.data_ram[27][23] ),
    .S0(_06933_),
    .S1(_07819_),
    .X(_08444_));
 sky130_fd_sc_hd__o22a_1 _21156_ (.A1(_06922_),
    .A2(_08443_),
    .B1(_08444_),
    .B2(_07866_),
    .X(_08445_));
 sky130_fd_sc_hd__o211a_1 _21157_ (.A1(_07862_),
    .A2(_08442_),
    .B1(_08445_),
    .C1(_06598_),
    .X(_08446_));
 sky130_fd_sc_hd__a31o_1 _21158_ (.A1(_08437_),
    .A2(_08438_),
    .A3(_08441_),
    .B1(_08446_),
    .X(_08447_));
 sky130_fd_sc_hd__mux2_1 _21159_ (.A0(\datamem.data_ram[2][23] ),
    .A1(\datamem.data_ram[3][23] ),
    .S(_07912_),
    .X(_08448_));
 sky130_fd_sc_hd__o221a_1 _21160_ (.A1(\datamem.data_ram[0][23] ),
    .A2(_06645_),
    .B1(_08448_),
    .B2(_06940_),
    .C1(_06676_),
    .X(_08449_));
 sky130_fd_sc_hd__mux2_1 _21161_ (.A0(\datamem.data_ram[4][23] ),
    .A1(\datamem.data_ram[5][23] ),
    .S(_07911_),
    .X(_08450_));
 sky130_fd_sc_hd__mux2_1 _21162_ (.A0(\datamem.data_ram[6][23] ),
    .A1(\datamem.data_ram[7][23] ),
    .S(_07911_),
    .X(_08451_));
 sky130_fd_sc_hd__mux2_1 _21163_ (.A0(_08450_),
    .A1(_08451_),
    .S(_07819_),
    .X(_08452_));
 sky130_fd_sc_hd__o22a_1 _21164_ (.A1(\datamem.data_ram[1][23] ),
    .A2(_07242_),
    .B1(_08452_),
    .B2(_07844_),
    .X(_08453_));
 sky130_fd_sc_hd__mux2_1 _21165_ (.A0(\datamem.data_ram[8][23] ),
    .A1(\datamem.data_ram[9][23] ),
    .S(_06933_),
    .X(_08454_));
 sky130_fd_sc_hd__mux2_1 _21166_ (.A0(\datamem.data_ram[10][23] ),
    .A1(\datamem.data_ram[11][23] ),
    .S(_06933_),
    .X(_08455_));
 sky130_fd_sc_hd__mux2_1 _21167_ (.A0(_08454_),
    .A1(_08455_),
    .S(_07819_),
    .X(_08456_));
 sky130_fd_sc_hd__mux2_1 _21168_ (.A0(\datamem.data_ram[12][23] ),
    .A1(\datamem.data_ram[13][23] ),
    .S(_07824_),
    .X(_08457_));
 sky130_fd_sc_hd__or2_1 _21169_ (.A(_06917_),
    .B(_08457_),
    .X(_08458_));
 sky130_fd_sc_hd__mux2_1 _21170_ (.A0(\datamem.data_ram[14][23] ),
    .A1(\datamem.data_ram[15][23] ),
    .S(_07824_),
    .X(_08459_));
 sky130_fd_sc_hd__o21a_1 _21171_ (.A1(_07859_),
    .A2(_08459_),
    .B1(_06598_),
    .X(_08460_));
 sky130_fd_sc_hd__o211a_1 _21172_ (.A1(_07866_),
    .A2(_08456_),
    .B1(_08458_),
    .C1(_08460_),
    .X(_08461_));
 sky130_fd_sc_hd__a211o_1 _21173_ (.A1(_08449_),
    .A2(_08453_),
    .B1(_08461_),
    .C1(_06594_),
    .X(_08462_));
 sky130_fd_sc_hd__a22o_1 _21174_ (.A1(_06714_),
    .A2(_08447_),
    .B1(_08462_),
    .B2(_07177_),
    .X(_08463_));
 sky130_fd_sc_hd__o211ai_4 _21175_ (.A1(_07903_),
    .A2(_08422_),
    .B1(_08436_),
    .C1(_08463_),
    .Y(_08464_));
 sky130_fd_sc_hd__mux2_1 _21176_ (.A0(_08408_),
    .A1(_08464_),
    .S(_06911_),
    .X(_08465_));
 sky130_fd_sc_hd__mux2_1 _21177_ (.A0(_08354_),
    .A1(_08465_),
    .S(_06588_),
    .X(_08466_));
 sky130_fd_sc_hd__or2_1 _21178_ (.A(_06580_),
    .B(_08465_),
    .X(_08467_));
 sky130_fd_sc_hd__buf_2 _21179_ (.A(_06582_),
    .X(_08468_));
 sky130_fd_sc_hd__or2_1 _21180_ (.A(_08468_),
    .B(_08408_),
    .X(_08469_));
 sky130_fd_sc_hd__o211ai_2 _21181_ (.A1(_06583_),
    .A2(_08466_),
    .B1(_08467_),
    .C1(_08469_),
    .Y(_04444_));
 sky130_fd_sc_hd__o21a_1 _21182_ (.A1(\rvcpu.dp.plem.funct3M[0] ),
    .A2(\rvcpu.dp.plem.funct3M[2] ),
    .B1(\rvcpu.dp.plem.funct3M[1] ),
    .X(_00000_));
 sky130_fd_sc_hd__nor3_1 _21183_ (.A(\rvcpu.dp.plem.funct3M[0] ),
    .B(\rvcpu.dp.plem.funct3M[1] ),
    .C(\rvcpu.dp.plem.funct3M[2] ),
    .Y(_08470_));
 sky130_fd_sc_hd__o21ba_1 _21184_ (.A1(net118),
    .A2(_08470_),
    .B1_N(_08466_),
    .X(_08471_));
 sky130_fd_sc_hd__o22ai_1 _21185_ (.A1(_06910_),
    .A2(_06580_),
    .B1(_08468_),
    .B2(_06909_),
    .Y(_08472_));
 sky130_fd_sc_hd__or2_1 _21186_ (.A(_08471_),
    .B(_08472_),
    .X(_08473_));
 sky130_fd_sc_hd__clkbuf_1 _21187_ (.A(_08473_),
    .X(_04445_));
 sky130_fd_sc_hd__o22ai_1 _21188_ (.A1(_07277_),
    .A2(_07119_),
    .B1(_07070_),
    .B2(_06915_),
    .Y(_08474_));
 sky130_fd_sc_hd__or2_1 _21189_ (.A(_08471_),
    .B(_08474_),
    .X(_08475_));
 sky130_fd_sc_hd__clkbuf_1 _21190_ (.A(_08475_),
    .X(_04446_));
 sky130_fd_sc_hd__o22a_1 _21191_ (.A1(_06915_),
    .A2(_07368_),
    .B1(_07413_),
    .B2(_07277_),
    .X(_08476_));
 sky130_fd_sc_hd__or2b_1 _21192_ (.A(_08471_),
    .B_N(_08476_),
    .X(_08477_));
 sky130_fd_sc_hd__clkbuf_1 _21193_ (.A(_08477_),
    .X(_04416_));
 sky130_fd_sc_hd__o22ai_1 _21194_ (.A1(_07277_),
    .A2(net37),
    .B1(_07461_),
    .B2(_06915_),
    .Y(_08478_));
 sky130_fd_sc_hd__or2_1 _21195_ (.A(_08471_),
    .B(_08478_),
    .X(_08479_));
 sky130_fd_sc_hd__clkbuf_1 _21196_ (.A(_08479_),
    .X(_04417_));
 sky130_fd_sc_hd__o22ai_1 _21197_ (.A1(_07277_),
    .A2(_07737_),
    .B1(_07691_),
    .B2(_06915_),
    .Y(_08480_));
 sky130_fd_sc_hd__or2_1 _21198_ (.A(_08471_),
    .B(_08480_),
    .X(_08481_));
 sky130_fd_sc_hd__clkbuf_1 _21199_ (.A(_08481_),
    .X(_04418_));
 sky130_fd_sc_hd__o22a_1 _21200_ (.A1(_08468_),
    .A2(_07920_),
    .B1(_07965_),
    .B2(_06580_),
    .X(_08482_));
 sky130_fd_sc_hd__or2b_1 _21201_ (.A(_08471_),
    .B_N(_08482_),
    .X(_08483_));
 sky130_fd_sc_hd__clkbuf_1 _21202_ (.A(_08483_),
    .X(_04419_));
 sky130_fd_sc_hd__o22ai_1 _21203_ (.A1(_06915_),
    .A2(_08123_),
    .B1(_08182_),
    .B2(_07277_),
    .Y(_08484_));
 sky130_fd_sc_hd__or2_1 _21204_ (.A(_08471_),
    .B(_08484_),
    .X(_08485_));
 sky130_fd_sc_hd__clkbuf_1 _21205_ (.A(_08485_),
    .X(_04420_));
 sky130_fd_sc_hd__nor2_1 _21206_ (.A(_06580_),
    .B(_08354_),
    .Y(_08486_));
 sky130_fd_sc_hd__a211o_1 _21207_ (.A1(_06987_),
    .A2(_08298_),
    .B1(_08471_),
    .C1(_08486_),
    .X(_04421_));
 sky130_fd_sc_hd__buf_2 _21208_ (.A(_08468_),
    .X(_08487_));
 sky130_fd_sc_hd__or2_4 _21209_ (.A(\rvcpu.dp.plem.funct3M[2] ),
    .B(_06580_),
    .X(_08488_));
 sky130_fd_sc_hd__o21ba_1 _21210_ (.A1(_08354_),
    .A2(_08488_),
    .B1_N(_08471_),
    .X(_08489_));
 sky130_fd_sc_hd__clkbuf_2 _21211_ (.A(_08489_),
    .X(_08490_));
 sky130_fd_sc_hd__o21ai_1 _21212_ (.A1(_08487_),
    .A2(_06799_),
    .B1(_08490_),
    .Y(_04422_));
 sky130_fd_sc_hd__o21ai_1 _21213_ (.A1(_08487_),
    .A2(_07226_),
    .B1(_08490_),
    .Y(_04423_));
 sky130_fd_sc_hd__o21ai_1 _21214_ (.A1(_08487_),
    .A2(_07276_),
    .B1(_08490_),
    .Y(_04424_));
 sky130_fd_sc_hd__o21ai_1 _21215_ (.A1(_08487_),
    .A2(_07597_),
    .B1(_08490_),
    .Y(_04425_));
 sky130_fd_sc_hd__o21ai_1 _21216_ (.A1(_08487_),
    .A2(_07781_),
    .B1(_08490_),
    .Y(_04427_));
 sky130_fd_sc_hd__o21ai_1 _21217_ (.A1(_08487_),
    .A2(_07857_),
    .B1(_08490_),
    .Y(_04428_));
 sky130_fd_sc_hd__o21ai_1 _21218_ (.A1(_08487_),
    .A2(_08240_),
    .B1(_08490_),
    .Y(_04429_));
 sky130_fd_sc_hd__o21ai_1 _21219_ (.A1(_08487_),
    .A2(_08464_),
    .B1(_08490_),
    .Y(_04430_));
 sky130_fd_sc_hd__o21ai_1 _21220_ (.A1(_06862_),
    .A2(_08487_),
    .B1(_08490_),
    .Y(_04431_));
 sky130_fd_sc_hd__o21ai_1 _21221_ (.A1(_08487_),
    .A2(_07070_),
    .B1(_08490_),
    .Y(_04432_));
 sky130_fd_sc_hd__o21ai_1 _21222_ (.A1(_08468_),
    .A2(_07368_),
    .B1(_08489_),
    .Y(_04433_));
 sky130_fd_sc_hd__o21ai_1 _21223_ (.A1(_08468_),
    .A2(_07461_),
    .B1(_08489_),
    .Y(_04434_));
 sky130_fd_sc_hd__o21ai_1 _21224_ (.A1(_08468_),
    .A2(_07691_),
    .B1(_08489_),
    .Y(_04435_));
 sky130_fd_sc_hd__o21ai_1 _21225_ (.A1(_08468_),
    .A2(net36),
    .B1(_08489_),
    .Y(_04436_));
 sky130_fd_sc_hd__o21ai_1 _21226_ (.A1(_08468_),
    .A2(_08123_),
    .B1(_08489_),
    .Y(_04438_));
 sky130_fd_sc_hd__o21ai_1 _21227_ (.A1(_08468_),
    .A2(_08353_),
    .B1(_08489_),
    .Y(_04439_));
 sky130_fd_sc_hd__or4_1 _21228_ (.A(\datamem.data_ram[53][14] ),
    .B(\datamem.data_ram[52][14] ),
    .C(\datamem.data_ram[52][7] ),
    .D(\datamem.data_ram[53][7] ),
    .X(_08491_));
 sky130_fd_sc_hd__or4_2 _21229_ (.A(\datamem.data_ram[52][6] ),
    .B(\datamem.data_ram[53][6] ),
    .C(\datamem.data_ram[52][30] ),
    .D(\datamem.data_ram[52][22] ),
    .X(_08492_));
 sky130_fd_sc_hd__or4_1 _21230_ (.A(\datamem.data_ram[52][29] ),
    .B(\datamem.data_ram[52][21] ),
    .C(\datamem.data_ram[53][13] ),
    .D(\datamem.data_ram[52][13] ),
    .X(_08493_));
 sky130_fd_sc_hd__or4_1 _21231_ (.A(\datamem.data_ram[52][31] ),
    .B(\datamem.data_ram[52][23] ),
    .C(\datamem.data_ram[53][15] ),
    .D(\datamem.data_ram[52][15] ),
    .X(_08494_));
 sky130_fd_sc_hd__or3_1 _21232_ (.A(_08492_),
    .B(_08493_),
    .C(_08494_),
    .X(_08495_));
 sky130_fd_sc_hd__or4b_1 _21233_ (.A(\datamem.data_ram[52][27] ),
    .B(\datamem.data_ram[52][19] ),
    .C(\datamem.data_ram[53][11] ),
    .D_N(\datamem.data_ram[52][11] ),
    .X(_08496_));
 sky130_fd_sc_hd__nand2_1 _21234_ (.A(\datamem.data_ram[52][10] ),
    .B(\datamem.data_ram[52][3] ),
    .Y(_08497_));
 sky130_fd_sc_hd__or4_1 _21235_ (.A(\datamem.data_ram[53][10] ),
    .B(\datamem.data_ram[53][3] ),
    .C(_08496_),
    .D(_08497_),
    .X(_08498_));
 sky130_fd_sc_hd__nand2_2 _21236_ (.A(\datamem.data_ram[52][12] ),
    .B(\datamem.data_ram[53][12] ),
    .Y(_08499_));
 sky130_fd_sc_hd__and4_1 _21237_ (.A(\datamem.data_ram[52][4] ),
    .B(\datamem.data_ram[53][4] ),
    .C(\datamem.data_ram[52][28] ),
    .D(\datamem.data_ram[52][20] ),
    .X(_08500_));
 sky130_fd_sc_hd__or4b_2 _21238_ (.A(\datamem.data_ram[52][5] ),
    .B(\datamem.data_ram[53][5] ),
    .C(_08499_),
    .D_N(_08500_),
    .X(_08501_));
 sky130_fd_sc_hd__or4b_1 _21239_ (.A(\datamem.data_ram[53][8] ),
    .B(\datamem.data_ram[52][8] ),
    .C(\datamem.data_ram[52][1] ),
    .D_N(\datamem.data_ram[53][1] ),
    .X(_08502_));
 sky130_fd_sc_hd__nand2_1 _21240_ (.A(\datamem.data_ram[52][24] ),
    .B(\datamem.data_ram[52][16] ),
    .Y(_08503_));
 sky130_fd_sc_hd__or4_2 _21241_ (.A(\datamem.data_ram[52][0] ),
    .B(\datamem.data_ram[53][0] ),
    .C(_08502_),
    .D(_08503_),
    .X(_08504_));
 sky130_fd_sc_hd__nand2_1 _21242_ (.A(\datamem.data_ram[52][17] ),
    .B(\datamem.data_ram[52][9] ),
    .Y(_08505_));
 sky130_fd_sc_hd__and4b_1 _21243_ (.A_N(\datamem.data_ram[53][2] ),
    .B(\datamem.data_ram[52][26] ),
    .C(\datamem.data_ram[52][18] ),
    .D(\datamem.data_ram[52][2] ),
    .X(_08506_));
 sky130_fd_sc_hd__or4b_1 _21244_ (.A(\datamem.data_ram[52][25] ),
    .B(_08505_),
    .C(\datamem.data_ram[53][9] ),
    .D_N(_08506_),
    .X(_08507_));
 sky130_fd_sc_hd__or4_1 _21245_ (.A(_08498_),
    .B(_08501_),
    .C(_08504_),
    .D(_08507_),
    .X(_08508_));
 sky130_fd_sc_hd__nor3_1 _21246_ (.A(_08491_),
    .B(_08495_),
    .C(_08508_),
    .Y(net34));
 sky130_fd_sc_hd__inv_2 _21247_ (.A(\rvcpu.dp.plfd.InstrD[19] ),
    .Y(_08509_));
 sky130_fd_sc_hd__buf_2 _21248_ (.A(_08509_),
    .X(_08510_));
 sky130_fd_sc_hd__buf_2 _21249_ (.A(_08510_),
    .X(_08511_));
 sky130_fd_sc_hd__clkbuf_4 _21250_ (.A(\rvcpu.dp.plfd.InstrD[18] ),
    .X(_08512_));
 sky130_fd_sc_hd__clkbuf_4 _21251_ (.A(_08512_),
    .X(_08513_));
 sky130_fd_sc_hd__clkbuf_4 _21252_ (.A(\rvcpu.dp.plfd.InstrD[17] ),
    .X(_08514_));
 sky130_fd_sc_hd__buf_2 _21253_ (.A(_08514_),
    .X(_08515_));
 sky130_fd_sc_hd__buf_6 _21254_ (.A(\rvcpu.dp.plfd.InstrD[15] ),
    .X(_08516_));
 sky130_fd_sc_hd__clkbuf_8 _21255_ (.A(_08516_),
    .X(_08517_));
 sky130_fd_sc_hd__buf_4 _21256_ (.A(\rvcpu.dp.plfd.InstrD[16] ),
    .X(_08518_));
 sky130_fd_sc_hd__buf_4 _21257_ (.A(_08518_),
    .X(_08519_));
 sky130_fd_sc_hd__mux4_1 _21258_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][0] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][0] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][0] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][0] ),
    .S0(_08517_),
    .S1(_08519_),
    .X(_08520_));
 sky130_fd_sc_hd__nor2_1 _21259_ (.A(_08515_),
    .B(_08520_),
    .Y(_08521_));
 sky130_fd_sc_hd__inv_2 _21260_ (.A(\rvcpu.dp.plfd.InstrD[17] ),
    .Y(_08522_));
 sky130_fd_sc_hd__clkbuf_4 _21261_ (.A(_08522_),
    .X(_08523_));
 sky130_fd_sc_hd__clkbuf_8 _21262_ (.A(\rvcpu.dp.plfd.InstrD[15] ),
    .X(_08524_));
 sky130_fd_sc_hd__clkbuf_8 _21263_ (.A(_08524_),
    .X(_08525_));
 sky130_fd_sc_hd__buf_4 _21264_ (.A(\rvcpu.dp.plfd.InstrD[16] ),
    .X(_08526_));
 sky130_fd_sc_hd__clkbuf_8 _21265_ (.A(_08526_),
    .X(_08527_));
 sky130_fd_sc_hd__clkbuf_8 _21266_ (.A(_08527_),
    .X(_08528_));
 sky130_fd_sc_hd__mux4_1 _21267_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][0] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][0] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][0] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][0] ),
    .S0(_08525_),
    .S1(_08528_),
    .X(_08529_));
 sky130_fd_sc_hd__nor2_1 _21268_ (.A(_08523_),
    .B(_08529_),
    .Y(_08530_));
 sky130_fd_sc_hd__clkbuf_4 _21269_ (.A(_08522_),
    .X(_08531_));
 sky130_fd_sc_hd__clkbuf_4 _21270_ (.A(_08531_),
    .X(_08532_));
 sky130_fd_sc_hd__clkbuf_8 _21271_ (.A(\rvcpu.dp.plfd.InstrD[16] ),
    .X(_08533_));
 sky130_fd_sc_hd__buf_6 _21272_ (.A(_08533_),
    .X(_08534_));
 sky130_fd_sc_hd__buf_4 _21273_ (.A(\rvcpu.dp.plfd.InstrD[15] ),
    .X(_08535_));
 sky130_fd_sc_hd__clkbuf_8 _21274_ (.A(_08535_),
    .X(_08536_));
 sky130_fd_sc_hd__clkbuf_8 _21275_ (.A(_08536_),
    .X(_08537_));
 sky130_fd_sc_hd__mux4_1 _21276_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][0] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][0] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][0] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][0] ),
    .S0(_08534_),
    .S1(_08537_),
    .X(_08538_));
 sky130_fd_sc_hd__nor2_1 _21277_ (.A(_08532_),
    .B(_08538_),
    .Y(_08539_));
 sky130_fd_sc_hd__buf_4 _21278_ (.A(\rvcpu.dp.plfd.InstrD[17] ),
    .X(_08540_));
 sky130_fd_sc_hd__clkbuf_4 _21279_ (.A(_08540_),
    .X(_08541_));
 sky130_fd_sc_hd__buf_4 _21280_ (.A(_08541_),
    .X(_08542_));
 sky130_fd_sc_hd__mux4_1 _21281_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][0] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][0] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][0] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][0] ),
    .S0(_08525_),
    .S1(_08528_),
    .X(_08543_));
 sky130_fd_sc_hd__o21ai_1 _21282_ (.A1(_08542_),
    .A2(_08543_),
    .B1(_08513_),
    .Y(_08544_));
 sky130_fd_sc_hd__o32a_1 _21283_ (.A1(_08513_),
    .A2(_08521_),
    .A3(_08530_),
    .B1(_08539_),
    .B2(_08544_),
    .X(_08545_));
 sky130_fd_sc_hd__nor2_1 _21284_ (.A(_08511_),
    .B(_08545_),
    .Y(_08546_));
 sky130_fd_sc_hd__clkbuf_4 _21285_ (.A(_08532_),
    .X(_08547_));
 sky130_fd_sc_hd__clkbuf_8 _21286_ (.A(\rvcpu.dp.plfd.InstrD[15] ),
    .X(_08548_));
 sky130_fd_sc_hd__buf_6 _21287_ (.A(_08548_),
    .X(_08549_));
 sky130_fd_sc_hd__buf_4 _21288_ (.A(_08549_),
    .X(_08550_));
 sky130_fd_sc_hd__clkbuf_8 _21289_ (.A(_08550_),
    .X(_08551_));
 sky130_fd_sc_hd__buf_4 _21290_ (.A(\rvcpu.dp.plfd.InstrD[16] ),
    .X(_08552_));
 sky130_fd_sc_hd__buf_4 _21291_ (.A(_08552_),
    .X(_08553_));
 sky130_fd_sc_hd__clkbuf_4 _21292_ (.A(_08553_),
    .X(_08554_));
 sky130_fd_sc_hd__buf_4 _21293_ (.A(_08554_),
    .X(_08555_));
 sky130_fd_sc_hd__mux4_1 _21294_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][0] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][0] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][0] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][0] ),
    .S0(_08551_),
    .S1(_08555_),
    .X(_08556_));
 sky130_fd_sc_hd__inv_2 _21295_ (.A(\rvcpu.dp.plfd.InstrD[18] ),
    .Y(_08557_));
 sky130_fd_sc_hd__nor2_4 _21296_ (.A(\rvcpu.dp.plfd.InstrD[19] ),
    .B(_08557_),
    .Y(_08558_));
 sky130_fd_sc_hd__clkbuf_8 _21297_ (.A(\rvcpu.dp.plfd.InstrD[16] ),
    .X(_08559_));
 sky130_fd_sc_hd__buf_4 _21298_ (.A(_08559_),
    .X(_08560_));
 sky130_fd_sc_hd__clkbuf_4 _21299_ (.A(_08536_),
    .X(_08561_));
 sky130_fd_sc_hd__mux4_1 _21300_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][0] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][0] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][0] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][0] ),
    .S0(_08560_),
    .S1(_08561_),
    .X(_08562_));
 sky130_fd_sc_hd__or2_1 _21301_ (.A(_08542_),
    .B(_08562_),
    .X(_08563_));
 sky130_fd_sc_hd__o211a_1 _21302_ (.A1(_08547_),
    .A2(_08556_),
    .B1(_08558_),
    .C1(_08563_),
    .X(_08564_));
 sky130_fd_sc_hd__clkbuf_4 _21303_ (.A(_08532_),
    .X(_08565_));
 sky130_fd_sc_hd__clkbuf_8 _21304_ (.A(_08549_),
    .X(_08566_));
 sky130_fd_sc_hd__buf_8 _21305_ (.A(_08566_),
    .X(_08567_));
 sky130_fd_sc_hd__clkbuf_8 _21306_ (.A(_08552_),
    .X(_08568_));
 sky130_fd_sc_hd__buf_4 _21307_ (.A(_08568_),
    .X(_08569_));
 sky130_fd_sc_hd__buf_6 _21308_ (.A(_08569_),
    .X(_08570_));
 sky130_fd_sc_hd__mux4_1 _21309_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][0] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][0] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][0] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][0] ),
    .S0(_08567_),
    .S1(_08570_),
    .X(_08571_));
 sky130_fd_sc_hd__clkbuf_8 _21310_ (.A(_08541_),
    .X(_08572_));
 sky130_fd_sc_hd__mux4_1 _21311_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][0] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][0] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][0] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][0] ),
    .S0(_08566_),
    .S1(_08569_),
    .X(_08573_));
 sky130_fd_sc_hd__or2_1 _21312_ (.A(_08572_),
    .B(_08573_),
    .X(_08574_));
 sky130_fd_sc_hd__nor2_4 _21313_ (.A(\rvcpu.dp.plfd.InstrD[19] ),
    .B(_08512_),
    .Y(_08575_));
 sky130_fd_sc_hd__clkbuf_4 _21314_ (.A(_08575_),
    .X(_08576_));
 sky130_fd_sc_hd__o211a_1 _21315_ (.A1(_08565_),
    .A2(_08571_),
    .B1(_08574_),
    .C1(_08576_),
    .X(_08577_));
 sky130_fd_sc_hd__clkbuf_8 _21316_ (.A(_08517_),
    .X(_08578_));
 sky130_fd_sc_hd__or2_2 _21317_ (.A(\rvcpu.dp.plfd.InstrD[19] ),
    .B(\rvcpu.dp.plfd.InstrD[18] ),
    .X(_08579_));
 sky130_fd_sc_hd__inv_2 _21318_ (.A(\rvcpu.dp.plfd.InstrD[15] ),
    .Y(_08580_));
 sky130_fd_sc_hd__inv_2 _21319_ (.A(\rvcpu.dp.plfd.InstrD[16] ),
    .Y(_08581_));
 sky130_fd_sc_hd__inv_2 _21320_ (.A(\rvcpu.dp.plde.RdE[3] ),
    .Y(_08582_));
 sky130_fd_sc_hd__a22o_1 _21321_ (.A1(\rvcpu.dp.plfd.InstrD[18] ),
    .A2(_08582_),
    .B1(\rvcpu.dp.plde.RdE[4] ),
    .B2(_08509_),
    .X(_08583_));
 sky130_fd_sc_hd__a221o_1 _21322_ (.A1(_08580_),
    .A2(\rvcpu.dp.plde.RdE[0] ),
    .B1(\rvcpu.dp.plde.RdE[1] ),
    .B2(_08581_),
    .C1(_08583_),
    .X(_08584_));
 sky130_fd_sc_hd__xnor2_1 _21323_ (.A(\rvcpu.dp.plfd.InstrD[17] ),
    .B(\rvcpu.dp.plde.RdE[2] ),
    .Y(_08585_));
 sky130_fd_sc_hd__o22a_1 _21324_ (.A1(_08580_),
    .A2(\rvcpu.dp.plde.RdE[0] ),
    .B1(_08582_),
    .B2(\rvcpu.dp.plfd.InstrD[18] ),
    .X(_08586_));
 sky130_fd_sc_hd__o221a_1 _21325_ (.A1(_08581_),
    .A2(\rvcpu.dp.plde.RdE[1] ),
    .B1(\rvcpu.dp.plde.RdE[4] ),
    .B2(_08509_),
    .C1(_08586_),
    .X(_08587_));
 sky130_fd_sc_hd__and3b_2 _21326_ (.A_N(_08584_),
    .B(_08585_),
    .C(_08587_),
    .X(_08588_));
 sky130_fd_sc_hd__inv_2 _21327_ (.A(\rvcpu.dp.plfd.InstrD[24] ),
    .Y(_08589_));
 sky130_fd_sc_hd__xor2_1 _21328_ (.A(\rvcpu.dp.plfd.InstrD[22] ),
    .B(\rvcpu.dp.plde.RdE[2] ),
    .X(_08590_));
 sky130_fd_sc_hd__a221o_1 _21329_ (.A1(\rvcpu.dp.plfd.InstrD[23] ),
    .A2(_08582_),
    .B1(\rvcpu.dp.plde.RdE[4] ),
    .B2(_08589_),
    .C1(_08590_),
    .X(_08591_));
 sky130_fd_sc_hd__clkbuf_8 _21330_ (.A(\rvcpu.dp.plfd.InstrD[20] ),
    .X(_08592_));
 sky130_fd_sc_hd__xnor2_1 _21331_ (.A(_08592_),
    .B(\rvcpu.dp.plde.RdE[0] ),
    .Y(_08593_));
 sky130_fd_sc_hd__o221a_1 _21332_ (.A1(\rvcpu.dp.plfd.InstrD[23] ),
    .A2(_08582_),
    .B1(\rvcpu.dp.plde.RdE[4] ),
    .B2(_08589_),
    .C1(_08593_),
    .X(_08594_));
 sky130_fd_sc_hd__buf_4 _21333_ (.A(\rvcpu.dp.plfd.InstrD[21] ),
    .X(_08595_));
 sky130_fd_sc_hd__xnor2_1 _21334_ (.A(_08595_),
    .B(\rvcpu.dp.plde.RdE[1] ),
    .Y(_08596_));
 sky130_fd_sc_hd__and3b_2 _21335_ (.A_N(_08591_),
    .B(_08594_),
    .C(_08596_),
    .X(_08597_));
 sky130_fd_sc_hd__o21ai_4 _21336_ (.A1(_08588_),
    .A2(_08597_),
    .B1(\rvcpu.dp.hu.ResultSrcE0 ),
    .Y(_08598_));
 sky130_fd_sc_hd__or4_1 _21337_ (.A(\rvcpu.ALUResultE[23] ),
    .B(_06294_),
    .C(_06305_),
    .D(\rvcpu.ALUResultE[29] ),
    .X(_08599_));
 sky130_fd_sc_hd__or4_1 _21338_ (.A(\rvcpu.ALUResultE[1] ),
    .B(\rvcpu.ALUResultE[2] ),
    .C(\rvcpu.ALUResultE[3] ),
    .D(\rvcpu.ALUResultE[4] ),
    .X(_08600_));
 sky130_fd_sc_hd__or4_1 _21339_ (.A(\rvcpu.ALUResultE[5] ),
    .B(\rvcpu.ALUResultE[6] ),
    .C(\rvcpu.ALUResultE[7] ),
    .D(_08600_),
    .X(_08601_));
 sky130_fd_sc_hd__or3_1 _21340_ (.A(\rvcpu.ALUResultE[8] ),
    .B(\rvcpu.ALUResultE[9] ),
    .C(_08601_),
    .X(_08602_));
 sky130_fd_sc_hd__or4_1 _21341_ (.A(\rvcpu.ALUResultE[10] ),
    .B(\rvcpu.ALUResultE[12] ),
    .C(\rvcpu.ALUResultE[16] ),
    .D(_08602_),
    .X(_08603_));
 sky130_fd_sc_hd__or2_1 _21342_ (.A(\rvcpu.ALUResultE[11] ),
    .B(\rvcpu.ALUResultE[13] ),
    .X(_08604_));
 sky130_fd_sc_hd__or4_1 _21343_ (.A(\rvcpu.ALUResultE[14] ),
    .B(\rvcpu.ALUResultE[17] ),
    .C(_08603_),
    .D(_08604_),
    .X(_08605_));
 sky130_fd_sc_hd__a211o_1 _21344_ (.A1(_05239_),
    .A2(_06195_),
    .B1(_06209_),
    .C1(\rvcpu.ALUResultE[18] ),
    .X(_08606_));
 sky130_fd_sc_hd__or4_1 _21345_ (.A(_06122_),
    .B(_06130_),
    .C(\rvcpu.ALUResultE[24] ),
    .D(_08606_),
    .X(_08607_));
 sky130_fd_sc_hd__or4_1 _21346_ (.A(\rvcpu.ALUResultE[19] ),
    .B(\rvcpu.ALUResultE[21] ),
    .C(_08605_),
    .D(_08607_),
    .X(_08608_));
 sky130_fd_sc_hd__or4_1 _21347_ (.A(\rvcpu.ALUResultE[22] ),
    .B(\rvcpu.ALUResultE[25] ),
    .C(\rvcpu.ALUResultE[26] ),
    .D(\rvcpu.ALUResultE[28] ),
    .X(_08609_));
 sky130_fd_sc_hd__or4_1 _21348_ (.A(_05747_),
    .B(_05794_),
    .C(_08608_),
    .D(_08609_),
    .X(_08610_));
 sky130_fd_sc_hd__or4_1 _21349_ (.A(\rvcpu.ALUResultE[31] ),
    .B(\rvcpu.ALUResultE[30] ),
    .C(_08599_),
    .D(_08610_),
    .X(_08611_));
 sky130_fd_sc_hd__or4bb_1 _21350_ (.A(\rvcpu.dp.plde.funct3E[2] ),
    .B(\rvcpu.dp.plde.funct3E[1] ),
    .C_N(_08611_),
    .D_N(\rvcpu.dp.plde.funct3E[0] ),
    .X(_08612_));
 sky130_fd_sc_hd__or3_1 _21351_ (.A(\rvcpu.dp.plde.funct3E[2] ),
    .B(\rvcpu.dp.plde.funct3E[0] ),
    .C(\rvcpu.dp.plde.funct3E[1] ),
    .X(_08613_));
 sky130_fd_sc_hd__or4bb_1 _21352_ (.A(\rvcpu.dp.plde.funct3E[0] ),
    .B(\rvcpu.dp.plde.funct3E[1] ),
    .C_N(\rvcpu.ALUResultE[31] ),
    .D_N(\rvcpu.dp.plde.funct3E[2] ),
    .X(_08614_));
 sky130_fd_sc_hd__nand2_1 _21353_ (.A(\rvcpu.dp.plde.funct3E[0] ),
    .B(\rvcpu.dp.Cout ),
    .Y(_08615_));
 sky130_fd_sc_hd__o211a_1 _21354_ (.A1(\rvcpu.dp.plde.funct3E[0] ),
    .A2(\rvcpu.dp.Cout ),
    .B1(\rvcpu.dp.plde.funct3E[1] ),
    .C1(\rvcpu.dp.plde.funct3E[2] ),
    .X(_08616_));
 sky130_fd_sc_hd__nand3b_1 _21355_ (.A_N(\rvcpu.dp.plde.funct3E[1] ),
    .B(\rvcpu.dp.plde.funct3E[0] ),
    .C(\rvcpu.dp.plde.funct3E[2] ),
    .Y(_08617_));
 sky130_fd_sc_hd__o2bb2a_1 _21356_ (.A1_N(_08615_),
    .A2_N(_08616_),
    .B1(\rvcpu.ALUResultE[31] ),
    .B2(_08617_),
    .X(_08618_));
 sky130_fd_sc_hd__o211a_1 _21357_ (.A1(_08611_),
    .A2(_08613_),
    .B1(_08614_),
    .C1(_08618_),
    .X(_08619_));
 sky130_fd_sc_hd__a21bo_2 _21358_ (.A1(_08612_),
    .A2(_08619_),
    .B1_N(\rvcpu.dp.plde.BranchE ),
    .X(_08620_));
 sky130_fd_sc_hd__nor2_2 _21359_ (.A(\rvcpu.dp.plde.JumpE ),
    .B(\rvcpu.dp.plde.JalrE ),
    .Y(_08621_));
 sky130_fd_sc_hd__and3_4 _21360_ (.A(_08598_),
    .B(_08620_),
    .C(_08621_),
    .X(_08622_));
 sky130_fd_sc_hd__o41a_1 _21361_ (.A1(_08514_),
    .A2(_08569_),
    .A3(_08578_),
    .A4(_08579_),
    .B1(_08622_),
    .X(_08623_));
 sky130_fd_sc_hd__buf_2 _21362_ (.A(_08623_),
    .X(_08624_));
 sky130_fd_sc_hd__buf_2 _21363_ (.A(_08624_),
    .X(_08625_));
 sky130_fd_sc_hd__o31a_1 _21364_ (.A1(_08546_),
    .A2(_08564_),
    .A3(_08577_),
    .B1(_08625_),
    .X(_01028_));
 sky130_fd_sc_hd__buf_2 _21365_ (.A(_08557_),
    .X(_08626_));
 sky130_fd_sc_hd__buf_2 _21366_ (.A(_08626_),
    .X(_08627_));
 sky130_fd_sc_hd__clkbuf_8 _21367_ (.A(_08535_),
    .X(_08628_));
 sky130_fd_sc_hd__buf_4 _21368_ (.A(_08552_),
    .X(_08629_));
 sky130_fd_sc_hd__mux4_1 _21369_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][1] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][1] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][1] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][1] ),
    .S0(_08628_),
    .S1(_08629_),
    .X(_08630_));
 sky130_fd_sc_hd__buf_4 _21370_ (.A(_08535_),
    .X(_08631_));
 sky130_fd_sc_hd__buf_4 _21371_ (.A(_08559_),
    .X(_08632_));
 sky130_fd_sc_hd__mux4_1 _21372_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][1] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][1] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][1] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][1] ),
    .S0(_08631_),
    .S1(_08632_),
    .X(_08633_));
 sky130_fd_sc_hd__mux2_1 _21373_ (.A0(_08630_),
    .A1(_08633_),
    .S(_08541_),
    .X(_08634_));
 sky130_fd_sc_hd__buf_4 _21374_ (.A(_08559_),
    .X(_08635_));
 sky130_fd_sc_hd__buf_4 _21375_ (.A(_08535_),
    .X(_08636_));
 sky130_fd_sc_hd__buf_4 _21376_ (.A(_08636_),
    .X(_08637_));
 sky130_fd_sc_hd__mux4_1 _21377_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][1] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][1] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][1] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][1] ),
    .S0(_08635_),
    .S1(_08637_),
    .X(_08638_));
 sky130_fd_sc_hd__nor2_1 _21378_ (.A(_08532_),
    .B(_08638_),
    .Y(_08639_));
 sky130_fd_sc_hd__mux4_1 _21379_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][1] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][1] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][1] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][1] ),
    .S0(_08517_),
    .S1(_08519_),
    .X(_08640_));
 sky130_fd_sc_hd__o21ai_1 _21380_ (.A1(_08515_),
    .A2(_08640_),
    .B1(_08513_),
    .Y(_08641_));
 sky130_fd_sc_hd__o2bb2a_1 _21381_ (.A1_N(_08627_),
    .A2_N(_08634_),
    .B1(_08639_),
    .B2(_08641_),
    .X(_08642_));
 sky130_fd_sc_hd__nor2_1 _21382_ (.A(_08511_),
    .B(_08642_),
    .Y(_08643_));
 sky130_fd_sc_hd__mux4_1 _21383_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][1] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][1] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][1] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][1] ),
    .S0(_08551_),
    .S1(_08555_),
    .X(_08644_));
 sky130_fd_sc_hd__mux4_1 _21384_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][1] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][1] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][1] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][1] ),
    .S0(_08550_),
    .S1(_08554_),
    .X(_08645_));
 sky130_fd_sc_hd__or2_1 _21385_ (.A(_08542_),
    .B(_08645_),
    .X(_08646_));
 sky130_fd_sc_hd__o211a_1 _21386_ (.A1(_08547_),
    .A2(_08644_),
    .B1(_08646_),
    .C1(_08575_),
    .X(_08647_));
 sky130_fd_sc_hd__mux4_1 _21387_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][1] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][1] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][1] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][1] ),
    .S0(_08567_),
    .S1(_08570_),
    .X(_08648_));
 sky130_fd_sc_hd__buf_6 _21388_ (.A(_08533_),
    .X(_08649_));
 sky130_fd_sc_hd__mux4_1 _21389_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][1] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][1] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][1] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][1] ),
    .S0(_08649_),
    .S1(_08537_),
    .X(_08650_));
 sky130_fd_sc_hd__or2_1 _21390_ (.A(_08572_),
    .B(_08650_),
    .X(_08651_));
 sky130_fd_sc_hd__buf_2 _21391_ (.A(_08558_),
    .X(_08652_));
 sky130_fd_sc_hd__o211a_1 _21392_ (.A1(_08565_),
    .A2(_08648_),
    .B1(_08651_),
    .C1(_08652_),
    .X(_08653_));
 sky130_fd_sc_hd__o31a_1 _21393_ (.A1(_08643_),
    .A2(_08647_),
    .A3(_08653_),
    .B1(_08625_),
    .X(_01029_));
 sky130_fd_sc_hd__mux4_1 _21394_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][2] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][2] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][2] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][2] ),
    .S0(_08628_),
    .S1(_08629_),
    .X(_08654_));
 sky130_fd_sc_hd__mux4_1 _21395_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][2] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][2] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][2] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][2] ),
    .S0(_08631_),
    .S1(_08632_),
    .X(_08655_));
 sky130_fd_sc_hd__mux2_1 _21396_ (.A0(_08654_),
    .A1(_08655_),
    .S(_08541_),
    .X(_08656_));
 sky130_fd_sc_hd__mux4_1 _21397_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][2] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][2] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][2] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][2] ),
    .S0(_08635_),
    .S1(_08637_),
    .X(_08657_));
 sky130_fd_sc_hd__nor2_1 _21398_ (.A(_08532_),
    .B(_08657_),
    .Y(_08658_));
 sky130_fd_sc_hd__mux4_1 _21399_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][2] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][2] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][2] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][2] ),
    .S0(_08517_),
    .S1(_08519_),
    .X(_08659_));
 sky130_fd_sc_hd__o21ai_1 _21400_ (.A1(_08515_),
    .A2(_08659_),
    .B1(_08513_),
    .Y(_08660_));
 sky130_fd_sc_hd__o2bb2a_1 _21401_ (.A1_N(_08627_),
    .A2_N(_08656_),
    .B1(_08658_),
    .B2(_08660_),
    .X(_08661_));
 sky130_fd_sc_hd__nor2_1 _21402_ (.A(_08511_),
    .B(_08661_),
    .Y(_08662_));
 sky130_fd_sc_hd__clkbuf_4 _21403_ (.A(_08532_),
    .X(_08663_));
 sky130_fd_sc_hd__mux4_1 _21404_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][2] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][2] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][2] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][2] ),
    .S0(_08551_),
    .S1(_08555_),
    .X(_08664_));
 sky130_fd_sc_hd__mux4_1 _21405_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][2] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][2] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][2] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][2] ),
    .S0(_08560_),
    .S1(_08561_),
    .X(_08665_));
 sky130_fd_sc_hd__or2_1 _21406_ (.A(_08542_),
    .B(_08665_),
    .X(_08666_));
 sky130_fd_sc_hd__o211a_1 _21407_ (.A1(_08663_),
    .A2(_08664_),
    .B1(_08666_),
    .C1(_08652_),
    .X(_08667_));
 sky130_fd_sc_hd__mux4_1 _21408_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][2] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][2] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][2] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][2] ),
    .S0(_08567_),
    .S1(_08570_),
    .X(_08668_));
 sky130_fd_sc_hd__mux4_1 _21409_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][2] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][2] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][2] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][2] ),
    .S0(_08566_),
    .S1(_08569_),
    .X(_08669_));
 sky130_fd_sc_hd__or2_1 _21410_ (.A(_08572_),
    .B(_08669_),
    .X(_08670_));
 sky130_fd_sc_hd__o211a_1 _21411_ (.A1(_08565_),
    .A2(_08668_),
    .B1(_08670_),
    .C1(_08576_),
    .X(_08671_));
 sky130_fd_sc_hd__o31a_1 _21412_ (.A1(_08662_),
    .A2(_08667_),
    .A3(_08671_),
    .B1(_08625_),
    .X(_01030_));
 sky130_fd_sc_hd__buf_2 _21413_ (.A(_08623_),
    .X(_08672_));
 sky130_fd_sc_hd__buf_4 _21414_ (.A(\rvcpu.dp.plfd.InstrD[17] ),
    .X(_08673_));
 sky130_fd_sc_hd__mux4_2 _21415_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][3] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][3] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][3] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][3] ),
    .S0(_08549_),
    .S1(_08527_),
    .X(_08674_));
 sky130_fd_sc_hd__or2_1 _21416_ (.A(_08673_),
    .B(_08674_),
    .X(_08675_));
 sky130_fd_sc_hd__mux4_1 _21417_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][3] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][3] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][3] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][3] ),
    .S0(_08533_),
    .S1(_08636_),
    .X(_08676_));
 sky130_fd_sc_hd__o21a_1 _21418_ (.A1(_08531_),
    .A2(_08676_),
    .B1(_08512_),
    .X(_08677_));
 sky130_fd_sc_hd__mux4_1 _21419_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][3] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][3] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][3] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][3] ),
    .S0(_08524_),
    .S1(_08527_),
    .X(_08678_));
 sky130_fd_sc_hd__mux4_1 _21420_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][3] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][3] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][3] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][3] ),
    .S0(_08524_),
    .S1(_08527_),
    .X(_08679_));
 sky130_fd_sc_hd__mux2_1 _21421_ (.A0(_08678_),
    .A1(_08679_),
    .S(_08514_),
    .X(_08680_));
 sky130_fd_sc_hd__a221o_1 _21422_ (.A1(_08675_),
    .A2(_08677_),
    .B1(_08680_),
    .B2(_08626_),
    .C1(_08510_),
    .X(_08681_));
 sky130_fd_sc_hd__clkbuf_4 _21423_ (.A(_08523_),
    .X(_08682_));
 sky130_fd_sc_hd__buf_4 _21424_ (.A(_08628_),
    .X(_08683_));
 sky130_fd_sc_hd__buf_4 _21425_ (.A(_08560_),
    .X(_08684_));
 sky130_fd_sc_hd__mux4_1 _21426_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][3] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][3] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][3] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][3] ),
    .S0(_08683_),
    .S1(_08684_),
    .X(_08685_));
 sky130_fd_sc_hd__buf_4 _21427_ (.A(_08540_),
    .X(_08686_));
 sky130_fd_sc_hd__buf_6 _21428_ (.A(_08535_),
    .X(_08687_));
 sky130_fd_sc_hd__mux4_1 _21429_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][3] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][3] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][3] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][3] ),
    .S0(_08687_),
    .S1(_08649_),
    .X(_08688_));
 sky130_fd_sc_hd__clkbuf_4 _21430_ (.A(_08579_),
    .X(_08689_));
 sky130_fd_sc_hd__a21o_1 _21431_ (.A1(_08686_),
    .A2(_08688_),
    .B1(_08689_),
    .X(_08690_));
 sky130_fd_sc_hd__a21o_1 _21432_ (.A1(_08682_),
    .A2(_08685_),
    .B1(_08690_),
    .X(_08691_));
 sky130_fd_sc_hd__clkbuf_4 _21433_ (.A(_08523_),
    .X(_08692_));
 sky130_fd_sc_hd__clkbuf_8 _21434_ (.A(_08533_),
    .X(_08693_));
 sky130_fd_sc_hd__mux4_1 _21435_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][3] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][3] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][3] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][3] ),
    .S0(_08693_),
    .S1(_08578_),
    .X(_08694_));
 sky130_fd_sc_hd__buf_2 _21436_ (.A(_08540_),
    .X(_08695_));
 sky130_fd_sc_hd__clkbuf_8 _21437_ (.A(_08535_),
    .X(_08696_));
 sky130_fd_sc_hd__mux4_1 _21438_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][3] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][3] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][3] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][3] ),
    .S0(_08696_),
    .S1(_08568_),
    .X(_08697_));
 sky130_fd_sc_hd__and2_1 _21439_ (.A(_08695_),
    .B(_08697_),
    .X(_08698_));
 sky130_fd_sc_hd__nand2_2 _21440_ (.A(_08509_),
    .B(_08512_),
    .Y(_08699_));
 sky130_fd_sc_hd__clkbuf_4 _21441_ (.A(_08699_),
    .X(_08700_));
 sky130_fd_sc_hd__a211o_1 _21442_ (.A1(_08692_),
    .A2(_08694_),
    .B1(_08698_),
    .C1(_08700_),
    .X(_08701_));
 sky130_fd_sc_hd__and4_1 _21443_ (.A(_08672_),
    .B(_08681_),
    .C(_08691_),
    .D(_08701_),
    .X(_08702_));
 sky130_fd_sc_hd__clkbuf_1 _21444_ (.A(_08702_),
    .X(_01031_));
 sky130_fd_sc_hd__buf_4 _21445_ (.A(_08535_),
    .X(_08703_));
 sky130_fd_sc_hd__mux4_1 _21446_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][4] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][4] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][4] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][4] ),
    .S0(_08703_),
    .S1(_08629_),
    .X(_08704_));
 sky130_fd_sc_hd__mux4_1 _21447_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][4] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][4] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][4] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][4] ),
    .S0(_08631_),
    .S1(_08632_),
    .X(_08705_));
 sky130_fd_sc_hd__mux2_1 _21448_ (.A0(_08704_),
    .A1(_08705_),
    .S(_08541_),
    .X(_08706_));
 sky130_fd_sc_hd__mux4_1 _21449_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][4] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][4] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][4] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][4] ),
    .S0(_08635_),
    .S1(_08637_),
    .X(_08707_));
 sky130_fd_sc_hd__nor2_1 _21450_ (.A(_08532_),
    .B(_08707_),
    .Y(_08708_));
 sky130_fd_sc_hd__mux4_1 _21451_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][4] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][4] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][4] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][4] ),
    .S0(_08517_),
    .S1(_08519_),
    .X(_08709_));
 sky130_fd_sc_hd__o21ai_1 _21452_ (.A1(_08515_),
    .A2(_08709_),
    .B1(_08513_),
    .Y(_08710_));
 sky130_fd_sc_hd__o2bb2a_1 _21453_ (.A1_N(_08627_),
    .A2_N(_08706_),
    .B1(_08708_),
    .B2(_08710_),
    .X(_08711_));
 sky130_fd_sc_hd__nor2_1 _21454_ (.A(_08511_),
    .B(_08711_),
    .Y(_08712_));
 sky130_fd_sc_hd__mux4_1 _21455_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][4] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][4] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][4] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][4] ),
    .S0(_08551_),
    .S1(_08555_),
    .X(_08713_));
 sky130_fd_sc_hd__mux4_1 _21456_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][4] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][4] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][4] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][4] ),
    .S0(_08550_),
    .S1(_08554_),
    .X(_08714_));
 sky130_fd_sc_hd__or2_1 _21457_ (.A(_08542_),
    .B(_08714_),
    .X(_08715_));
 sky130_fd_sc_hd__o211a_1 _21458_ (.A1(_08663_),
    .A2(_08713_),
    .B1(_08715_),
    .C1(_08575_),
    .X(_08716_));
 sky130_fd_sc_hd__mux4_1 _21459_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][4] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][4] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][4] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][4] ),
    .S0(_08567_),
    .S1(_08570_),
    .X(_08717_));
 sky130_fd_sc_hd__mux4_1 _21460_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][4] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][4] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][4] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][4] ),
    .S0(_08649_),
    .S1(_08537_),
    .X(_08718_));
 sky130_fd_sc_hd__or2_1 _21461_ (.A(_08572_),
    .B(_08718_),
    .X(_08719_));
 sky130_fd_sc_hd__o211a_1 _21462_ (.A1(_08565_),
    .A2(_08717_),
    .B1(_08719_),
    .C1(_08652_),
    .X(_08720_));
 sky130_fd_sc_hd__o31a_1 _21463_ (.A1(_08712_),
    .A2(_08716_),
    .A3(_08720_),
    .B1(_08625_),
    .X(_01032_));
 sky130_fd_sc_hd__buf_4 _21464_ (.A(_08559_),
    .X(_08721_));
 sky130_fd_sc_hd__mux4_1 _21465_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][5] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][5] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][5] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][5] ),
    .S0(_08703_),
    .S1(_08721_),
    .X(_08722_));
 sky130_fd_sc_hd__mux4_1 _21466_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][5] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][5] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][5] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][5] ),
    .S0(_08631_),
    .S1(_08632_),
    .X(_08723_));
 sky130_fd_sc_hd__mux2_1 _21467_ (.A0(_08722_),
    .A1(_08723_),
    .S(_08541_),
    .X(_08724_));
 sky130_fd_sc_hd__clkbuf_4 _21468_ (.A(_08531_),
    .X(_08725_));
 sky130_fd_sc_hd__mux4_1 _21469_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][5] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][5] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][5] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][5] ),
    .S0(_08635_),
    .S1(_08637_),
    .X(_08726_));
 sky130_fd_sc_hd__nor2_1 _21470_ (.A(_08725_),
    .B(_08726_),
    .Y(_08727_));
 sky130_fd_sc_hd__mux4_1 _21471_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][5] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][5] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][5] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][5] ),
    .S0(_08517_),
    .S1(_08519_),
    .X(_08728_));
 sky130_fd_sc_hd__o21ai_1 _21472_ (.A1(_08515_),
    .A2(_08728_),
    .B1(_08513_),
    .Y(_08729_));
 sky130_fd_sc_hd__o2bb2a_1 _21473_ (.A1_N(_08627_),
    .A2_N(_08724_),
    .B1(_08727_),
    .B2(_08729_),
    .X(_08730_));
 sky130_fd_sc_hd__nor2_1 _21474_ (.A(_08511_),
    .B(_08730_),
    .Y(_08731_));
 sky130_fd_sc_hd__mux4_1 _21475_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][5] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][5] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][5] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][5] ),
    .S0(_08551_),
    .S1(_08555_),
    .X(_08732_));
 sky130_fd_sc_hd__mux4_1 _21476_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][5] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][5] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][5] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][5] ),
    .S0(_08560_),
    .S1(_08561_),
    .X(_08733_));
 sky130_fd_sc_hd__or2_1 _21477_ (.A(_08542_),
    .B(_08733_),
    .X(_08734_));
 sky130_fd_sc_hd__o211a_1 _21478_ (.A1(_08663_),
    .A2(_08732_),
    .B1(_08734_),
    .C1(_08652_),
    .X(_08735_));
 sky130_fd_sc_hd__mux4_1 _21479_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][5] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][5] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][5] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][5] ),
    .S0(_08567_),
    .S1(_08570_),
    .X(_08736_));
 sky130_fd_sc_hd__mux4_1 _21480_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][5] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][5] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][5] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][5] ),
    .S0(_08566_),
    .S1(_08569_),
    .X(_08737_));
 sky130_fd_sc_hd__or2_1 _21481_ (.A(_08572_),
    .B(_08737_),
    .X(_08738_));
 sky130_fd_sc_hd__o211a_1 _21482_ (.A1(_08565_),
    .A2(_08736_),
    .B1(_08738_),
    .C1(_08576_),
    .X(_08739_));
 sky130_fd_sc_hd__o31a_1 _21483_ (.A1(_08731_),
    .A2(_08735_),
    .A3(_08739_),
    .B1(_08625_),
    .X(_01033_));
 sky130_fd_sc_hd__mux4_1 _21484_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][6] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][6] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][6] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][6] ),
    .S0(_08703_),
    .S1(_08721_),
    .X(_08740_));
 sky130_fd_sc_hd__mux4_1 _21485_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][6] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][6] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][6] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][6] ),
    .S0(_08631_),
    .S1(_08632_),
    .X(_08741_));
 sky130_fd_sc_hd__buf_2 _21486_ (.A(\rvcpu.dp.plfd.InstrD[17] ),
    .X(_08742_));
 sky130_fd_sc_hd__buf_4 _21487_ (.A(_08742_),
    .X(_08743_));
 sky130_fd_sc_hd__mux2_2 _21488_ (.A0(_08740_),
    .A1(_08741_),
    .S(_08743_),
    .X(_08744_));
 sky130_fd_sc_hd__mux4_1 _21489_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][6] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][6] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][6] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][6] ),
    .S0(_08635_),
    .S1(_08637_),
    .X(_08745_));
 sky130_fd_sc_hd__nor2_1 _21490_ (.A(_08725_),
    .B(_08745_),
    .Y(_08746_));
 sky130_fd_sc_hd__mux4_1 _21491_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][6] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][6] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][6] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][6] ),
    .S0(_08517_),
    .S1(_08519_),
    .X(_08747_));
 sky130_fd_sc_hd__buf_2 _21492_ (.A(_08512_),
    .X(_08748_));
 sky130_fd_sc_hd__o21ai_1 _21493_ (.A1(_08515_),
    .A2(_08747_),
    .B1(_08748_),
    .Y(_08749_));
 sky130_fd_sc_hd__o2bb2a_1 _21494_ (.A1_N(_08627_),
    .A2_N(_08744_),
    .B1(_08746_),
    .B2(_08749_),
    .X(_08750_));
 sky130_fd_sc_hd__nor2_1 _21495_ (.A(_08511_),
    .B(_08750_),
    .Y(_08751_));
 sky130_fd_sc_hd__mux4_1 _21496_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][6] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][6] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][6] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][6] ),
    .S0(_08551_),
    .S1(_08555_),
    .X(_08752_));
 sky130_fd_sc_hd__mux4_1 _21497_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][6] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][6] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][6] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][6] ),
    .S0(_08560_),
    .S1(_08561_),
    .X(_08753_));
 sky130_fd_sc_hd__or2_1 _21498_ (.A(_08542_),
    .B(_08753_),
    .X(_08754_));
 sky130_fd_sc_hd__o211a_1 _21499_ (.A1(_08663_),
    .A2(_08752_),
    .B1(_08754_),
    .C1(_08652_),
    .X(_08755_));
 sky130_fd_sc_hd__mux4_1 _21500_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][6] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][6] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][6] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][6] ),
    .S0(_08567_),
    .S1(_08570_),
    .X(_08756_));
 sky130_fd_sc_hd__mux4_1 _21501_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][6] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][6] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][6] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][6] ),
    .S0(_08566_),
    .S1(_08569_),
    .X(_08757_));
 sky130_fd_sc_hd__or2_1 _21502_ (.A(_08572_),
    .B(_08757_),
    .X(_08758_));
 sky130_fd_sc_hd__o211a_1 _21503_ (.A1(_08565_),
    .A2(_08756_),
    .B1(_08758_),
    .C1(_08576_),
    .X(_08759_));
 sky130_fd_sc_hd__o31a_1 _21504_ (.A1(_08751_),
    .A2(_08755_),
    .A3(_08759_),
    .B1(_08625_),
    .X(_01034_));
 sky130_fd_sc_hd__mux4_1 _21505_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][7] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][7] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][7] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][7] ),
    .S0(_08703_),
    .S1(_08721_),
    .X(_08760_));
 sky130_fd_sc_hd__mux4_1 _21506_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][7] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][7] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][7] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][7] ),
    .S0(_08631_),
    .S1(_08632_),
    .X(_08761_));
 sky130_fd_sc_hd__mux2_2 _21507_ (.A0(_08760_),
    .A1(_08761_),
    .S(_08743_),
    .X(_08762_));
 sky130_fd_sc_hd__mux4_1 _21508_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][7] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][7] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][7] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][7] ),
    .S0(_08635_),
    .S1(_08637_),
    .X(_08763_));
 sky130_fd_sc_hd__nor2_1 _21509_ (.A(_08725_),
    .B(_08763_),
    .Y(_08764_));
 sky130_fd_sc_hd__mux4_1 _21510_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][7] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][7] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][7] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][7] ),
    .S0(_08517_),
    .S1(_08519_),
    .X(_08765_));
 sky130_fd_sc_hd__o21ai_1 _21511_ (.A1(_08686_),
    .A2(_08765_),
    .B1(_08748_),
    .Y(_08766_));
 sky130_fd_sc_hd__o2bb2a_1 _21512_ (.A1_N(_08627_),
    .A2_N(_08762_),
    .B1(_08764_),
    .B2(_08766_),
    .X(_08767_));
 sky130_fd_sc_hd__nor2_1 _21513_ (.A(_08511_),
    .B(_08767_),
    .Y(_08768_));
 sky130_fd_sc_hd__mux4_1 _21514_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][7] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][7] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][7] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][7] ),
    .S0(_08551_),
    .S1(_08555_),
    .X(_08769_));
 sky130_fd_sc_hd__mux4_1 _21515_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][7] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][7] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][7] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][7] ),
    .S0(_08550_),
    .S1(_08554_),
    .X(_08770_));
 sky130_fd_sc_hd__or2_1 _21516_ (.A(_08542_),
    .B(_08770_),
    .X(_08771_));
 sky130_fd_sc_hd__o211a_1 _21517_ (.A1(_08663_),
    .A2(_08769_),
    .B1(_08771_),
    .C1(_08575_),
    .X(_08772_));
 sky130_fd_sc_hd__mux4_2 _21518_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][7] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][7] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][7] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][7] ),
    .S0(_08567_),
    .S1(_08570_),
    .X(_08773_));
 sky130_fd_sc_hd__mux4_1 _21519_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][7] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][7] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][7] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][7] ),
    .S0(_08649_),
    .S1(_08537_),
    .X(_08774_));
 sky130_fd_sc_hd__or2_1 _21520_ (.A(_08572_),
    .B(_08774_),
    .X(_08775_));
 sky130_fd_sc_hd__o211a_1 _21521_ (.A1(_08565_),
    .A2(_08773_),
    .B1(_08775_),
    .C1(_08652_),
    .X(_08776_));
 sky130_fd_sc_hd__o31a_1 _21522_ (.A1(_08768_),
    .A2(_08772_),
    .A3(_08776_),
    .B1(_08625_),
    .X(_01035_));
 sky130_fd_sc_hd__mux4_1 _21523_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][8] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][8] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][8] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][8] ),
    .S0(_08703_),
    .S1(_08721_),
    .X(_08777_));
 sky130_fd_sc_hd__clkbuf_8 _21524_ (.A(_08535_),
    .X(_08778_));
 sky130_fd_sc_hd__mux4_1 _21525_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][8] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][8] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][8] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][8] ),
    .S0(_08778_),
    .S1(_08632_),
    .X(_08779_));
 sky130_fd_sc_hd__mux2_2 _21526_ (.A0(_08777_),
    .A1(_08779_),
    .S(_08743_),
    .X(_08780_));
 sky130_fd_sc_hd__mux4_1 _21527_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][8] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][8] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][8] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][8] ),
    .S0(_08635_),
    .S1(_08637_),
    .X(_08781_));
 sky130_fd_sc_hd__nor2_1 _21528_ (.A(_08725_),
    .B(_08781_),
    .Y(_08782_));
 sky130_fd_sc_hd__mux4_1 _21529_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][8] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][8] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][8] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][8] ),
    .S0(_08517_),
    .S1(_08519_),
    .X(_08783_));
 sky130_fd_sc_hd__o21ai_1 _21530_ (.A1(_08686_),
    .A2(_08783_),
    .B1(_08748_),
    .Y(_08784_));
 sky130_fd_sc_hd__o2bb2a_1 _21531_ (.A1_N(_08627_),
    .A2_N(_08780_),
    .B1(_08782_),
    .B2(_08784_),
    .X(_08785_));
 sky130_fd_sc_hd__nor2_1 _21532_ (.A(_08511_),
    .B(_08785_),
    .Y(_08786_));
 sky130_fd_sc_hd__mux4_1 _21533_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][8] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][8] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][8] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][8] ),
    .S0(_08551_),
    .S1(_08555_),
    .X(_08787_));
 sky130_fd_sc_hd__mux4_1 _21534_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][8] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][8] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][8] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][8] ),
    .S0(_08550_),
    .S1(_08554_),
    .X(_08788_));
 sky130_fd_sc_hd__or2_1 _21535_ (.A(_08542_),
    .B(_08788_),
    .X(_08789_));
 sky130_fd_sc_hd__o211a_1 _21536_ (.A1(_08663_),
    .A2(_08787_),
    .B1(_08789_),
    .C1(_08575_),
    .X(_08790_));
 sky130_fd_sc_hd__mux4_2 _21537_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][8] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][8] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][8] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][8] ),
    .S0(_08567_),
    .S1(_08570_),
    .X(_08791_));
 sky130_fd_sc_hd__mux4_1 _21538_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][8] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][8] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][8] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][8] ),
    .S0(_08649_),
    .S1(_08537_),
    .X(_08792_));
 sky130_fd_sc_hd__or2_1 _21539_ (.A(_08572_),
    .B(_08792_),
    .X(_08793_));
 sky130_fd_sc_hd__o211a_1 _21540_ (.A1(_08565_),
    .A2(_08791_),
    .B1(_08793_),
    .C1(_08652_),
    .X(_08794_));
 sky130_fd_sc_hd__o31a_1 _21541_ (.A1(_08786_),
    .A2(_08790_),
    .A3(_08794_),
    .B1(_08625_),
    .X(_01036_));
 sky130_fd_sc_hd__buf_2 _21542_ (.A(_08557_),
    .X(_08795_));
 sky130_fd_sc_hd__mux4_2 _21543_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][9] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][9] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][9] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][9] ),
    .S0(_08524_),
    .S1(_08527_),
    .X(_08796_));
 sky130_fd_sc_hd__or2_1 _21544_ (.A(_08673_),
    .B(_08796_),
    .X(_08797_));
 sky130_fd_sc_hd__buf_2 _21545_ (.A(_08522_),
    .X(_08798_));
 sky130_fd_sc_hd__clkbuf_8 _21546_ (.A(\rvcpu.dp.plfd.InstrD[15] ),
    .X(_08799_));
 sky130_fd_sc_hd__buf_4 _21547_ (.A(_08526_),
    .X(_08800_));
 sky130_fd_sc_hd__mux4_2 _21548_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][9] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][9] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][9] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][9] ),
    .S0(_08799_),
    .S1(_08800_),
    .X(_08801_));
 sky130_fd_sc_hd__or2_1 _21549_ (.A(_08798_),
    .B(_08801_),
    .X(_08802_));
 sky130_fd_sc_hd__mux4_1 _21550_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][9] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][9] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][9] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][9] ),
    .S0(_08559_),
    .S1(_08636_),
    .X(_08803_));
 sky130_fd_sc_hd__mux4_1 _21551_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][9] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][9] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][9] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][9] ),
    .S0(_08548_),
    .S1(_08526_),
    .X(_08804_));
 sky130_fd_sc_hd__or2_1 _21552_ (.A(_08742_),
    .B(_08804_),
    .X(_08805_));
 sky130_fd_sc_hd__clkbuf_4 _21553_ (.A(\rvcpu.dp.plfd.InstrD[18] ),
    .X(_08806_));
 sky130_fd_sc_hd__o211a_1 _21554_ (.A1(_08531_),
    .A2(_08803_),
    .B1(_08805_),
    .C1(_08806_),
    .X(_08807_));
 sky130_fd_sc_hd__clkbuf_4 _21555_ (.A(_08509_),
    .X(_08808_));
 sky130_fd_sc_hd__a311o_1 _21556_ (.A1(_08795_),
    .A2(_08797_),
    .A3(_08802_),
    .B1(_08807_),
    .C1(_08808_),
    .X(_08809_));
 sky130_fd_sc_hd__buf_4 _21557_ (.A(_08628_),
    .X(_08810_));
 sky130_fd_sc_hd__clkbuf_4 _21558_ (.A(_08560_),
    .X(_08811_));
 sky130_fd_sc_hd__mux4_1 _21559_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][9] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][9] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][9] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][9] ),
    .S0(_08810_),
    .S1(_08811_),
    .X(_08812_));
 sky130_fd_sc_hd__clkbuf_4 _21560_ (.A(_08540_),
    .X(_08813_));
 sky130_fd_sc_hd__mux4_1 _21561_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][9] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][9] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][9] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][9] ),
    .S0(_08687_),
    .S1(_08649_),
    .X(_08814_));
 sky130_fd_sc_hd__a21o_1 _21562_ (.A1(_08813_),
    .A2(_08814_),
    .B1(_08689_),
    .X(_08815_));
 sky130_fd_sc_hd__a21o_1 _21563_ (.A1(_08682_),
    .A2(_08812_),
    .B1(_08815_),
    .X(_08816_));
 sky130_fd_sc_hd__clkbuf_4 _21564_ (.A(_08523_),
    .X(_08817_));
 sky130_fd_sc_hd__buf_4 _21565_ (.A(_08525_),
    .X(_08818_));
 sky130_fd_sc_hd__mux4_1 _21566_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][9] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][9] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][9] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][9] ),
    .S0(_08693_),
    .S1(_08818_),
    .X(_08819_));
 sky130_fd_sc_hd__mux4_1 _21567_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][9] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][9] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][9] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][9] ),
    .S0(_08696_),
    .S1(_08568_),
    .X(_08820_));
 sky130_fd_sc_hd__and2_1 _21568_ (.A(_08695_),
    .B(_08820_),
    .X(_08821_));
 sky130_fd_sc_hd__a211o_1 _21569_ (.A1(_08817_),
    .A2(_08819_),
    .B1(_08821_),
    .C1(_08700_),
    .X(_08822_));
 sky130_fd_sc_hd__and4_1 _21570_ (.A(_08672_),
    .B(_08809_),
    .C(_08816_),
    .D(_08822_),
    .X(_08823_));
 sky130_fd_sc_hd__clkbuf_1 _21571_ (.A(_08823_),
    .X(_01037_));
 sky130_fd_sc_hd__mux4_1 _21572_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][10] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][10] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][10] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][10] ),
    .S0(_08703_),
    .S1(_08721_),
    .X(_08824_));
 sky130_fd_sc_hd__buf_4 _21573_ (.A(_08552_),
    .X(_08825_));
 sky130_fd_sc_hd__mux4_1 _21574_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][10] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][10] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][10] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][10] ),
    .S0(_08778_),
    .S1(_08825_),
    .X(_08826_));
 sky130_fd_sc_hd__mux2_2 _21575_ (.A0(_08824_),
    .A1(_08826_),
    .S(_08743_),
    .X(_08827_));
 sky130_fd_sc_hd__mux4_1 _21576_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][10] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][10] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][10] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][10] ),
    .S0(_08629_),
    .S1(_08637_),
    .X(_08828_));
 sky130_fd_sc_hd__nor2_1 _21577_ (.A(_08725_),
    .B(_08828_),
    .Y(_08829_));
 sky130_fd_sc_hd__mux4_1 _21578_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][10] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][10] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][10] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][10] ),
    .S0(_08536_),
    .S1(_08519_),
    .X(_08830_));
 sky130_fd_sc_hd__o21ai_1 _21579_ (.A1(_08686_),
    .A2(_08830_),
    .B1(_08748_),
    .Y(_08831_));
 sky130_fd_sc_hd__o2bb2a_1 _21580_ (.A1_N(_08627_),
    .A2_N(_08827_),
    .B1(_08829_),
    .B2(_08831_),
    .X(_08832_));
 sky130_fd_sc_hd__nor2_1 _21581_ (.A(_08511_),
    .B(_08832_),
    .Y(_08833_));
 sky130_fd_sc_hd__mux4_1 _21582_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][10] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][10] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][10] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][10] ),
    .S0(_08551_),
    .S1(_08555_),
    .X(_08834_));
 sky130_fd_sc_hd__clkbuf_4 _21583_ (.A(_08673_),
    .X(_08835_));
 sky130_fd_sc_hd__mux4_1 _21584_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][10] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][10] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][10] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][10] ),
    .S0(_08550_),
    .S1(_08528_),
    .X(_08836_));
 sky130_fd_sc_hd__or2_1 _21585_ (.A(_08835_),
    .B(_08836_),
    .X(_08837_));
 sky130_fd_sc_hd__o211a_1 _21586_ (.A1(_08663_),
    .A2(_08834_),
    .B1(_08837_),
    .C1(_08575_),
    .X(_08838_));
 sky130_fd_sc_hd__buf_6 _21587_ (.A(_08566_),
    .X(_08839_));
 sky130_fd_sc_hd__clkbuf_8 _21588_ (.A(_08569_),
    .X(_08840_));
 sky130_fd_sc_hd__mux4_1 _21589_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][10] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][10] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][10] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][10] ),
    .S0(_08839_),
    .S1(_08840_),
    .X(_08841_));
 sky130_fd_sc_hd__clkbuf_4 _21590_ (.A(_08673_),
    .X(_08842_));
 sky130_fd_sc_hd__mux4_1 _21591_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][10] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][10] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][10] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][10] ),
    .S0(_08649_),
    .S1(_08537_),
    .X(_08843_));
 sky130_fd_sc_hd__or2_1 _21592_ (.A(_08842_),
    .B(_08843_),
    .X(_08844_));
 sky130_fd_sc_hd__o211a_1 _21593_ (.A1(_08565_),
    .A2(_08841_),
    .B1(_08844_),
    .C1(_08652_),
    .X(_08845_));
 sky130_fd_sc_hd__o31a_1 _21594_ (.A1(_08833_),
    .A2(_08838_),
    .A3(_08845_),
    .B1(_08625_),
    .X(_01038_));
 sky130_fd_sc_hd__mux4_1 _21595_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][11] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][11] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][11] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][11] ),
    .S0(_08524_),
    .S1(_08527_),
    .X(_08846_));
 sky130_fd_sc_hd__or2_1 _21596_ (.A(_08514_),
    .B(_08846_),
    .X(_08847_));
 sky130_fd_sc_hd__mux4_2 _21597_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][11] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][11] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][11] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][11] ),
    .S0(_08799_),
    .S1(_08800_),
    .X(_08848_));
 sky130_fd_sc_hd__or2_1 _21598_ (.A(_08798_),
    .B(_08848_),
    .X(_08849_));
 sky130_fd_sc_hd__mux4_1 _21599_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][11] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][11] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][11] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][11] ),
    .S0(_08559_),
    .S1(_08636_),
    .X(_08850_));
 sky130_fd_sc_hd__mux4_1 _21600_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][11] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][11] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][11] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][11] ),
    .S0(_08548_),
    .S1(_08526_),
    .X(_08851_));
 sky130_fd_sc_hd__or2_1 _21601_ (.A(_08742_),
    .B(_08851_),
    .X(_08852_));
 sky130_fd_sc_hd__o211a_1 _21602_ (.A1(_08531_),
    .A2(_08850_),
    .B1(_08852_),
    .C1(_08806_),
    .X(_08853_));
 sky130_fd_sc_hd__a311o_1 _21603_ (.A1(_08795_),
    .A2(_08847_),
    .A3(_08849_),
    .B1(_08853_),
    .C1(_08808_),
    .X(_08854_));
 sky130_fd_sc_hd__mux4_1 _21604_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][11] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][11] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][11] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][11] ),
    .S0(_08810_),
    .S1(_08811_),
    .X(_08855_));
 sky130_fd_sc_hd__buf_4 _21605_ (.A(_08533_),
    .X(_08856_));
 sky130_fd_sc_hd__mux4_1 _21606_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][11] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][11] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][11] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][11] ),
    .S0(_08687_),
    .S1(_08856_),
    .X(_08857_));
 sky130_fd_sc_hd__a21o_1 _21607_ (.A1(_08813_),
    .A2(_08857_),
    .B1(_08689_),
    .X(_08858_));
 sky130_fd_sc_hd__a21o_1 _21608_ (.A1(_08682_),
    .A2(_08855_),
    .B1(_08858_),
    .X(_08859_));
 sky130_fd_sc_hd__mux4_1 _21609_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][11] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][11] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][11] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][11] ),
    .S0(_08693_),
    .S1(_08818_),
    .X(_08860_));
 sky130_fd_sc_hd__mux4_1 _21610_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][11] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][11] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][11] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][11] ),
    .S0(_08696_),
    .S1(_08568_),
    .X(_08861_));
 sky130_fd_sc_hd__and2_1 _21611_ (.A(_08695_),
    .B(_08861_),
    .X(_08862_));
 sky130_fd_sc_hd__a211o_1 _21612_ (.A1(_08817_),
    .A2(_08860_),
    .B1(_08862_),
    .C1(_08700_),
    .X(_08863_));
 sky130_fd_sc_hd__and4_1 _21613_ (.A(_08672_),
    .B(_08854_),
    .C(_08859_),
    .D(_08863_),
    .X(_08864_));
 sky130_fd_sc_hd__clkbuf_1 _21614_ (.A(_08864_),
    .X(_01039_));
 sky130_fd_sc_hd__mux4_1 _21615_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][12] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][12] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][12] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][12] ),
    .S0(_08516_),
    .S1(_08518_),
    .X(_08865_));
 sky130_fd_sc_hd__mux4_1 _21616_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][12] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][12] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][12] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][12] ),
    .S0(_08516_),
    .S1(_08518_),
    .X(_08866_));
 sky130_fd_sc_hd__mux2_1 _21617_ (.A0(_08865_),
    .A1(_08866_),
    .S(_08540_),
    .X(_08867_));
 sky130_fd_sc_hd__mux4_1 _21618_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][12] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][12] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][12] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][12] ),
    .S0(_08549_),
    .S1(_08553_),
    .X(_08868_));
 sky130_fd_sc_hd__or2_1 _21619_ (.A(_08673_),
    .B(_08868_),
    .X(_08869_));
 sky130_fd_sc_hd__mux4_1 _21620_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][12] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][12] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][12] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][12] ),
    .S0(_08533_),
    .S1(_08536_),
    .X(_08870_));
 sky130_fd_sc_hd__o21a_1 _21621_ (.A1(_08531_),
    .A2(_08870_),
    .B1(_08806_),
    .X(_08871_));
 sky130_fd_sc_hd__a221o_1 _21622_ (.A1(_08626_),
    .A2(_08867_),
    .B1(_08869_),
    .B2(_08871_),
    .C1(_08808_),
    .X(_08872_));
 sky130_fd_sc_hd__mux4_2 _21623_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][12] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][12] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][12] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][12] ),
    .S0(_08534_),
    .S1(_08537_),
    .X(_08873_));
 sky130_fd_sc_hd__mux4_1 _21624_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][12] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][12] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][12] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][12] ),
    .S0(_08549_),
    .S1(_08553_),
    .X(_08874_));
 sky130_fd_sc_hd__and2_1 _21625_ (.A(_08541_),
    .B(_08874_),
    .X(_08875_));
 sky130_fd_sc_hd__a211o_1 _21626_ (.A1(_08532_),
    .A2(_08873_),
    .B1(_08875_),
    .C1(_08699_),
    .X(_08876_));
 sky130_fd_sc_hd__mux4_1 _21627_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][12] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][12] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][12] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][12] ),
    .S0(_08683_),
    .S1(_08684_),
    .X(_08877_));
 sky130_fd_sc_hd__mux4_1 _21628_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][12] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][12] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][12] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][12] ),
    .S0(_08687_),
    .S1(_08649_),
    .X(_08878_));
 sky130_fd_sc_hd__a21o_1 _21629_ (.A1(_08686_),
    .A2(_08878_),
    .B1(_08689_),
    .X(_08879_));
 sky130_fd_sc_hd__a21o_1 _21630_ (.A1(_08682_),
    .A2(_08877_),
    .B1(_08879_),
    .X(_08880_));
 sky130_fd_sc_hd__and4_1 _21631_ (.A(_08672_),
    .B(_08872_),
    .C(_08876_),
    .D(_08880_),
    .X(_08881_));
 sky130_fd_sc_hd__clkbuf_1 _21632_ (.A(_08881_),
    .X(_01040_));
 sky130_fd_sc_hd__mux4_1 _21633_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][13] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][13] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][13] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][13] ),
    .S0(_08524_),
    .S1(_08800_),
    .X(_08882_));
 sky130_fd_sc_hd__or2_1 _21634_ (.A(_08514_),
    .B(_08882_),
    .X(_08883_));
 sky130_fd_sc_hd__mux4_2 _21635_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][13] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][13] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][13] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][13] ),
    .S0(_08799_),
    .S1(_08800_),
    .X(_08884_));
 sky130_fd_sc_hd__or2_1 _21636_ (.A(_08798_),
    .B(_08884_),
    .X(_08885_));
 sky130_fd_sc_hd__mux4_1 _21637_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][13] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][13] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][13] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][13] ),
    .S0(_08559_),
    .S1(_08636_),
    .X(_08886_));
 sky130_fd_sc_hd__mux4_1 _21638_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][13] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][13] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][13] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][13] ),
    .S0(_08548_),
    .S1(_08526_),
    .X(_08887_));
 sky130_fd_sc_hd__or2_1 _21639_ (.A(_08742_),
    .B(_08887_),
    .X(_08888_));
 sky130_fd_sc_hd__o211a_1 _21640_ (.A1(_08531_),
    .A2(_08886_),
    .B1(_08888_),
    .C1(_08806_),
    .X(_08889_));
 sky130_fd_sc_hd__a311o_1 _21641_ (.A1(_08795_),
    .A2(_08883_),
    .A3(_08885_),
    .B1(_08889_),
    .C1(_08808_),
    .X(_08890_));
 sky130_fd_sc_hd__mux4_1 _21642_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][13] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][13] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][13] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][13] ),
    .S0(_08810_),
    .S1(_08811_),
    .X(_08891_));
 sky130_fd_sc_hd__mux4_1 _21643_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][13] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][13] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][13] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][13] ),
    .S0(_08687_),
    .S1(_08856_),
    .X(_08892_));
 sky130_fd_sc_hd__a21o_1 _21644_ (.A1(_08813_),
    .A2(_08892_),
    .B1(_08689_),
    .X(_08893_));
 sky130_fd_sc_hd__a21o_1 _21645_ (.A1(_08692_),
    .A2(_08891_),
    .B1(_08893_),
    .X(_08894_));
 sky130_fd_sc_hd__mux4_1 _21646_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][13] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][13] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][13] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][13] ),
    .S0(_08693_),
    .S1(_08818_),
    .X(_08895_));
 sky130_fd_sc_hd__mux4_1 _21647_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][13] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][13] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][13] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][13] ),
    .S0(_08696_),
    .S1(_08568_),
    .X(_08896_));
 sky130_fd_sc_hd__and2_1 _21648_ (.A(_08695_),
    .B(_08896_),
    .X(_08897_));
 sky130_fd_sc_hd__a211o_1 _21649_ (.A1(_08817_),
    .A2(_08895_),
    .B1(_08897_),
    .C1(_08700_),
    .X(_08898_));
 sky130_fd_sc_hd__and4_1 _21650_ (.A(_08672_),
    .B(_08890_),
    .C(_08894_),
    .D(_08898_),
    .X(_08899_));
 sky130_fd_sc_hd__clkbuf_1 _21651_ (.A(_08899_),
    .X(_01041_));
 sky130_fd_sc_hd__mux4_1 _21652_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][14] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][14] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][14] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][14] ),
    .S0(_08524_),
    .S1(_08527_),
    .X(_08900_));
 sky130_fd_sc_hd__or2_1 _21653_ (.A(_08673_),
    .B(_08900_),
    .X(_08901_));
 sky130_fd_sc_hd__mux4_1 _21654_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][14] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][14] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][14] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][14] ),
    .S0(_08533_),
    .S1(_08636_),
    .X(_08902_));
 sky130_fd_sc_hd__o21a_1 _21655_ (.A1(_08531_),
    .A2(_08902_),
    .B1(_08512_),
    .X(_08903_));
 sky130_fd_sc_hd__mux4_1 _21656_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][14] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][14] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][14] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][14] ),
    .S0(_08524_),
    .S1(_08527_),
    .X(_08904_));
 sky130_fd_sc_hd__mux4_1 _21657_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][14] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][14] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][14] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][14] ),
    .S0(_08524_),
    .S1(_08527_),
    .X(_08905_));
 sky130_fd_sc_hd__mux2_1 _21658_ (.A0(_08904_),
    .A1(_08905_),
    .S(_08540_),
    .X(_08906_));
 sky130_fd_sc_hd__a221o_1 _21659_ (.A1(_08901_),
    .A2(_08903_),
    .B1(_08906_),
    .B2(_08626_),
    .C1(_08808_),
    .X(_08907_));
 sky130_fd_sc_hd__mux4_1 _21660_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][14] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][14] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][14] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][14] ),
    .S0(_08810_),
    .S1(_08811_),
    .X(_08908_));
 sky130_fd_sc_hd__mux4_1 _21661_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][14] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][14] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][14] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][14] ),
    .S0(_08687_),
    .S1(_08856_),
    .X(_08909_));
 sky130_fd_sc_hd__a21o_1 _21662_ (.A1(_08813_),
    .A2(_08909_),
    .B1(_08689_),
    .X(_08910_));
 sky130_fd_sc_hd__a21o_1 _21663_ (.A1(_08692_),
    .A2(_08908_),
    .B1(_08910_),
    .X(_08911_));
 sky130_fd_sc_hd__mux4_2 _21664_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][14] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][14] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][14] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][14] ),
    .S0(_08693_),
    .S1(_08818_),
    .X(_08912_));
 sky130_fd_sc_hd__mux4_1 _21665_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][14] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][14] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][14] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][14] ),
    .S0(_08696_),
    .S1(_08568_),
    .X(_08913_));
 sky130_fd_sc_hd__and2_1 _21666_ (.A(_08695_),
    .B(_08913_),
    .X(_08914_));
 sky130_fd_sc_hd__a211o_1 _21667_ (.A1(_08817_),
    .A2(_08912_),
    .B1(_08914_),
    .C1(_08700_),
    .X(_08915_));
 sky130_fd_sc_hd__and4_1 _21668_ (.A(_08672_),
    .B(_08907_),
    .C(_08911_),
    .D(_08915_),
    .X(_08916_));
 sky130_fd_sc_hd__clkbuf_1 _21669_ (.A(_08916_),
    .X(_01042_));
 sky130_fd_sc_hd__mux4_2 _21670_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][15] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][15] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][15] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][15] ),
    .S0(_08799_),
    .S1(_08800_),
    .X(_08917_));
 sky130_fd_sc_hd__or2_1 _21671_ (.A(_08514_),
    .B(_08917_),
    .X(_08918_));
 sky130_fd_sc_hd__mux4_2 _21672_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][15] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][15] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][15] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][15] ),
    .S0(_08799_),
    .S1(_08800_),
    .X(_08919_));
 sky130_fd_sc_hd__or2_1 _21673_ (.A(_08798_),
    .B(_08919_),
    .X(_08920_));
 sky130_fd_sc_hd__mux4_1 _21674_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][15] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][15] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][15] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][15] ),
    .S0(_08559_),
    .S1(_08636_),
    .X(_08921_));
 sky130_fd_sc_hd__mux4_1 _21675_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][15] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][15] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][15] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][15] ),
    .S0(_08548_),
    .S1(_08526_),
    .X(_08922_));
 sky130_fd_sc_hd__or2_1 _21676_ (.A(_08742_),
    .B(_08922_),
    .X(_08923_));
 sky130_fd_sc_hd__o211a_1 _21677_ (.A1(_08798_),
    .A2(_08921_),
    .B1(_08923_),
    .C1(_08806_),
    .X(_08924_));
 sky130_fd_sc_hd__a311o_1 _21678_ (.A1(_08795_),
    .A2(_08918_),
    .A3(_08920_),
    .B1(_08924_),
    .C1(_08808_),
    .X(_08925_));
 sky130_fd_sc_hd__mux4_1 _21679_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][15] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][15] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][15] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][15] ),
    .S0(_08810_),
    .S1(_08811_),
    .X(_08926_));
 sky130_fd_sc_hd__mux4_1 _21680_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][15] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][15] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][15] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][15] ),
    .S0(_08687_),
    .S1(_08856_),
    .X(_08927_));
 sky130_fd_sc_hd__a21o_1 _21681_ (.A1(_08813_),
    .A2(_08927_),
    .B1(_08689_),
    .X(_08928_));
 sky130_fd_sc_hd__a21o_1 _21682_ (.A1(_08692_),
    .A2(_08926_),
    .B1(_08928_),
    .X(_08929_));
 sky130_fd_sc_hd__mux4_1 _21683_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][15] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][15] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][15] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][15] ),
    .S0(_08534_),
    .S1(_08818_),
    .X(_08930_));
 sky130_fd_sc_hd__mux4_1 _21684_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][15] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][15] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][15] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][15] ),
    .S0(_08696_),
    .S1(_08568_),
    .X(_08931_));
 sky130_fd_sc_hd__and2_1 _21685_ (.A(_08695_),
    .B(_08931_),
    .X(_08932_));
 sky130_fd_sc_hd__a211o_1 _21686_ (.A1(_08817_),
    .A2(_08930_),
    .B1(_08932_),
    .C1(_08700_),
    .X(_08933_));
 sky130_fd_sc_hd__and4_1 _21687_ (.A(_08672_),
    .B(_08925_),
    .C(_08929_),
    .D(_08933_),
    .X(_08934_));
 sky130_fd_sc_hd__clkbuf_1 _21688_ (.A(_08934_),
    .X(_01043_));
 sky130_fd_sc_hd__mux4_1 _21689_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][16] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][16] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][16] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][16] ),
    .S0(_08703_),
    .S1(_08721_),
    .X(_08935_));
 sky130_fd_sc_hd__mux4_1 _21690_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][16] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][16] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][16] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][16] ),
    .S0(_08778_),
    .S1(_08825_),
    .X(_08936_));
 sky130_fd_sc_hd__mux2_1 _21691_ (.A0(_08935_),
    .A1(_08936_),
    .S(_08743_),
    .X(_08937_));
 sky130_fd_sc_hd__mux4_1 _21692_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][16] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][16] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][16] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][16] ),
    .S0(_08525_),
    .S1(_08528_),
    .X(_08938_));
 sky130_fd_sc_hd__nor2_1 _21693_ (.A(_08515_),
    .B(_08938_),
    .Y(_08939_));
 sky130_fd_sc_hd__mux4_1 _21694_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][16] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][16] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][16] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][16] ),
    .S0(_08568_),
    .S1(_08683_),
    .X(_08940_));
 sky130_fd_sc_hd__o21ai_1 _21695_ (.A1(_08523_),
    .A2(_08940_),
    .B1(_08748_),
    .Y(_08941_));
 sky130_fd_sc_hd__o2bb2a_1 _21696_ (.A1_N(_08627_),
    .A2_N(_08937_),
    .B1(_08939_),
    .B2(_08941_),
    .X(_08942_));
 sky130_fd_sc_hd__nor2_1 _21697_ (.A(_08511_),
    .B(_08942_),
    .Y(_08943_));
 sky130_fd_sc_hd__mux4_1 _21698_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][16] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][16] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][16] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][16] ),
    .S0(_08551_),
    .S1(_08555_),
    .X(_08944_));
 sky130_fd_sc_hd__mux4_1 _21699_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][16] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][16] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][16] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][16] ),
    .S0(_08560_),
    .S1(_08561_),
    .X(_08945_));
 sky130_fd_sc_hd__or2_1 _21700_ (.A(_08835_),
    .B(_08945_),
    .X(_08946_));
 sky130_fd_sc_hd__o211a_1 _21701_ (.A1(_08663_),
    .A2(_08944_),
    .B1(_08946_),
    .C1(_08558_),
    .X(_08947_));
 sky130_fd_sc_hd__mux4_1 _21702_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][16] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][16] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][16] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][16] ),
    .S0(_08839_),
    .S1(_08840_),
    .X(_08948_));
 sky130_fd_sc_hd__mux4_1 _21703_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][16] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][16] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][16] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][16] ),
    .S0(_08566_),
    .S1(_08569_),
    .X(_08949_));
 sky130_fd_sc_hd__or2_1 _21704_ (.A(_08842_),
    .B(_08949_),
    .X(_08950_));
 sky130_fd_sc_hd__o211a_1 _21705_ (.A1(_08565_),
    .A2(_08948_),
    .B1(_08950_),
    .C1(_08576_),
    .X(_08951_));
 sky130_fd_sc_hd__o31a_1 _21706_ (.A1(_08943_),
    .A2(_08947_),
    .A3(_08951_),
    .B1(_08625_),
    .X(_01044_));
 sky130_fd_sc_hd__mux4_1 _21707_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][17] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][17] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][17] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][17] ),
    .S0(_08703_),
    .S1(_08721_),
    .X(_08952_));
 sky130_fd_sc_hd__mux4_1 _21708_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][17] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][17] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][17] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][17] ),
    .S0(_08778_),
    .S1(_08825_),
    .X(_08953_));
 sky130_fd_sc_hd__mux2_1 _21709_ (.A0(_08952_),
    .A1(_08953_),
    .S(_08743_),
    .X(_08954_));
 sky130_fd_sc_hd__mux4_1 _21710_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][17] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][17] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][17] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][17] ),
    .S0(_08629_),
    .S1(_08683_),
    .X(_08955_));
 sky130_fd_sc_hd__nor2_1 _21711_ (.A(_08725_),
    .B(_08955_),
    .Y(_08956_));
 sky130_fd_sc_hd__mux4_1 _21712_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][17] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][17] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][17] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][17] ),
    .S0(_08536_),
    .S1(_08693_),
    .X(_08957_));
 sky130_fd_sc_hd__o21ai_1 _21713_ (.A1(_08686_),
    .A2(_08957_),
    .B1(_08748_),
    .Y(_08958_));
 sky130_fd_sc_hd__o2bb2a_1 _21714_ (.A1_N(_08627_),
    .A2_N(_08954_),
    .B1(_08956_),
    .B2(_08958_),
    .X(_08959_));
 sky130_fd_sc_hd__nor2_1 _21715_ (.A(_08510_),
    .B(_08959_),
    .Y(_08960_));
 sky130_fd_sc_hd__mux4_1 _21716_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][17] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][17] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][17] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][17] ),
    .S0(_08578_),
    .S1(_08684_),
    .X(_08961_));
 sky130_fd_sc_hd__mux4_1 _21717_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][17] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][17] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][17] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][17] ),
    .S0(_08525_),
    .S1(_08528_),
    .X(_08962_));
 sky130_fd_sc_hd__or2_1 _21718_ (.A(_08835_),
    .B(_08962_),
    .X(_08963_));
 sky130_fd_sc_hd__o211a_1 _21719_ (.A1(_08663_),
    .A2(_08961_),
    .B1(_08963_),
    .C1(_08575_),
    .X(_08964_));
 sky130_fd_sc_hd__mux4_2 _21720_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][17] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][17] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][17] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][17] ),
    .S0(_08839_),
    .S1(_08840_),
    .X(_08965_));
 sky130_fd_sc_hd__mux4_2 _21721_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][17] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][17] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][17] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][17] ),
    .S0(_08649_),
    .S1(_08537_),
    .X(_08966_));
 sky130_fd_sc_hd__or2_1 _21722_ (.A(_08842_),
    .B(_08966_),
    .X(_08967_));
 sky130_fd_sc_hd__o211a_1 _21723_ (.A1(_08547_),
    .A2(_08965_),
    .B1(_08967_),
    .C1(_08652_),
    .X(_08968_));
 sky130_fd_sc_hd__o31a_1 _21724_ (.A1(_08960_),
    .A2(_08964_),
    .A3(_08968_),
    .B1(_08624_),
    .X(_01045_));
 sky130_fd_sc_hd__mux4_1 _21725_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][18] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][18] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][18] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][18] ),
    .S0(_08703_),
    .S1(_08721_),
    .X(_08969_));
 sky130_fd_sc_hd__mux4_1 _21726_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][18] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][18] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][18] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][18] ),
    .S0(_08778_),
    .S1(_08825_),
    .X(_08970_));
 sky130_fd_sc_hd__mux2_2 _21727_ (.A0(_08969_),
    .A1(_08970_),
    .S(_08743_),
    .X(_08971_));
 sky130_fd_sc_hd__mux4_1 _21728_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][18] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][18] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][18] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][18] ),
    .S0(_08629_),
    .S1(_08683_),
    .X(_08972_));
 sky130_fd_sc_hd__nor2_1 _21729_ (.A(_08725_),
    .B(_08972_),
    .Y(_08973_));
 sky130_fd_sc_hd__mux4_1 _21730_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][18] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][18] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][18] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][18] ),
    .S0(_08536_),
    .S1(_08693_),
    .X(_08974_));
 sky130_fd_sc_hd__o21ai_1 _21731_ (.A1(_08686_),
    .A2(_08974_),
    .B1(_08748_),
    .Y(_08975_));
 sky130_fd_sc_hd__o2bb2a_1 _21732_ (.A1_N(_08795_),
    .A2_N(_08971_),
    .B1(_08973_),
    .B2(_08975_),
    .X(_08976_));
 sky130_fd_sc_hd__nor2_1 _21733_ (.A(_08510_),
    .B(_08976_),
    .Y(_08977_));
 sky130_fd_sc_hd__mux4_1 _21734_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][18] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][18] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][18] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][18] ),
    .S0(_08578_),
    .S1(_08684_),
    .X(_08978_));
 sky130_fd_sc_hd__mux4_1 _21735_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][18] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][18] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][18] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][18] ),
    .S0(_08560_),
    .S1(_08561_),
    .X(_08979_));
 sky130_fd_sc_hd__or2_1 _21736_ (.A(_08835_),
    .B(_08979_),
    .X(_08980_));
 sky130_fd_sc_hd__o211a_1 _21737_ (.A1(_08663_),
    .A2(_08978_),
    .B1(_08980_),
    .C1(_08558_),
    .X(_08981_));
 sky130_fd_sc_hd__mux4_1 _21738_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][18] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][18] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][18] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][18] ),
    .S0(_08839_),
    .S1(_08840_),
    .X(_08982_));
 sky130_fd_sc_hd__mux4_1 _21739_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][18] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][18] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][18] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][18] ),
    .S0(_08566_),
    .S1(_08569_),
    .X(_08983_));
 sky130_fd_sc_hd__or2_1 _21740_ (.A(_08842_),
    .B(_08983_),
    .X(_08984_));
 sky130_fd_sc_hd__o211a_1 _21741_ (.A1(_08547_),
    .A2(_08982_),
    .B1(_08984_),
    .C1(_08576_),
    .X(_08985_));
 sky130_fd_sc_hd__o31a_1 _21742_ (.A1(_08977_),
    .A2(_08981_),
    .A3(_08985_),
    .B1(_08624_),
    .X(_01046_));
 sky130_fd_sc_hd__mux4_2 _21743_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][19] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][19] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][19] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][19] ),
    .S0(_08799_),
    .S1(_08800_),
    .X(_08986_));
 sky130_fd_sc_hd__or2_1 _21744_ (.A(_08514_),
    .B(_08986_),
    .X(_08987_));
 sky130_fd_sc_hd__mux4_2 _21745_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][19] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][19] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][19] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][19] ),
    .S0(_08799_),
    .S1(_08518_),
    .X(_08988_));
 sky130_fd_sc_hd__or2_1 _21746_ (.A(_08798_),
    .B(_08988_),
    .X(_08989_));
 sky130_fd_sc_hd__mux4_1 _21747_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][19] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][19] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][19] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][19] ),
    .S0(_08559_),
    .S1(_08636_),
    .X(_08990_));
 sky130_fd_sc_hd__mux4_1 _21748_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][19] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][19] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][19] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][19] ),
    .S0(_08548_),
    .S1(_08526_),
    .X(_08991_));
 sky130_fd_sc_hd__or2_1 _21749_ (.A(_08742_),
    .B(_08991_),
    .X(_08992_));
 sky130_fd_sc_hd__o211a_1 _21750_ (.A1(_08798_),
    .A2(_08990_),
    .B1(_08992_),
    .C1(_08806_),
    .X(_08993_));
 sky130_fd_sc_hd__a311o_1 _21751_ (.A1(_08626_),
    .A2(_08987_),
    .A3(_08989_),
    .B1(_08993_),
    .C1(_08808_),
    .X(_08994_));
 sky130_fd_sc_hd__mux4_1 _21752_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][19] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][19] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][19] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][19] ),
    .S0(_08810_),
    .S1(_08811_),
    .X(_08995_));
 sky130_fd_sc_hd__mux4_1 _21753_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][19] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][19] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][19] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][19] ),
    .S0(_08687_),
    .S1(_08856_),
    .X(_08996_));
 sky130_fd_sc_hd__a21o_1 _21754_ (.A1(_08813_),
    .A2(_08996_),
    .B1(_08689_),
    .X(_08997_));
 sky130_fd_sc_hd__a21o_1 _21755_ (.A1(_08692_),
    .A2(_08995_),
    .B1(_08997_),
    .X(_08998_));
 sky130_fd_sc_hd__mux4_1 _21756_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][19] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][19] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][19] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][19] ),
    .S0(_08534_),
    .S1(_08818_),
    .X(_08999_));
 sky130_fd_sc_hd__mux4_1 _21757_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][19] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][19] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][19] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][19] ),
    .S0(_08696_),
    .S1(_08553_),
    .X(_09000_));
 sky130_fd_sc_hd__and2_1 _21758_ (.A(_08695_),
    .B(_09000_),
    .X(_09001_));
 sky130_fd_sc_hd__a211o_1 _21759_ (.A1(_08817_),
    .A2(_08999_),
    .B1(_09001_),
    .C1(_08700_),
    .X(_09002_));
 sky130_fd_sc_hd__and4_1 _21760_ (.A(_08672_),
    .B(_08994_),
    .C(_08998_),
    .D(_09002_),
    .X(_09003_));
 sky130_fd_sc_hd__clkbuf_1 _21761_ (.A(_09003_),
    .X(_01047_));
 sky130_fd_sc_hd__mux4_1 _21762_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][20] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][20] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][20] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][20] ),
    .S0(_08799_),
    .S1(_08800_),
    .X(_09004_));
 sky130_fd_sc_hd__or2_1 _21763_ (.A(_08514_),
    .B(_09004_),
    .X(_09005_));
 sky130_fd_sc_hd__mux4_2 _21764_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][20] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][20] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][20] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][20] ),
    .S0(_08516_),
    .S1(_08518_),
    .X(_09006_));
 sky130_fd_sc_hd__or2_1 _21765_ (.A(_08522_),
    .B(_09006_),
    .X(_09007_));
 sky130_fd_sc_hd__mux4_1 _21766_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][20] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][20] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][20] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][20] ),
    .S0(_08559_),
    .S1(_08636_),
    .X(_09008_));
 sky130_fd_sc_hd__mux4_1 _21767_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][20] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][20] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][20] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][20] ),
    .S0(_08548_),
    .S1(_08526_),
    .X(_09009_));
 sky130_fd_sc_hd__or2_1 _21768_ (.A(_08742_),
    .B(_09009_),
    .X(_09010_));
 sky130_fd_sc_hd__o211a_1 _21769_ (.A1(_08798_),
    .A2(_09008_),
    .B1(_09010_),
    .C1(_08512_),
    .X(_09011_));
 sky130_fd_sc_hd__a311o_1 _21770_ (.A1(_08626_),
    .A2(_09005_),
    .A3(_09007_),
    .B1(_09011_),
    .C1(_08808_),
    .X(_09012_));
 sky130_fd_sc_hd__mux4_1 _21771_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][20] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][20] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][20] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][20] ),
    .S0(_08810_),
    .S1(_08811_),
    .X(_09013_));
 sky130_fd_sc_hd__mux4_1 _21772_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][20] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][20] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][20] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][20] ),
    .S0(_08628_),
    .S1(_08856_),
    .X(_09014_));
 sky130_fd_sc_hd__a21o_1 _21773_ (.A1(_08813_),
    .A2(_09014_),
    .B1(_08689_),
    .X(_09015_));
 sky130_fd_sc_hd__a21o_1 _21774_ (.A1(_08692_),
    .A2(_09013_),
    .B1(_09015_),
    .X(_09016_));
 sky130_fd_sc_hd__mux4_1 _21775_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][20] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][20] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][20] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][20] ),
    .S0(_08534_),
    .S1(_08818_),
    .X(_09017_));
 sky130_fd_sc_hd__mux4_1 _21776_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][20] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][20] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][20] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][20] ),
    .S0(_08696_),
    .S1(_08553_),
    .X(_09018_));
 sky130_fd_sc_hd__and2_1 _21777_ (.A(_08695_),
    .B(_09018_),
    .X(_09019_));
 sky130_fd_sc_hd__a211o_1 _21778_ (.A1(_08817_),
    .A2(_09017_),
    .B1(_09019_),
    .C1(_08700_),
    .X(_09020_));
 sky130_fd_sc_hd__and4_1 _21779_ (.A(_08672_),
    .B(_09012_),
    .C(_09016_),
    .D(_09020_),
    .X(_09021_));
 sky130_fd_sc_hd__clkbuf_1 _21780_ (.A(_09021_),
    .X(_01048_));
 sky130_fd_sc_hd__mux4_1 _21781_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][21] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][21] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][21] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][21] ),
    .S0(_08703_),
    .S1(_08721_),
    .X(_09022_));
 sky130_fd_sc_hd__mux4_1 _21782_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][21] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][21] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][21] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][21] ),
    .S0(_08778_),
    .S1(_08825_),
    .X(_09023_));
 sky130_fd_sc_hd__mux2_1 _21783_ (.A0(_09022_),
    .A1(_09023_),
    .S(_08743_),
    .X(_09024_));
 sky130_fd_sc_hd__mux4_1 _21784_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][21] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][21] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][21] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][21] ),
    .S0(_08629_),
    .S1(_08683_),
    .X(_09025_));
 sky130_fd_sc_hd__nor2_1 _21785_ (.A(_08725_),
    .B(_09025_),
    .Y(_09026_));
 sky130_fd_sc_hd__mux4_1 _21786_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][21] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][21] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][21] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][21] ),
    .S0(_08536_),
    .S1(_08693_),
    .X(_09027_));
 sky130_fd_sc_hd__o21ai_1 _21787_ (.A1(_08686_),
    .A2(_09027_),
    .B1(_08748_),
    .Y(_09028_));
 sky130_fd_sc_hd__o2bb2a_1 _21788_ (.A1_N(_08795_),
    .A2_N(_09024_),
    .B1(_09026_),
    .B2(_09028_),
    .X(_09029_));
 sky130_fd_sc_hd__nor2_1 _21789_ (.A(_08510_),
    .B(_09029_),
    .Y(_09030_));
 sky130_fd_sc_hd__mux4_1 _21790_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][21] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][21] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][21] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][21] ),
    .S0(_08578_),
    .S1(_08684_),
    .X(_09031_));
 sky130_fd_sc_hd__mux4_1 _21791_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][21] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][21] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][21] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][21] ),
    .S0(_08560_),
    .S1(_08561_),
    .X(_09032_));
 sky130_fd_sc_hd__or2_1 _21792_ (.A(_08835_),
    .B(_09032_),
    .X(_09033_));
 sky130_fd_sc_hd__o211a_1 _21793_ (.A1(_08682_),
    .A2(_09031_),
    .B1(_09033_),
    .C1(_08558_),
    .X(_09034_));
 sky130_fd_sc_hd__mux4_1 _21794_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][21] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][21] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][21] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][21] ),
    .S0(_08839_),
    .S1(_08840_),
    .X(_09035_));
 sky130_fd_sc_hd__mux4_1 _21795_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][21] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][21] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][21] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][21] ),
    .S0(_08566_),
    .S1(_08554_),
    .X(_09036_));
 sky130_fd_sc_hd__or2_1 _21796_ (.A(_08842_),
    .B(_09036_),
    .X(_09037_));
 sky130_fd_sc_hd__o211a_1 _21797_ (.A1(_08547_),
    .A2(_09035_),
    .B1(_09037_),
    .C1(_08576_),
    .X(_09038_));
 sky130_fd_sc_hd__o31a_1 _21798_ (.A1(_09030_),
    .A2(_09034_),
    .A3(_09038_),
    .B1(_08624_),
    .X(_01049_));
 sky130_fd_sc_hd__mux4_1 _21799_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][22] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][22] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][22] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][22] ),
    .S0(_08799_),
    .S1(_08800_),
    .X(_09039_));
 sky130_fd_sc_hd__or2_1 _21800_ (.A(_08514_),
    .B(_09039_),
    .X(_09040_));
 sky130_fd_sc_hd__mux4_1 _21801_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][22] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][22] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][22] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][22] ),
    .S0(_08516_),
    .S1(_08518_),
    .X(_09041_));
 sky130_fd_sc_hd__or2_1 _21802_ (.A(_08522_),
    .B(_09041_),
    .X(_09042_));
 sky130_fd_sc_hd__mux4_1 _21803_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][22] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][22] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][22] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][22] ),
    .S0(_08552_),
    .S1(_08687_),
    .X(_09043_));
 sky130_fd_sc_hd__mux4_1 _21804_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][22] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][22] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][22] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][22] ),
    .S0(\rvcpu.dp.plfd.InstrD[15] ),
    .S1(_08526_),
    .X(_09044_));
 sky130_fd_sc_hd__or2_1 _21805_ (.A(_08742_),
    .B(_09044_),
    .X(_09045_));
 sky130_fd_sc_hd__o211a_1 _21806_ (.A1(_08798_),
    .A2(_09043_),
    .B1(_09045_),
    .C1(_08512_),
    .X(_09046_));
 sky130_fd_sc_hd__a311o_1 _21807_ (.A1(_08626_),
    .A2(_09040_),
    .A3(_09042_),
    .B1(_09046_),
    .C1(_08509_),
    .X(_09047_));
 sky130_fd_sc_hd__mux4_1 _21808_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][22] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][22] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][22] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][22] ),
    .S0(_08810_),
    .S1(_08811_),
    .X(_09048_));
 sky130_fd_sc_hd__mux4_1 _21809_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][22] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][22] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][22] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][22] ),
    .S0(_08628_),
    .S1(_08856_),
    .X(_09049_));
 sky130_fd_sc_hd__a21o_1 _21810_ (.A1(_08813_),
    .A2(_09049_),
    .B1(_08689_),
    .X(_09050_));
 sky130_fd_sc_hd__a21o_1 _21811_ (.A1(_08692_),
    .A2(_09048_),
    .B1(_09050_),
    .X(_09051_));
 sky130_fd_sc_hd__mux4_1 _21812_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][22] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][22] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][22] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][22] ),
    .S0(_08534_),
    .S1(_08818_),
    .X(_09052_));
 sky130_fd_sc_hd__mux4_1 _21813_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][22] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][22] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][22] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][22] ),
    .S0(_08696_),
    .S1(_08553_),
    .X(_09053_));
 sky130_fd_sc_hd__and2_1 _21814_ (.A(_08695_),
    .B(_09053_),
    .X(_09054_));
 sky130_fd_sc_hd__a211o_1 _21815_ (.A1(_08817_),
    .A2(_09052_),
    .B1(_09054_),
    .C1(_08700_),
    .X(_09055_));
 sky130_fd_sc_hd__and4_1 _21816_ (.A(_08672_),
    .B(_09047_),
    .C(_09051_),
    .D(_09055_),
    .X(_09056_));
 sky130_fd_sc_hd__clkbuf_1 _21817_ (.A(_09056_),
    .X(_01050_));
 sky130_fd_sc_hd__mux4_1 _21818_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][23] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][23] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][23] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][23] ),
    .S0(_08631_),
    .S1(_08721_),
    .X(_09057_));
 sky130_fd_sc_hd__mux4_1 _21819_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][23] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][23] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][23] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][23] ),
    .S0(_08778_),
    .S1(_08825_),
    .X(_09058_));
 sky130_fd_sc_hd__mux2_1 _21820_ (.A0(_09057_),
    .A1(_09058_),
    .S(_08743_),
    .X(_09059_));
 sky130_fd_sc_hd__mux4_1 _21821_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][23] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][23] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][23] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][23] ),
    .S0(_08525_),
    .S1(_08528_),
    .X(_09060_));
 sky130_fd_sc_hd__nor2_1 _21822_ (.A(_08515_),
    .B(_09060_),
    .Y(_09061_));
 sky130_fd_sc_hd__mux4_1 _21823_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][23] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][23] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][23] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][23] ),
    .S0(_08568_),
    .S1(_08683_),
    .X(_09062_));
 sky130_fd_sc_hd__o21ai_1 _21824_ (.A1(_08523_),
    .A2(_09062_),
    .B1(_08748_),
    .Y(_09063_));
 sky130_fd_sc_hd__o2bb2a_1 _21825_ (.A1_N(_08795_),
    .A2_N(_09059_),
    .B1(_09061_),
    .B2(_09063_),
    .X(_09064_));
 sky130_fd_sc_hd__nor2_1 _21826_ (.A(_08510_),
    .B(_09064_),
    .Y(_09065_));
 sky130_fd_sc_hd__mux4_1 _21827_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][23] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][23] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][23] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][23] ),
    .S0(_08578_),
    .S1(_08684_),
    .X(_09066_));
 sky130_fd_sc_hd__mux4_1 _21828_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][23] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][23] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][23] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][23] ),
    .S0(_08560_),
    .S1(_08561_),
    .X(_09067_));
 sky130_fd_sc_hd__or2_1 _21829_ (.A(_08835_),
    .B(_09067_),
    .X(_09068_));
 sky130_fd_sc_hd__o211a_1 _21830_ (.A1(_08682_),
    .A2(_09066_),
    .B1(_09068_),
    .C1(_08558_),
    .X(_09069_));
 sky130_fd_sc_hd__mux4_1 _21831_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][23] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][23] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][23] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][23] ),
    .S0(_08839_),
    .S1(_08840_),
    .X(_09070_));
 sky130_fd_sc_hd__mux4_1 _21832_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][23] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][23] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][23] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][23] ),
    .S0(_08550_),
    .S1(_08554_),
    .X(_09071_));
 sky130_fd_sc_hd__or2_1 _21833_ (.A(_08842_),
    .B(_09071_),
    .X(_09072_));
 sky130_fd_sc_hd__o211a_1 _21834_ (.A1(_08547_),
    .A2(_09070_),
    .B1(_09072_),
    .C1(_08576_),
    .X(_09073_));
 sky130_fd_sc_hd__o31a_1 _21835_ (.A1(_09065_),
    .A2(_09069_),
    .A3(_09073_),
    .B1(_08624_),
    .X(_01051_));
 sky130_fd_sc_hd__mux4_1 _21836_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][24] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][24] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][24] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][24] ),
    .S0(_08517_),
    .S1(_08519_),
    .X(_09074_));
 sky130_fd_sc_hd__nor2_1 _21837_ (.A(_08515_),
    .B(_09074_),
    .Y(_09075_));
 sky130_fd_sc_hd__mux4_1 _21838_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][24] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][24] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][24] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][24] ),
    .S0(_08525_),
    .S1(_08528_),
    .X(_09076_));
 sky130_fd_sc_hd__nor2_1 _21839_ (.A(_08523_),
    .B(_09076_),
    .Y(_09077_));
 sky130_fd_sc_hd__mux4_1 _21840_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][24] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][24] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][24] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][24] ),
    .S0(_08534_),
    .S1(_08537_),
    .X(_09078_));
 sky130_fd_sc_hd__nor2_1 _21841_ (.A(_08532_),
    .B(_09078_),
    .Y(_09079_));
 sky130_fd_sc_hd__mux4_1 _21842_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][24] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][24] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][24] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][24] ),
    .S0(_08525_),
    .S1(_08528_),
    .X(_09080_));
 sky130_fd_sc_hd__o21ai_1 _21843_ (.A1(_08542_),
    .A2(_09080_),
    .B1(_08513_),
    .Y(_09081_));
 sky130_fd_sc_hd__o32a_1 _21844_ (.A1(_08513_),
    .A2(_09075_),
    .A3(_09077_),
    .B1(_09079_),
    .B2(_09081_),
    .X(_09082_));
 sky130_fd_sc_hd__nor2_1 _21845_ (.A(_08510_),
    .B(_09082_),
    .Y(_09083_));
 sky130_fd_sc_hd__mux4_2 _21846_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][24] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][24] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][24] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][24] ),
    .S0(_08578_),
    .S1(_08684_),
    .X(_09084_));
 sky130_fd_sc_hd__mux4_1 _21847_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][24] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][24] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][24] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][24] ),
    .S0(_08635_),
    .S1(_08561_),
    .X(_09085_));
 sky130_fd_sc_hd__or2_1 _21848_ (.A(_08835_),
    .B(_09085_),
    .X(_09086_));
 sky130_fd_sc_hd__o211a_1 _21849_ (.A1(_08682_),
    .A2(_09084_),
    .B1(_09086_),
    .C1(_08558_),
    .X(_09087_));
 sky130_fd_sc_hd__mux4_1 _21850_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][24] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][24] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][24] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][24] ),
    .S0(_08839_),
    .S1(_08840_),
    .X(_09088_));
 sky130_fd_sc_hd__mux4_1 _21851_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][24] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][24] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][24] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][24] ),
    .S0(_08550_),
    .S1(_08554_),
    .X(_09089_));
 sky130_fd_sc_hd__or2_1 _21852_ (.A(_08842_),
    .B(_09089_),
    .X(_09090_));
 sky130_fd_sc_hd__o211a_1 _21853_ (.A1(_08547_),
    .A2(_09088_),
    .B1(_09090_),
    .C1(_08576_),
    .X(_09091_));
 sky130_fd_sc_hd__o31a_1 _21854_ (.A1(_09083_),
    .A2(_09087_),
    .A3(_09091_),
    .B1(_08624_),
    .X(_01052_));
 sky130_fd_sc_hd__mux4_1 _21855_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][25] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][25] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][25] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][25] ),
    .S0(_08631_),
    .S1(_08632_),
    .X(_09092_));
 sky130_fd_sc_hd__mux4_1 _21856_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][25] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][25] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][25] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][25] ),
    .S0(_08778_),
    .S1(_08825_),
    .X(_09093_));
 sky130_fd_sc_hd__mux2_1 _21857_ (.A0(_09092_),
    .A1(_09093_),
    .S(_08743_),
    .X(_09094_));
 sky130_fd_sc_hd__mux4_1 _21858_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][25] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][25] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][25] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][25] ),
    .S0(_08525_),
    .S1(_08528_),
    .X(_09095_));
 sky130_fd_sc_hd__nor2_1 _21859_ (.A(_08515_),
    .B(_09095_),
    .Y(_09096_));
 sky130_fd_sc_hd__mux4_1 _21860_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][25] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][25] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][25] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][25] ),
    .S0(_08568_),
    .S1(_08683_),
    .X(_09097_));
 sky130_fd_sc_hd__o21ai_1 _21861_ (.A1(_08523_),
    .A2(_09097_),
    .B1(_08748_),
    .Y(_09098_));
 sky130_fd_sc_hd__o2bb2a_1 _21862_ (.A1_N(_08795_),
    .A2_N(_09094_),
    .B1(_09096_),
    .B2(_09098_),
    .X(_09099_));
 sky130_fd_sc_hd__nor2_1 _21863_ (.A(_08510_),
    .B(_09099_),
    .Y(_09100_));
 sky130_fd_sc_hd__mux4_1 _21864_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][25] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][25] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][25] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][25] ),
    .S0(_08578_),
    .S1(_08684_),
    .X(_09101_));
 sky130_fd_sc_hd__mux4_1 _21865_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][25] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][25] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][25] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][25] ),
    .S0(_08635_),
    .S1(_08637_),
    .X(_09102_));
 sky130_fd_sc_hd__or2_1 _21866_ (.A(_08835_),
    .B(_09102_),
    .X(_09103_));
 sky130_fd_sc_hd__o211a_1 _21867_ (.A1(_08682_),
    .A2(_09101_),
    .B1(_09103_),
    .C1(_08558_),
    .X(_09104_));
 sky130_fd_sc_hd__mux4_1 _21868_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][25] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][25] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][25] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][25] ),
    .S0(_08839_),
    .S1(_08840_),
    .X(_09105_));
 sky130_fd_sc_hd__mux4_1 _21869_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][25] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][25] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][25] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][25] ),
    .S0(_08550_),
    .S1(_08554_),
    .X(_09106_));
 sky130_fd_sc_hd__or2_1 _21870_ (.A(_08842_),
    .B(_09106_),
    .X(_09107_));
 sky130_fd_sc_hd__o211a_1 _21871_ (.A1(_08547_),
    .A2(_09105_),
    .B1(_09107_),
    .C1(_08576_),
    .X(_09108_));
 sky130_fd_sc_hd__o31a_1 _21872_ (.A1(_09100_),
    .A2(_09104_),
    .A3(_09108_),
    .B1(_08624_),
    .X(_01053_));
 sky130_fd_sc_hd__mux4_1 _21873_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][26] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][26] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][26] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][26] ),
    .S0(_08631_),
    .S1(_08632_),
    .X(_09109_));
 sky130_fd_sc_hd__mux4_1 _21874_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][26] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][26] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][26] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][26] ),
    .S0(_08778_),
    .S1(_08825_),
    .X(_09110_));
 sky130_fd_sc_hd__mux2_1 _21875_ (.A0(_09109_),
    .A1(_09110_),
    .S(_08673_),
    .X(_09111_));
 sky130_fd_sc_hd__mux4_1 _21876_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][26] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][26] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][26] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][26] ),
    .S0(_08629_),
    .S1(_08683_),
    .X(_09112_));
 sky130_fd_sc_hd__nor2_1 _21877_ (.A(_08725_),
    .B(_09112_),
    .Y(_09113_));
 sky130_fd_sc_hd__mux4_1 _21878_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][26] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][26] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][26] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][26] ),
    .S0(_08536_),
    .S1(_08693_),
    .X(_09114_));
 sky130_fd_sc_hd__o21ai_1 _21879_ (.A1(_08686_),
    .A2(_09114_),
    .B1(_08806_),
    .Y(_09115_));
 sky130_fd_sc_hd__o2bb2a_1 _21880_ (.A1_N(_08795_),
    .A2_N(_09111_),
    .B1(_09113_),
    .B2(_09115_),
    .X(_09116_));
 sky130_fd_sc_hd__nor2_1 _21881_ (.A(_08510_),
    .B(_09116_),
    .Y(_09117_));
 sky130_fd_sc_hd__mux4_1 _21882_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][26] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][26] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][26] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][26] ),
    .S0(_08578_),
    .S1(_08684_),
    .X(_09118_));
 sky130_fd_sc_hd__mux4_1 _21883_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][26] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][26] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][26] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][26] ),
    .S0(_08635_),
    .S1(_08637_),
    .X(_09119_));
 sky130_fd_sc_hd__or2_1 _21884_ (.A(_08835_),
    .B(_09119_),
    .X(_09120_));
 sky130_fd_sc_hd__o211a_1 _21885_ (.A1(_08682_),
    .A2(_09118_),
    .B1(_09120_),
    .C1(_08558_),
    .X(_09121_));
 sky130_fd_sc_hd__mux4_1 _21886_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][26] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][26] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][26] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][26] ),
    .S0(_08839_),
    .S1(_08840_),
    .X(_09122_));
 sky130_fd_sc_hd__mux4_1 _21887_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][26] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][26] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][26] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][26] ),
    .S0(_08550_),
    .S1(_08554_),
    .X(_09123_));
 sky130_fd_sc_hd__or2_1 _21888_ (.A(_08842_),
    .B(_09123_),
    .X(_09124_));
 sky130_fd_sc_hd__o211a_1 _21889_ (.A1(_08547_),
    .A2(_09122_),
    .B1(_09124_),
    .C1(_08575_),
    .X(_09125_));
 sky130_fd_sc_hd__o31a_1 _21890_ (.A1(_09117_),
    .A2(_09121_),
    .A3(_09125_),
    .B1(_08624_),
    .X(_01054_));
 sky130_fd_sc_hd__mux4_1 _21891_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][27] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][27] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][27] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][27] ),
    .S0(_08799_),
    .S1(_08800_),
    .X(_09126_));
 sky130_fd_sc_hd__or2_1 _21892_ (.A(_08514_),
    .B(_09126_),
    .X(_09127_));
 sky130_fd_sc_hd__mux4_1 _21893_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][27] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][27] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][27] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][27] ),
    .S0(_08516_),
    .S1(_08518_),
    .X(_09128_));
 sky130_fd_sc_hd__or2_1 _21894_ (.A(_08522_),
    .B(_09128_),
    .X(_09129_));
 sky130_fd_sc_hd__mux4_1 _21895_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][27] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][27] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][27] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][27] ),
    .S0(_08552_),
    .S1(_08687_),
    .X(_09130_));
 sky130_fd_sc_hd__mux4_1 _21896_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][27] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][27] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][27] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][27] ),
    .S0(\rvcpu.dp.plfd.InstrD[15] ),
    .S1(_08526_),
    .X(_09131_));
 sky130_fd_sc_hd__or2_1 _21897_ (.A(_08742_),
    .B(_09131_),
    .X(_09132_));
 sky130_fd_sc_hd__o211a_1 _21898_ (.A1(_08798_),
    .A2(_09130_),
    .B1(_09132_),
    .C1(_08512_),
    .X(_09133_));
 sky130_fd_sc_hd__a311o_1 _21899_ (.A1(_08626_),
    .A2(_09127_),
    .A3(_09129_),
    .B1(_09133_),
    .C1(_08509_),
    .X(_09134_));
 sky130_fd_sc_hd__mux4_1 _21900_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][27] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][27] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][27] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][27] ),
    .S0(_08810_),
    .S1(_08811_),
    .X(_09135_));
 sky130_fd_sc_hd__mux4_1 _21901_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][27] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][27] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][27] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][27] ),
    .S0(_08628_),
    .S1(_08856_),
    .X(_09136_));
 sky130_fd_sc_hd__a21o_1 _21902_ (.A1(_08813_),
    .A2(_09136_),
    .B1(_08579_),
    .X(_09137_));
 sky130_fd_sc_hd__a21o_1 _21903_ (.A1(_08692_),
    .A2(_09135_),
    .B1(_09137_),
    .X(_09138_));
 sky130_fd_sc_hd__mux4_1 _21904_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][27] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][27] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][27] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][27] ),
    .S0(_08534_),
    .S1(_08818_),
    .X(_09139_));
 sky130_fd_sc_hd__mux4_1 _21905_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][27] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][27] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][27] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][27] ),
    .S0(_08549_),
    .S1(_08553_),
    .X(_09140_));
 sky130_fd_sc_hd__and2_1 _21906_ (.A(_08541_),
    .B(_09140_),
    .X(_09141_));
 sky130_fd_sc_hd__a211o_1 _21907_ (.A1(_08817_),
    .A2(_09139_),
    .B1(_09141_),
    .C1(_08700_),
    .X(_09142_));
 sky130_fd_sc_hd__and4_1 _21908_ (.A(_08623_),
    .B(_09134_),
    .C(_09138_),
    .D(_09142_),
    .X(_09143_));
 sky130_fd_sc_hd__clkbuf_1 _21909_ (.A(_09143_),
    .X(_01055_));
 sky130_fd_sc_hd__mux4_1 _21910_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][28] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][28] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][28] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][28] ),
    .S0(_08516_),
    .S1(_08518_),
    .X(_09144_));
 sky130_fd_sc_hd__mux4_1 _21911_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][28] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][28] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][28] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][28] ),
    .S0(_08516_),
    .S1(_08518_),
    .X(_09145_));
 sky130_fd_sc_hd__mux2_1 _21912_ (.A0(_09144_),
    .A1(_09145_),
    .S(_08540_),
    .X(_09146_));
 sky130_fd_sc_hd__mux4_1 _21913_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][28] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][28] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][28] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][28] ),
    .S0(_08549_),
    .S1(_08553_),
    .X(_09147_));
 sky130_fd_sc_hd__or2_1 _21914_ (.A(_08673_),
    .B(_09147_),
    .X(_09148_));
 sky130_fd_sc_hd__mux4_2 _21915_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][28] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][28] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][28] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][28] ),
    .S0(_08533_),
    .S1(_08536_),
    .X(_09149_));
 sky130_fd_sc_hd__o21a_1 _21916_ (.A1(_08531_),
    .A2(_09149_),
    .B1(_08806_),
    .X(_09150_));
 sky130_fd_sc_hd__a221o_1 _21917_ (.A1(_08626_),
    .A2(_09146_),
    .B1(_09148_),
    .B2(_09150_),
    .C1(_08808_),
    .X(_09151_));
 sky130_fd_sc_hd__mux4_1 _21918_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][28] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][28] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][28] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][28] ),
    .S0(_08810_),
    .S1(_08811_),
    .X(_09152_));
 sky130_fd_sc_hd__mux4_1 _21919_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][28] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][28] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][28] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][28] ),
    .S0(_08628_),
    .S1(_08856_),
    .X(_09153_));
 sky130_fd_sc_hd__a21o_1 _21920_ (.A1(_08813_),
    .A2(_09153_),
    .B1(_08579_),
    .X(_09154_));
 sky130_fd_sc_hd__a21o_1 _21921_ (.A1(_08692_),
    .A2(_09152_),
    .B1(_09154_),
    .X(_09155_));
 sky130_fd_sc_hd__mux4_1 _21922_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][28] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][28] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][28] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][28] ),
    .S0(_08534_),
    .S1(_08818_),
    .X(_09156_));
 sky130_fd_sc_hd__mux4_1 _21923_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][28] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][28] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][28] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][28] ),
    .S0(_08549_),
    .S1(_08553_),
    .X(_09157_));
 sky130_fd_sc_hd__and2_1 _21924_ (.A(_08541_),
    .B(_09157_),
    .X(_09158_));
 sky130_fd_sc_hd__a211o_1 _21925_ (.A1(_08817_),
    .A2(_09156_),
    .B1(_09158_),
    .C1(_08699_),
    .X(_09159_));
 sky130_fd_sc_hd__and4_1 _21926_ (.A(_08623_),
    .B(_09151_),
    .C(_09155_),
    .D(_09159_),
    .X(_09160_));
 sky130_fd_sc_hd__clkbuf_1 _21927_ (.A(_09160_),
    .X(_01056_));
 sky130_fd_sc_hd__mux4_1 _21928_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][29] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][29] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][29] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][29] ),
    .S0(_08631_),
    .S1(_08632_),
    .X(_09161_));
 sky130_fd_sc_hd__mux4_1 _21929_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][29] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][29] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][29] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][29] ),
    .S0(_08778_),
    .S1(_08825_),
    .X(_09162_));
 sky130_fd_sc_hd__mux2_1 _21930_ (.A0(_09161_),
    .A1(_09162_),
    .S(_08673_),
    .X(_09163_));
 sky130_fd_sc_hd__mux4_1 _21931_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][29] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][29] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][29] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][29] ),
    .S0(_08629_),
    .S1(_08683_),
    .X(_09164_));
 sky130_fd_sc_hd__nor2_1 _21932_ (.A(_08725_),
    .B(_09164_),
    .Y(_09165_));
 sky130_fd_sc_hd__mux4_1 _21933_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][29] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][29] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][29] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][29] ),
    .S0(_08536_),
    .S1(_08693_),
    .X(_09166_));
 sky130_fd_sc_hd__o21ai_1 _21934_ (.A1(_08686_),
    .A2(_09166_),
    .B1(_08806_),
    .Y(_09167_));
 sky130_fd_sc_hd__o2bb2a_1 _21935_ (.A1_N(_08795_),
    .A2_N(_09163_),
    .B1(_09165_),
    .B2(_09167_),
    .X(_09168_));
 sky130_fd_sc_hd__nor2_1 _21936_ (.A(_08510_),
    .B(_09168_),
    .Y(_09169_));
 sky130_fd_sc_hd__mux4_1 _21937_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][29] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][29] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][29] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][29] ),
    .S0(_08578_),
    .S1(_08684_),
    .X(_09170_));
 sky130_fd_sc_hd__mux4_1 _21938_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][29] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][29] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][29] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][29] ),
    .S0(_08525_),
    .S1(_08528_),
    .X(_09171_));
 sky130_fd_sc_hd__or2_1 _21939_ (.A(_08835_),
    .B(_09171_),
    .X(_09172_));
 sky130_fd_sc_hd__o211a_1 _21940_ (.A1(_08682_),
    .A2(_09170_),
    .B1(_09172_),
    .C1(_08575_),
    .X(_09173_));
 sky130_fd_sc_hd__mux4_1 _21941_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][29] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][29] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][29] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][29] ),
    .S0(_08839_),
    .S1(_08840_),
    .X(_09174_));
 sky130_fd_sc_hd__mux4_1 _21942_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][29] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][29] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][29] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][29] ),
    .S0(_08649_),
    .S1(_08561_),
    .X(_09175_));
 sky130_fd_sc_hd__or2_1 _21943_ (.A(_08842_),
    .B(_09175_),
    .X(_09176_));
 sky130_fd_sc_hd__o211a_1 _21944_ (.A1(_08547_),
    .A2(_09174_),
    .B1(_09176_),
    .C1(_08652_),
    .X(_09177_));
 sky130_fd_sc_hd__o31a_1 _21945_ (.A1(_09169_),
    .A2(_09173_),
    .A3(_09177_),
    .B1(_08624_),
    .X(_01057_));
 sky130_fd_sc_hd__mux4_1 _21946_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][30] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][30] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][30] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][30] ),
    .S0(_08516_),
    .S1(_08518_),
    .X(_09178_));
 sky130_fd_sc_hd__mux4_1 _21947_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][30] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][30] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][30] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][30] ),
    .S0(_08535_),
    .S1(_08533_),
    .X(_09179_));
 sky130_fd_sc_hd__mux2_1 _21948_ (.A0(_09178_),
    .A1(_09179_),
    .S(_08540_),
    .X(_09180_));
 sky130_fd_sc_hd__mux4_2 _21949_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][30] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][30] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][30] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][30] ),
    .S0(_08549_),
    .S1(_08527_),
    .X(_09181_));
 sky130_fd_sc_hd__or2_1 _21950_ (.A(_08673_),
    .B(_09181_),
    .X(_09182_));
 sky130_fd_sc_hd__mux4_2 _21951_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][30] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][30] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][30] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][30] ),
    .S0(_08533_),
    .S1(_08636_),
    .X(_09183_));
 sky130_fd_sc_hd__o21a_1 _21952_ (.A1(_08531_),
    .A2(_09183_),
    .B1(_08806_),
    .X(_09184_));
 sky130_fd_sc_hd__a221o_1 _21953_ (.A1(_08626_),
    .A2(_09180_),
    .B1(_09182_),
    .B2(_09184_),
    .C1(_08808_),
    .X(_09185_));
 sky130_fd_sc_hd__mux4_1 _21954_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][30] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][30] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][30] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][30] ),
    .S0(_08566_),
    .S1(_08569_),
    .X(_09186_));
 sky130_fd_sc_hd__mux4_1 _21955_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][30] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][30] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][30] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][30] ),
    .S0(_08628_),
    .S1(_08856_),
    .X(_09187_));
 sky130_fd_sc_hd__a21o_1 _21956_ (.A1(_08695_),
    .A2(_09187_),
    .B1(_08579_),
    .X(_09188_));
 sky130_fd_sc_hd__a21o_1 _21957_ (.A1(_08692_),
    .A2(_09186_),
    .B1(_09188_),
    .X(_09189_));
 sky130_fd_sc_hd__mux4_1 _21958_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][30] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][30] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][30] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][30] ),
    .S0(_08534_),
    .S1(_08537_),
    .X(_09190_));
 sky130_fd_sc_hd__mux4_1 _21959_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][30] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][30] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][30] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][30] ),
    .S0(_08549_),
    .S1(_08553_),
    .X(_09191_));
 sky130_fd_sc_hd__and2_1 _21960_ (.A(_08541_),
    .B(_09191_),
    .X(_09192_));
 sky130_fd_sc_hd__a211o_1 _21961_ (.A1(_08532_),
    .A2(_09190_),
    .B1(_09192_),
    .C1(_08699_),
    .X(_09193_));
 sky130_fd_sc_hd__and4_1 _21962_ (.A(_08623_),
    .B(_09185_),
    .C(_09189_),
    .D(_09193_),
    .X(_09194_));
 sky130_fd_sc_hd__clkbuf_1 _21963_ (.A(_09194_),
    .X(_01058_));
 sky130_fd_sc_hd__mux4_2 _21964_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][31] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][31] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][31] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][31] ),
    .S0(_08548_),
    .S1(_08552_),
    .X(_09195_));
 sky130_fd_sc_hd__or2_1 _21965_ (.A(_08742_),
    .B(_09195_),
    .X(_09196_));
 sky130_fd_sc_hd__mux4_2 _21966_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][31] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][31] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][31] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][31] ),
    .S0(\rvcpu.dp.plfd.InstrD[16] ),
    .S1(_08516_),
    .X(_09197_));
 sky130_fd_sc_hd__o21a_1 _21967_ (.A1(_08522_),
    .A2(_09197_),
    .B1(_08512_),
    .X(_09198_));
 sky130_fd_sc_hd__mux4_1 _21968_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][31] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][31] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][31] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][31] ),
    .S0(_08548_),
    .S1(_08552_),
    .X(_09199_));
 sky130_fd_sc_hd__mux4_1 _21969_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][31] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][31] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][31] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][31] ),
    .S0(_08548_),
    .S1(_08552_),
    .X(_09200_));
 sky130_fd_sc_hd__mux2_1 _21970_ (.A0(_09199_),
    .A1(_09200_),
    .S(\rvcpu.dp.plfd.InstrD[17] ),
    .X(_09201_));
 sky130_fd_sc_hd__a22o_1 _21971_ (.A1(_09196_),
    .A2(_09198_),
    .B1(_09201_),
    .B2(_08557_),
    .X(_09202_));
 sky130_fd_sc_hd__mux4_1 _21972_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][31] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][31] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][31] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][31] ),
    .S0(_08696_),
    .S1(_08825_),
    .X(_09203_));
 sky130_fd_sc_hd__mux4_1 _21973_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][31] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][31] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][31] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][31] ),
    .S0(_08535_),
    .S1(_08552_),
    .X(_09204_));
 sky130_fd_sc_hd__or2_1 _21974_ (.A(_08540_),
    .B(_09204_),
    .X(_09205_));
 sky130_fd_sc_hd__o211a_1 _21975_ (.A1(_08523_),
    .A2(_09203_),
    .B1(_09205_),
    .C1(_08575_),
    .X(_09206_));
 sky130_fd_sc_hd__mux4_1 _21976_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][31] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][31] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][31] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][31] ),
    .S0(_08628_),
    .S1(_08629_),
    .X(_09207_));
 sky130_fd_sc_hd__mux4_1 _21977_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][31] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][31] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][31] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][31] ),
    .S0(\rvcpu.dp.plfd.InstrD[16] ),
    .S1(_08524_),
    .X(_09208_));
 sky130_fd_sc_hd__or2_1 _21978_ (.A(_08540_),
    .B(_09208_),
    .X(_09209_));
 sky130_fd_sc_hd__o211a_1 _21979_ (.A1(_08523_),
    .A2(_09207_),
    .B1(_09209_),
    .C1(_08558_),
    .X(_09210_));
 sky130_fd_sc_hd__a211o_1 _21980_ (.A1(\rvcpu.dp.plfd.InstrD[19] ),
    .A2(_09202_),
    .B1(_09206_),
    .C1(_09210_),
    .X(_09211_));
 sky130_fd_sc_hd__and2_1 _21981_ (.A(_08624_),
    .B(_09211_),
    .X(_09212_));
 sky130_fd_sc_hd__clkbuf_1 _21982_ (.A(_09212_),
    .X(_01059_));
 sky130_fd_sc_hd__nand2_2 _21983_ (.A(_06585_),
    .B(\rvcpu.dp.plem.MemWriteM ),
    .Y(_09213_));
 sky130_fd_sc_hd__or2_1 _21984_ (.A(_06582_),
    .B(_09213_),
    .X(_09214_));
 sky130_fd_sc_hd__buf_4 _21985_ (.A(_09214_),
    .X(_09215_));
 sky130_fd_sc_hd__inv_2 _21986_ (.A(_08488_),
    .Y(_09216_));
 sky130_fd_sc_hd__a21o_1 _21987_ (.A1(_05391_),
    .A2(net117),
    .B1(_09216_),
    .X(_09217_));
 sky130_fd_sc_hd__and3_1 _21988_ (.A(\rvcpu.dp.plem.MemWriteM ),
    .B(_06911_),
    .C(_09217_),
    .X(_09218_));
 sky130_fd_sc_hd__clkbuf_8 _21989_ (.A(_09218_),
    .X(_09219_));
 sky130_fd_sc_hd__nor2_8 _21990_ (.A(_06582_),
    .B(_09213_),
    .Y(_09220_));
 sky130_fd_sc_hd__clkbuf_4 _21991_ (.A(_09220_),
    .X(_09221_));
 sky130_fd_sc_hd__and2_1 _21992_ (.A(\rvcpu.dp.plem.WriteDataM[16] ),
    .B(_09221_),
    .X(_09222_));
 sky130_fd_sc_hd__a31o_4 _21993_ (.A1(\rvcpu.dp.plem.WriteDataM[0] ),
    .A2(_09215_),
    .A3(_09219_),
    .B1(_09222_),
    .X(_09223_));
 sky130_fd_sc_hd__clkbuf_2 _21994_ (.A(_09223_),
    .X(_09224_));
 sky130_fd_sc_hd__clkbuf_16 _21995_ (.A(_07159_),
    .X(_09225_));
 sky130_fd_sc_hd__buf_8 _21996_ (.A(_09225_),
    .X(_09226_));
 sky130_fd_sc_hd__nand2_8 _21997_ (.A(_06603_),
    .B(_08355_),
    .Y(_09227_));
 sky130_fd_sc_hd__nor2_8 _21998_ (.A(_09220_),
    .B(_09219_),
    .Y(_09228_));
 sky130_fd_sc_hd__nor2_8 _21999_ (.A(_09227_),
    .B(net104),
    .Y(_09229_));
 sky130_fd_sc_hd__buf_8 _22000_ (.A(_06591_),
    .X(_09230_));
 sky130_fd_sc_hd__buf_8 _22001_ (.A(_09230_),
    .X(_09231_));
 sky130_fd_sc_hd__a21oi_4 _22002_ (.A1(_09226_),
    .A2(_09229_),
    .B1(_09231_),
    .Y(_09232_));
 sky130_fd_sc_hd__mux2_1 _22003_ (.A0(_09224_),
    .A1(\datamem.data_ram[62][16] ),
    .S(_09232_),
    .X(_09233_));
 sky130_fd_sc_hd__clkbuf_1 _22004_ (.A(_09233_),
    .X(_01060_));
 sky130_fd_sc_hd__and2_1 _22005_ (.A(\rvcpu.dp.plem.WriteDataM[17] ),
    .B(_09221_),
    .X(_09234_));
 sky130_fd_sc_hd__a31o_4 _22006_ (.A1(\rvcpu.dp.plem.WriteDataM[1] ),
    .A2(_09215_),
    .A3(_09219_),
    .B1(_09234_),
    .X(_09235_));
 sky130_fd_sc_hd__clkbuf_2 _22007_ (.A(_09235_),
    .X(_09236_));
 sky130_fd_sc_hd__mux2_1 _22008_ (.A0(_09236_),
    .A1(\datamem.data_ram[62][17] ),
    .S(_09232_),
    .X(_09237_));
 sky130_fd_sc_hd__clkbuf_1 _22009_ (.A(_09237_),
    .X(_01061_));
 sky130_fd_sc_hd__and2_1 _22010_ (.A(\rvcpu.dp.plem.WriteDataM[18] ),
    .B(_09221_),
    .X(_09238_));
 sky130_fd_sc_hd__a31o_4 _22011_ (.A1(\rvcpu.dp.plem.WriteDataM[2] ),
    .A2(_09215_),
    .A3(_09219_),
    .B1(_09238_),
    .X(_09239_));
 sky130_fd_sc_hd__clkbuf_2 _22012_ (.A(_09239_),
    .X(_09240_));
 sky130_fd_sc_hd__mux2_1 _22013_ (.A0(_09240_),
    .A1(\datamem.data_ram[62][18] ),
    .S(_09232_),
    .X(_09241_));
 sky130_fd_sc_hd__clkbuf_1 _22014_ (.A(_09241_),
    .X(_01062_));
 sky130_fd_sc_hd__and2_1 _22015_ (.A(\rvcpu.dp.plem.WriteDataM[19] ),
    .B(_09221_),
    .X(_09242_));
 sky130_fd_sc_hd__a31o_4 _22016_ (.A1(\rvcpu.dp.plem.WriteDataM[3] ),
    .A2(_09215_),
    .A3(_09219_),
    .B1(_09242_),
    .X(_09243_));
 sky130_fd_sc_hd__clkbuf_2 _22017_ (.A(_09243_),
    .X(_09244_));
 sky130_fd_sc_hd__mux2_1 _22018_ (.A0(_09244_),
    .A1(\datamem.data_ram[62][19] ),
    .S(_09232_),
    .X(_09245_));
 sky130_fd_sc_hd__clkbuf_1 _22019_ (.A(_09245_),
    .X(_01063_));
 sky130_fd_sc_hd__and2_1 _22020_ (.A(\rvcpu.dp.plem.WriteDataM[20] ),
    .B(_09221_),
    .X(_09246_));
 sky130_fd_sc_hd__a31o_4 _22021_ (.A1(\rvcpu.dp.plem.WriteDataM[4] ),
    .A2(_09215_),
    .A3(_09219_),
    .B1(_09246_),
    .X(_09247_));
 sky130_fd_sc_hd__clkbuf_2 _22022_ (.A(_09247_),
    .X(_09248_));
 sky130_fd_sc_hd__mux2_1 _22023_ (.A0(_09248_),
    .A1(\datamem.data_ram[62][20] ),
    .S(_09232_),
    .X(_09249_));
 sky130_fd_sc_hd__clkbuf_1 _22024_ (.A(_09249_),
    .X(_01064_));
 sky130_fd_sc_hd__and2_1 _22025_ (.A(\rvcpu.dp.plem.WriteDataM[21] ),
    .B(_09220_),
    .X(_09250_));
 sky130_fd_sc_hd__a31o_4 _22026_ (.A1(\rvcpu.dp.plem.WriteDataM[5] ),
    .A2(_09215_),
    .A3(_09219_),
    .B1(_09250_),
    .X(_09251_));
 sky130_fd_sc_hd__clkbuf_2 _22027_ (.A(_09251_),
    .X(_09252_));
 sky130_fd_sc_hd__mux2_1 _22028_ (.A0(_09252_),
    .A1(\datamem.data_ram[62][21] ),
    .S(_09232_),
    .X(_09253_));
 sky130_fd_sc_hd__clkbuf_1 _22029_ (.A(_09253_),
    .X(_01065_));
 sky130_fd_sc_hd__and2_1 _22030_ (.A(\rvcpu.dp.plem.WriteDataM[22] ),
    .B(_09220_),
    .X(_09254_));
 sky130_fd_sc_hd__a31o_4 _22031_ (.A1(\rvcpu.dp.plem.WriteDataM[6] ),
    .A2(_09215_),
    .A3(_09219_),
    .B1(_09254_),
    .X(_09255_));
 sky130_fd_sc_hd__clkbuf_2 _22032_ (.A(_09255_),
    .X(_09256_));
 sky130_fd_sc_hd__mux2_1 _22033_ (.A0(_09256_),
    .A1(\datamem.data_ram[62][22] ),
    .S(_09232_),
    .X(_09257_));
 sky130_fd_sc_hd__clkbuf_1 _22034_ (.A(_09257_),
    .X(_01066_));
 sky130_fd_sc_hd__and2_1 _22035_ (.A(\rvcpu.dp.plem.WriteDataM[23] ),
    .B(_09220_),
    .X(_09258_));
 sky130_fd_sc_hd__a31o_4 _22036_ (.A1(\rvcpu.dp.plem.WriteDataM[7] ),
    .A2(_09215_),
    .A3(_09219_),
    .B1(_09258_),
    .X(_09259_));
 sky130_fd_sc_hd__clkbuf_2 _22037_ (.A(_09259_),
    .X(_09260_));
 sky130_fd_sc_hd__mux2_1 _22038_ (.A0(_09260_),
    .A1(\datamem.data_ram[62][23] ),
    .S(_09232_),
    .X(_09261_));
 sky130_fd_sc_hd__clkbuf_1 _22039_ (.A(_09261_),
    .X(_01067_));
 sky130_fd_sc_hd__nor2_2 _22040_ (.A(\rvcpu.dp.plem.ALUResultM[1] ),
    .B(_09213_),
    .Y(_09262_));
 sky130_fd_sc_hd__and3_1 _22041_ (.A(\rvcpu.dp.plem.ALUResultM[0] ),
    .B(net117),
    .C(_09262_),
    .X(_09263_));
 sky130_fd_sc_hd__buf_4 _22042_ (.A(_09263_),
    .X(_09264_));
 sky130_fd_sc_hd__a21o_4 _22043_ (.A1(_09216_),
    .A2(_09262_),
    .B1(_09220_),
    .X(_09265_));
 sky130_fd_sc_hd__a22o_4 _22044_ (.A1(\rvcpu.dp.plem.WriteDataM[0] ),
    .A2(_09264_),
    .B1(_09265_),
    .B2(\rvcpu.dp.plem.WriteDataM[8] ),
    .X(_09266_));
 sky130_fd_sc_hd__buf_2 _22045_ (.A(_09266_),
    .X(_09267_));
 sky130_fd_sc_hd__nor2_8 _22046_ (.A(_09264_),
    .B(_09265_),
    .Y(_09268_));
 sky130_fd_sc_hd__nor2_8 _22047_ (.A(_09227_),
    .B(net112),
    .Y(_09269_));
 sky130_fd_sc_hd__a21oi_4 _22048_ (.A1(_09226_),
    .A2(_09269_),
    .B1(_09231_),
    .Y(_09270_));
 sky130_fd_sc_hd__mux2_1 _22049_ (.A0(_09267_),
    .A1(\datamem.data_ram[62][8] ),
    .S(_09270_),
    .X(_09271_));
 sky130_fd_sc_hd__clkbuf_1 _22050_ (.A(_09271_),
    .X(_01068_));
 sky130_fd_sc_hd__a22o_4 _22051_ (.A1(\rvcpu.dp.plem.WriteDataM[1] ),
    .A2(_09264_),
    .B1(_09265_),
    .B2(\rvcpu.dp.plem.WriteDataM[9] ),
    .X(_09272_));
 sky130_fd_sc_hd__clkbuf_4 _22052_ (.A(_09272_),
    .X(_09273_));
 sky130_fd_sc_hd__mux2_1 _22053_ (.A0(_09273_),
    .A1(\datamem.data_ram[62][9] ),
    .S(_09270_),
    .X(_09274_));
 sky130_fd_sc_hd__clkbuf_1 _22054_ (.A(_09274_),
    .X(_01069_));
 sky130_fd_sc_hd__a22o_4 _22055_ (.A1(\rvcpu.dp.plem.WriteDataM[2] ),
    .A2(_09264_),
    .B1(_09265_),
    .B2(\rvcpu.dp.plem.WriteDataM[10] ),
    .X(_09275_));
 sky130_fd_sc_hd__buf_2 _22056_ (.A(_09275_),
    .X(_09276_));
 sky130_fd_sc_hd__mux2_1 _22057_ (.A0(_09276_),
    .A1(\datamem.data_ram[62][10] ),
    .S(_09270_),
    .X(_09277_));
 sky130_fd_sc_hd__clkbuf_1 _22058_ (.A(_09277_),
    .X(_01070_));
 sky130_fd_sc_hd__a22o_4 _22059_ (.A1(\rvcpu.dp.plem.WriteDataM[3] ),
    .A2(_09264_),
    .B1(_09265_),
    .B2(\rvcpu.dp.plem.WriteDataM[11] ),
    .X(_09278_));
 sky130_fd_sc_hd__buf_2 _22060_ (.A(_09278_),
    .X(_09279_));
 sky130_fd_sc_hd__mux2_1 _22061_ (.A0(_09279_),
    .A1(\datamem.data_ram[62][11] ),
    .S(_09270_),
    .X(_09280_));
 sky130_fd_sc_hd__clkbuf_1 _22062_ (.A(_09280_),
    .X(_01071_));
 sky130_fd_sc_hd__a22o_4 _22063_ (.A1(\rvcpu.dp.plem.WriteDataM[4] ),
    .A2(_09264_),
    .B1(_09265_),
    .B2(\rvcpu.dp.plem.WriteDataM[12] ),
    .X(_09281_));
 sky130_fd_sc_hd__buf_2 _22064_ (.A(_09281_),
    .X(_09282_));
 sky130_fd_sc_hd__mux2_1 _22065_ (.A0(_09282_),
    .A1(\datamem.data_ram[62][12] ),
    .S(_09270_),
    .X(_09283_));
 sky130_fd_sc_hd__clkbuf_1 _22066_ (.A(_09283_),
    .X(_01072_));
 sky130_fd_sc_hd__a22o_4 _22067_ (.A1(\rvcpu.dp.plem.WriteDataM[5] ),
    .A2(_09264_),
    .B1(_09265_),
    .B2(\rvcpu.dp.plem.WriteDataM[13] ),
    .X(_09284_));
 sky130_fd_sc_hd__buf_2 _22068_ (.A(_09284_),
    .X(_09285_));
 sky130_fd_sc_hd__mux2_1 _22069_ (.A0(_09285_),
    .A1(\datamem.data_ram[62][13] ),
    .S(_09270_),
    .X(_09286_));
 sky130_fd_sc_hd__clkbuf_1 _22070_ (.A(_09286_),
    .X(_01073_));
 sky130_fd_sc_hd__a22o_4 _22071_ (.A1(\rvcpu.dp.plem.WriteDataM[6] ),
    .A2(_09264_),
    .B1(_09265_),
    .B2(\rvcpu.dp.plem.WriteDataM[14] ),
    .X(_09287_));
 sky130_fd_sc_hd__buf_2 _22072_ (.A(_09287_),
    .X(_09288_));
 sky130_fd_sc_hd__mux2_1 _22073_ (.A0(_09288_),
    .A1(\datamem.data_ram[62][14] ),
    .S(_09270_),
    .X(_09289_));
 sky130_fd_sc_hd__clkbuf_1 _22074_ (.A(_09289_),
    .X(_01074_));
 sky130_fd_sc_hd__a22o_4 _22075_ (.A1(\rvcpu.dp.plem.WriteDataM[7] ),
    .A2(_09264_),
    .B1(_09265_),
    .B2(\rvcpu.dp.plem.WriteDataM[15] ),
    .X(_09290_));
 sky130_fd_sc_hd__clkbuf_2 _22076_ (.A(_09290_),
    .X(_09291_));
 sky130_fd_sc_hd__mux2_1 _22077_ (.A0(_09291_),
    .A1(\datamem.data_ram[62][15] ),
    .S(_09270_),
    .X(_09292_));
 sky130_fd_sc_hd__clkbuf_1 _22078_ (.A(_09292_),
    .X(_01075_));
 sky130_fd_sc_hd__and4_2 _22079_ (.A(\rvcpu.dp.plem.MemWriteM ),
    .B(\rvcpu.dp.plem.ALUResultM[0] ),
    .C(_06911_),
    .D(net117),
    .X(_09293_));
 sky130_fd_sc_hd__and3_1 _22080_ (.A(\rvcpu.dp.plem.MemWriteM ),
    .B(_06911_),
    .C(_09216_),
    .X(_09294_));
 sky130_fd_sc_hd__clkbuf_4 _22081_ (.A(_09294_),
    .X(_09295_));
 sky130_fd_sc_hd__a32o_1 _22082_ (.A1(\rvcpu.dp.plem.WriteDataM[0] ),
    .A2(_08488_),
    .A3(_09293_),
    .B1(_09295_),
    .B2(\rvcpu.dp.plem.WriteDataM[8] ),
    .X(_09296_));
 sky130_fd_sc_hd__mux2_8 _22083_ (.A0(\rvcpu.dp.plem.WriteDataM[24] ),
    .A1(_09296_),
    .S(_09215_),
    .X(_09297_));
 sky130_fd_sc_hd__clkbuf_2 _22084_ (.A(_09297_),
    .X(_09298_));
 sky130_fd_sc_hd__buf_6 _22085_ (.A(_07132_),
    .X(_09299_));
 sky130_fd_sc_hd__nor3_4 _22086_ (.A(_09220_),
    .B(_09293_),
    .C(_09295_),
    .Y(_09300_));
 sky130_fd_sc_hd__nor2_8 _22087_ (.A(_09227_),
    .B(net108),
    .Y(_09301_));
 sky130_fd_sc_hd__a21oi_4 _22088_ (.A1(_09299_),
    .A2(_09301_),
    .B1(_09231_),
    .Y(_09302_));
 sky130_fd_sc_hd__mux2_1 _22089_ (.A0(_09298_),
    .A1(\datamem.data_ram[61][24] ),
    .S(_09302_),
    .X(_09303_));
 sky130_fd_sc_hd__clkbuf_1 _22090_ (.A(_09303_),
    .X(_01076_));
 sky130_fd_sc_hd__a32o_1 _22091_ (.A1(\rvcpu.dp.plem.WriteDataM[1] ),
    .A2(_08488_),
    .A3(_09293_),
    .B1(_09295_),
    .B2(\rvcpu.dp.plem.WriteDataM[9] ),
    .X(_09304_));
 sky130_fd_sc_hd__mux2_8 _22092_ (.A0(\rvcpu.dp.plem.WriteDataM[25] ),
    .A1(_09304_),
    .S(_09215_),
    .X(_09305_));
 sky130_fd_sc_hd__buf_2 _22093_ (.A(_09305_),
    .X(_09306_));
 sky130_fd_sc_hd__mux2_1 _22094_ (.A0(_09306_),
    .A1(\datamem.data_ram[61][25] ),
    .S(_09302_),
    .X(_09307_));
 sky130_fd_sc_hd__clkbuf_1 _22095_ (.A(_09307_),
    .X(_01077_));
 sky130_fd_sc_hd__and3_1 _22096_ (.A(\rvcpu.dp.plem.WriteDataM[2] ),
    .B(_08488_),
    .C(_09293_),
    .X(_09308_));
 sky130_fd_sc_hd__a221o_4 _22097_ (.A1(\rvcpu.dp.plem.WriteDataM[26] ),
    .A2(_09221_),
    .B1(_09295_),
    .B2(\rvcpu.dp.plem.WriteDataM[10] ),
    .C1(_09308_),
    .X(_09309_));
 sky130_fd_sc_hd__clkbuf_2 _22098_ (.A(_09309_),
    .X(_09310_));
 sky130_fd_sc_hd__mux2_1 _22099_ (.A0(_09310_),
    .A1(\datamem.data_ram[61][26] ),
    .S(_09302_),
    .X(_09311_));
 sky130_fd_sc_hd__clkbuf_1 _22100_ (.A(_09311_),
    .X(_01078_));
 sky130_fd_sc_hd__and3_1 _22101_ (.A(\rvcpu.dp.plem.WriteDataM[3] ),
    .B(_08488_),
    .C(_09293_),
    .X(_09312_));
 sky130_fd_sc_hd__a221o_4 _22102_ (.A1(\rvcpu.dp.plem.WriteDataM[27] ),
    .A2(_09221_),
    .B1(_09295_),
    .B2(\rvcpu.dp.plem.WriteDataM[11] ),
    .C1(_09312_),
    .X(_09313_));
 sky130_fd_sc_hd__buf_2 _22103_ (.A(_09313_),
    .X(_09314_));
 sky130_fd_sc_hd__mux2_1 _22104_ (.A0(_09314_),
    .A1(\datamem.data_ram[61][27] ),
    .S(_09302_),
    .X(_09315_));
 sky130_fd_sc_hd__clkbuf_1 _22105_ (.A(_09315_),
    .X(_01079_));
 sky130_fd_sc_hd__a32o_1 _22106_ (.A1(\rvcpu.dp.plem.WriteDataM[4] ),
    .A2(_08488_),
    .A3(_09293_),
    .B1(_09295_),
    .B2(\rvcpu.dp.plem.WriteDataM[12] ),
    .X(_09316_));
 sky130_fd_sc_hd__mux2_8 _22107_ (.A0(\rvcpu.dp.plem.WriteDataM[28] ),
    .A1(_09316_),
    .S(_09214_),
    .X(_09317_));
 sky130_fd_sc_hd__clkbuf_2 _22108_ (.A(_09317_),
    .X(_09318_));
 sky130_fd_sc_hd__mux2_1 _22109_ (.A0(_09318_),
    .A1(\datamem.data_ram[61][28] ),
    .S(_09302_),
    .X(_09319_));
 sky130_fd_sc_hd__clkbuf_1 _22110_ (.A(_09319_),
    .X(_01080_));
 sky130_fd_sc_hd__and3_1 _22111_ (.A(\rvcpu.dp.plem.WriteDataM[5] ),
    .B(_08488_),
    .C(_09293_),
    .X(_09320_));
 sky130_fd_sc_hd__a221o_4 _22112_ (.A1(\rvcpu.dp.plem.WriteDataM[29] ),
    .A2(_09221_),
    .B1(_09295_),
    .B2(\rvcpu.dp.plem.WriteDataM[13] ),
    .C1(_09320_),
    .X(_09321_));
 sky130_fd_sc_hd__clkbuf_2 _22113_ (.A(_09321_),
    .X(_09322_));
 sky130_fd_sc_hd__mux2_1 _22114_ (.A0(_09322_),
    .A1(\datamem.data_ram[61][29] ),
    .S(_09302_),
    .X(_09323_));
 sky130_fd_sc_hd__clkbuf_1 _22115_ (.A(_09323_),
    .X(_01081_));
 sky130_fd_sc_hd__and3_1 _22116_ (.A(\rvcpu.dp.plem.WriteDataM[6] ),
    .B(_08488_),
    .C(_09293_),
    .X(_09324_));
 sky130_fd_sc_hd__a221o_4 _22117_ (.A1(\rvcpu.dp.plem.WriteDataM[30] ),
    .A2(_09221_),
    .B1(_09295_),
    .B2(\rvcpu.dp.plem.WriteDataM[14] ),
    .C1(_09324_),
    .X(_09325_));
 sky130_fd_sc_hd__clkbuf_2 _22118_ (.A(_09325_),
    .X(_09326_));
 sky130_fd_sc_hd__mux2_1 _22119_ (.A0(_09326_),
    .A1(\datamem.data_ram[61][30] ),
    .S(_09302_),
    .X(_09327_));
 sky130_fd_sc_hd__clkbuf_1 _22120_ (.A(_09327_),
    .X(_01082_));
 sky130_fd_sc_hd__and3_1 _22121_ (.A(\rvcpu.dp.plem.WriteDataM[7] ),
    .B(_08488_),
    .C(_09293_),
    .X(_09328_));
 sky130_fd_sc_hd__a221o_4 _22122_ (.A1(\rvcpu.dp.plem.WriteDataM[31] ),
    .A2(_09221_),
    .B1(_09295_),
    .B2(\rvcpu.dp.plem.WriteDataM[15] ),
    .C1(_09328_),
    .X(_09329_));
 sky130_fd_sc_hd__clkbuf_2 _22123_ (.A(_09329_),
    .X(_09330_));
 sky130_fd_sc_hd__mux2_1 _22124_ (.A0(_09330_),
    .A1(\datamem.data_ram[61][31] ),
    .S(_09302_),
    .X(_09331_));
 sky130_fd_sc_hd__clkbuf_1 _22125_ (.A(_09331_),
    .X(_01083_));
 sky130_fd_sc_hd__a21oi_4 _22126_ (.A1(_09299_),
    .A2(_09229_),
    .B1(_09231_),
    .Y(_09332_));
 sky130_fd_sc_hd__mux2_1 _22127_ (.A0(_09224_),
    .A1(\datamem.data_ram[61][16] ),
    .S(_09332_),
    .X(_09333_));
 sky130_fd_sc_hd__clkbuf_1 _22128_ (.A(_09333_),
    .X(_01084_));
 sky130_fd_sc_hd__mux2_1 _22129_ (.A0(_09236_),
    .A1(\datamem.data_ram[61][17] ),
    .S(_09332_),
    .X(_09334_));
 sky130_fd_sc_hd__clkbuf_1 _22130_ (.A(_09334_),
    .X(_01085_));
 sky130_fd_sc_hd__mux2_1 _22131_ (.A0(_09240_),
    .A1(\datamem.data_ram[61][18] ),
    .S(_09332_),
    .X(_09335_));
 sky130_fd_sc_hd__clkbuf_1 _22132_ (.A(_09335_),
    .X(_01086_));
 sky130_fd_sc_hd__mux2_1 _22133_ (.A0(_09244_),
    .A1(\datamem.data_ram[61][19] ),
    .S(_09332_),
    .X(_09336_));
 sky130_fd_sc_hd__clkbuf_1 _22134_ (.A(_09336_),
    .X(_01087_));
 sky130_fd_sc_hd__mux2_1 _22135_ (.A0(_09248_),
    .A1(\datamem.data_ram[61][20] ),
    .S(_09332_),
    .X(_09337_));
 sky130_fd_sc_hd__clkbuf_1 _22136_ (.A(_09337_),
    .X(_01088_));
 sky130_fd_sc_hd__mux2_1 _22137_ (.A0(_09252_),
    .A1(\datamem.data_ram[61][21] ),
    .S(_09332_),
    .X(_09338_));
 sky130_fd_sc_hd__clkbuf_1 _22138_ (.A(_09338_),
    .X(_01089_));
 sky130_fd_sc_hd__mux2_1 _22139_ (.A0(_09256_),
    .A1(\datamem.data_ram[61][22] ),
    .S(_09332_),
    .X(_09339_));
 sky130_fd_sc_hd__clkbuf_1 _22140_ (.A(_09339_),
    .X(_01090_));
 sky130_fd_sc_hd__mux2_1 _22141_ (.A0(_09260_),
    .A1(\datamem.data_ram[61][23] ),
    .S(_09332_),
    .X(_09340_));
 sky130_fd_sc_hd__clkbuf_1 _22142_ (.A(_09340_),
    .X(_01091_));
 sky130_fd_sc_hd__a21oi_1 _22143_ (.A1(_09299_),
    .A2(_09269_),
    .B1(_09231_),
    .Y(_09341_));
 sky130_fd_sc_hd__mux2_1 _22144_ (.A0(_09267_),
    .A1(\datamem.data_ram[61][8] ),
    .S(net62),
    .X(_09342_));
 sky130_fd_sc_hd__clkbuf_1 _22145_ (.A(_09342_),
    .X(_01092_));
 sky130_fd_sc_hd__mux2_1 _22146_ (.A0(_09273_),
    .A1(\datamem.data_ram[61][9] ),
    .S(net62),
    .X(_09343_));
 sky130_fd_sc_hd__clkbuf_1 _22147_ (.A(_09343_),
    .X(_01093_));
 sky130_fd_sc_hd__mux2_1 _22148_ (.A0(_09276_),
    .A1(\datamem.data_ram[61][10] ),
    .S(net62),
    .X(_09344_));
 sky130_fd_sc_hd__clkbuf_1 _22149_ (.A(_09344_),
    .X(_01094_));
 sky130_fd_sc_hd__mux2_1 _22150_ (.A0(_09279_),
    .A1(\datamem.data_ram[61][11] ),
    .S(net62),
    .X(_09345_));
 sky130_fd_sc_hd__clkbuf_1 _22151_ (.A(_09345_),
    .X(_01095_));
 sky130_fd_sc_hd__mux2_1 _22152_ (.A0(_09282_),
    .A1(\datamem.data_ram[61][12] ),
    .S(net62),
    .X(_09346_));
 sky130_fd_sc_hd__clkbuf_1 _22153_ (.A(_09346_),
    .X(_01096_));
 sky130_fd_sc_hd__mux2_1 _22154_ (.A0(_09285_),
    .A1(\datamem.data_ram[61][13] ),
    .S(net62),
    .X(_09347_));
 sky130_fd_sc_hd__clkbuf_1 _22155_ (.A(_09347_),
    .X(_01097_));
 sky130_fd_sc_hd__mux2_1 _22156_ (.A0(_09288_),
    .A1(\datamem.data_ram[61][14] ),
    .S(net62),
    .X(_09348_));
 sky130_fd_sc_hd__clkbuf_1 _22157_ (.A(_09348_),
    .X(_01098_));
 sky130_fd_sc_hd__mux2_1 _22158_ (.A0(_09291_),
    .A1(\datamem.data_ram[61][15] ),
    .S(net62),
    .X(_09349_));
 sky130_fd_sc_hd__clkbuf_1 _22159_ (.A(_09349_),
    .X(_01099_));
 sky130_fd_sc_hd__buf_12 _22160_ (.A(_07123_),
    .X(_09350_));
 sky130_fd_sc_hd__buf_8 _22161_ (.A(_09350_),
    .X(_09351_));
 sky130_fd_sc_hd__a21oi_4 _22162_ (.A1(_09351_),
    .A2(_09301_),
    .B1(_09231_),
    .Y(_09352_));
 sky130_fd_sc_hd__mux2_1 _22163_ (.A0(_09298_),
    .A1(\datamem.data_ram[60][24] ),
    .S(_09352_),
    .X(_09353_));
 sky130_fd_sc_hd__clkbuf_1 _22164_ (.A(_09353_),
    .X(_01100_));
 sky130_fd_sc_hd__mux2_1 _22165_ (.A0(_09306_),
    .A1(\datamem.data_ram[60][25] ),
    .S(_09352_),
    .X(_09354_));
 sky130_fd_sc_hd__clkbuf_1 _22166_ (.A(_09354_),
    .X(_01101_));
 sky130_fd_sc_hd__mux2_1 _22167_ (.A0(_09310_),
    .A1(\datamem.data_ram[60][26] ),
    .S(_09352_),
    .X(_09355_));
 sky130_fd_sc_hd__clkbuf_1 _22168_ (.A(_09355_),
    .X(_01102_));
 sky130_fd_sc_hd__mux2_1 _22169_ (.A0(_09314_),
    .A1(\datamem.data_ram[60][27] ),
    .S(_09352_),
    .X(_09356_));
 sky130_fd_sc_hd__clkbuf_1 _22170_ (.A(_09356_),
    .X(_01103_));
 sky130_fd_sc_hd__mux2_1 _22171_ (.A0(_09318_),
    .A1(\datamem.data_ram[60][28] ),
    .S(_09352_),
    .X(_09357_));
 sky130_fd_sc_hd__clkbuf_1 _22172_ (.A(_09357_),
    .X(_01104_));
 sky130_fd_sc_hd__mux2_1 _22173_ (.A0(_09322_),
    .A1(\datamem.data_ram[60][29] ),
    .S(_09352_),
    .X(_09358_));
 sky130_fd_sc_hd__clkbuf_1 _22174_ (.A(_09358_),
    .X(_01105_));
 sky130_fd_sc_hd__mux2_1 _22175_ (.A0(_09326_),
    .A1(\datamem.data_ram[60][30] ),
    .S(_09352_),
    .X(_09359_));
 sky130_fd_sc_hd__clkbuf_1 _22176_ (.A(_09359_),
    .X(_01106_));
 sky130_fd_sc_hd__mux2_1 _22177_ (.A0(_09330_),
    .A1(\datamem.data_ram[60][31] ),
    .S(_09352_),
    .X(_09360_));
 sky130_fd_sc_hd__clkbuf_1 _22178_ (.A(_09360_),
    .X(_01107_));
 sky130_fd_sc_hd__buf_8 _22179_ (.A(_09230_),
    .X(_09361_));
 sky130_fd_sc_hd__a21oi_4 _22180_ (.A1(_09351_),
    .A2(_09229_),
    .B1(_09361_),
    .Y(_09362_));
 sky130_fd_sc_hd__mux2_1 _22181_ (.A0(_09224_),
    .A1(\datamem.data_ram[60][16] ),
    .S(_09362_),
    .X(_09363_));
 sky130_fd_sc_hd__clkbuf_1 _22182_ (.A(_09363_),
    .X(_01108_));
 sky130_fd_sc_hd__mux2_1 _22183_ (.A0(_09236_),
    .A1(\datamem.data_ram[60][17] ),
    .S(_09362_),
    .X(_09364_));
 sky130_fd_sc_hd__clkbuf_1 _22184_ (.A(_09364_),
    .X(_01109_));
 sky130_fd_sc_hd__mux2_1 _22185_ (.A0(_09240_),
    .A1(\datamem.data_ram[60][18] ),
    .S(_09362_),
    .X(_09365_));
 sky130_fd_sc_hd__clkbuf_1 _22186_ (.A(_09365_),
    .X(_01110_));
 sky130_fd_sc_hd__mux2_1 _22187_ (.A0(_09244_),
    .A1(\datamem.data_ram[60][19] ),
    .S(_09362_),
    .X(_09366_));
 sky130_fd_sc_hd__clkbuf_1 _22188_ (.A(_09366_),
    .X(_01111_));
 sky130_fd_sc_hd__mux2_1 _22189_ (.A0(_09248_),
    .A1(\datamem.data_ram[60][20] ),
    .S(_09362_),
    .X(_09367_));
 sky130_fd_sc_hd__clkbuf_1 _22190_ (.A(_09367_),
    .X(_01112_));
 sky130_fd_sc_hd__mux2_1 _22191_ (.A0(_09252_),
    .A1(\datamem.data_ram[60][21] ),
    .S(_09362_),
    .X(_09368_));
 sky130_fd_sc_hd__clkbuf_1 _22192_ (.A(_09368_),
    .X(_01113_));
 sky130_fd_sc_hd__mux2_1 _22193_ (.A0(_09256_),
    .A1(\datamem.data_ram[60][22] ),
    .S(_09362_),
    .X(_09369_));
 sky130_fd_sc_hd__clkbuf_1 _22194_ (.A(_09369_),
    .X(_01114_));
 sky130_fd_sc_hd__mux2_1 _22195_ (.A0(_09260_),
    .A1(\datamem.data_ram[60][23] ),
    .S(_09362_),
    .X(_09370_));
 sky130_fd_sc_hd__clkbuf_1 _22196_ (.A(_09370_),
    .X(_01115_));
 sky130_fd_sc_hd__a21oi_4 _22197_ (.A1(_09351_),
    .A2(_09269_),
    .B1(_09361_),
    .Y(_09371_));
 sky130_fd_sc_hd__mux2_1 _22198_ (.A0(_09267_),
    .A1(\datamem.data_ram[60][8] ),
    .S(_09371_),
    .X(_09372_));
 sky130_fd_sc_hd__clkbuf_1 _22199_ (.A(_09372_),
    .X(_01116_));
 sky130_fd_sc_hd__mux2_1 _22200_ (.A0(_09273_),
    .A1(\datamem.data_ram[60][9] ),
    .S(_09371_),
    .X(_09373_));
 sky130_fd_sc_hd__clkbuf_1 _22201_ (.A(_09373_),
    .X(_01117_));
 sky130_fd_sc_hd__mux2_1 _22202_ (.A0(_09276_),
    .A1(\datamem.data_ram[60][10] ),
    .S(_09371_),
    .X(_09374_));
 sky130_fd_sc_hd__clkbuf_1 _22203_ (.A(_09374_),
    .X(_01118_));
 sky130_fd_sc_hd__mux2_1 _22204_ (.A0(_09279_),
    .A1(\datamem.data_ram[60][11] ),
    .S(_09371_),
    .X(_09375_));
 sky130_fd_sc_hd__clkbuf_1 _22205_ (.A(_09375_),
    .X(_01119_));
 sky130_fd_sc_hd__mux2_1 _22206_ (.A0(_09282_),
    .A1(\datamem.data_ram[60][12] ),
    .S(_09371_),
    .X(_09376_));
 sky130_fd_sc_hd__clkbuf_1 _22207_ (.A(_09376_),
    .X(_01120_));
 sky130_fd_sc_hd__mux2_1 _22208_ (.A0(_09285_),
    .A1(\datamem.data_ram[60][13] ),
    .S(_09371_),
    .X(_09377_));
 sky130_fd_sc_hd__clkbuf_1 _22209_ (.A(_09377_),
    .X(_01121_));
 sky130_fd_sc_hd__mux2_1 _22210_ (.A0(_09288_),
    .A1(\datamem.data_ram[60][14] ),
    .S(_09371_),
    .X(_09378_));
 sky130_fd_sc_hd__clkbuf_1 _22211_ (.A(_09378_),
    .X(_01122_));
 sky130_fd_sc_hd__mux2_1 _22212_ (.A0(_09291_),
    .A1(\datamem.data_ram[60][15] ),
    .S(_09371_),
    .X(_09379_));
 sky130_fd_sc_hd__clkbuf_1 _22213_ (.A(_09379_),
    .X(_01123_));
 sky130_fd_sc_hd__buf_4 _22214_ (.A(\rvcpu.dp.plfd.InstrD[22] ),
    .X(_09380_));
 sky130_fd_sc_hd__buf_4 _22215_ (.A(_08595_),
    .X(_09381_));
 sky130_fd_sc_hd__clkbuf_8 _22216_ (.A(_09381_),
    .X(_09382_));
 sky130_fd_sc_hd__clkbuf_4 _22217_ (.A(_09382_),
    .X(_09383_));
 sky130_fd_sc_hd__clkbuf_8 _22218_ (.A(_08592_),
    .X(_09384_));
 sky130_fd_sc_hd__buf_8 _22219_ (.A(_09384_),
    .X(_09385_));
 sky130_fd_sc_hd__buf_6 _22220_ (.A(_09385_),
    .X(_09386_));
 sky130_fd_sc_hd__or2_2 _22221_ (.A(\rvcpu.dp.plfd.InstrD[24] ),
    .B(\rvcpu.dp.plfd.InstrD[23] ),
    .X(_09387_));
 sky130_fd_sc_hd__o41a_1 _22222_ (.A1(_09380_),
    .A2(_09383_),
    .A3(_09386_),
    .A4(_09387_),
    .B1(_08622_),
    .X(_09388_));
 sky130_fd_sc_hd__clkbuf_4 _22223_ (.A(_09388_),
    .X(_09389_));
 sky130_fd_sc_hd__clkbuf_4 _22224_ (.A(\rvcpu.dp.plfd.InstrD[22] ),
    .X(_09390_));
 sky130_fd_sc_hd__clkbuf_4 _22225_ (.A(_09390_),
    .X(_09391_));
 sky130_fd_sc_hd__clkbuf_8 _22226_ (.A(_08592_),
    .X(_09392_));
 sky130_fd_sc_hd__buf_4 _22227_ (.A(_09392_),
    .X(_09393_));
 sky130_fd_sc_hd__buf_4 _22228_ (.A(_08595_),
    .X(_09394_));
 sky130_fd_sc_hd__buf_4 _22229_ (.A(_09394_),
    .X(_09395_));
 sky130_fd_sc_hd__mux4_1 _22230_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][0] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][0] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][0] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][0] ),
    .S0(_09393_),
    .S1(_09395_),
    .X(_09396_));
 sky130_fd_sc_hd__or2_1 _22231_ (.A(_09391_),
    .B(_09396_),
    .X(_09397_));
 sky130_fd_sc_hd__inv_2 _22232_ (.A(\rvcpu.dp.plfd.InstrD[22] ),
    .Y(_09398_));
 sky130_fd_sc_hd__buf_4 _22233_ (.A(_09398_),
    .X(_09399_));
 sky130_fd_sc_hd__clkbuf_8 _22234_ (.A(_08595_),
    .X(_09400_));
 sky130_fd_sc_hd__clkbuf_8 _22235_ (.A(_08592_),
    .X(_09401_));
 sky130_fd_sc_hd__buf_4 _22236_ (.A(_09401_),
    .X(_09402_));
 sky130_fd_sc_hd__mux4_1 _22237_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][0] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][0] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][0] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][0] ),
    .S0(_09400_),
    .S1(_09402_),
    .X(_09403_));
 sky130_fd_sc_hd__clkbuf_4 _22238_ (.A(\rvcpu.dp.plfd.InstrD[23] ),
    .X(_09404_));
 sky130_fd_sc_hd__o21a_1 _22239_ (.A1(_09399_),
    .A2(_09403_),
    .B1(_09404_),
    .X(_09405_));
 sky130_fd_sc_hd__buf_6 _22240_ (.A(_08592_),
    .X(_09406_));
 sky130_fd_sc_hd__mux4_1 _22241_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][0] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][0] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][0] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][0] ),
    .S0(_09406_),
    .S1(_09395_),
    .X(_09407_));
 sky130_fd_sc_hd__buf_4 _22242_ (.A(_09394_),
    .X(_09408_));
 sky130_fd_sc_hd__mux4_1 _22243_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][0] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][0] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][0] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][0] ),
    .S0(_09406_),
    .S1(_09408_),
    .X(_09409_));
 sky130_fd_sc_hd__mux2_1 _22244_ (.A0(_09407_),
    .A1(_09409_),
    .S(_09380_),
    .X(_09410_));
 sky130_fd_sc_hd__inv_2 _22245_ (.A(\rvcpu.dp.plfd.InstrD[23] ),
    .Y(_09411_));
 sky130_fd_sc_hd__clkbuf_4 _22246_ (.A(_09411_),
    .X(_09412_));
 sky130_fd_sc_hd__clkbuf_4 _22247_ (.A(_08589_),
    .X(_09413_));
 sky130_fd_sc_hd__a221o_1 _22248_ (.A1(_09397_),
    .A2(_09405_),
    .B1(_09410_),
    .B2(_09412_),
    .C1(_09413_),
    .X(_09414_));
 sky130_fd_sc_hd__buf_4 _22249_ (.A(_09399_),
    .X(_09415_));
 sky130_fd_sc_hd__buf_4 _22250_ (.A(_09401_),
    .X(_09416_));
 sky130_fd_sc_hd__clkbuf_8 _22251_ (.A(_09416_),
    .X(_09417_));
 sky130_fd_sc_hd__clkbuf_8 _22252_ (.A(_09400_),
    .X(_09418_));
 sky130_fd_sc_hd__clkbuf_8 _22253_ (.A(_09418_),
    .X(_09419_));
 sky130_fd_sc_hd__mux4_1 _22254_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][0] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][0] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][0] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][0] ),
    .S0(_09417_),
    .S1(_09419_),
    .X(_09420_));
 sky130_fd_sc_hd__clkbuf_8 _22255_ (.A(\rvcpu.dp.plfd.InstrD[22] ),
    .X(_09421_));
 sky130_fd_sc_hd__buf_4 _22256_ (.A(_09421_),
    .X(_09422_));
 sky130_fd_sc_hd__clkbuf_8 _22257_ (.A(_09401_),
    .X(_09423_));
 sky130_fd_sc_hd__clkbuf_8 _22258_ (.A(_09400_),
    .X(_09424_));
 sky130_fd_sc_hd__mux4_1 _22259_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][0] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][0] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][0] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][0] ),
    .S0(_09423_),
    .S1(_09424_),
    .X(_09425_));
 sky130_fd_sc_hd__clkbuf_4 _22260_ (.A(_09387_),
    .X(_09426_));
 sky130_fd_sc_hd__a21o_1 _22261_ (.A1(_09422_),
    .A2(_09425_),
    .B1(_09426_),
    .X(_09427_));
 sky130_fd_sc_hd__a21o_1 _22262_ (.A1(_09415_),
    .A2(_09420_),
    .B1(_09427_),
    .X(_09428_));
 sky130_fd_sc_hd__clkbuf_4 _22263_ (.A(_09399_),
    .X(_09429_));
 sky130_fd_sc_hd__buf_4 _22264_ (.A(_08595_),
    .X(_09430_));
 sky130_fd_sc_hd__clkbuf_8 _22265_ (.A(_09430_),
    .X(_09431_));
 sky130_fd_sc_hd__mux4_1 _22266_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][0] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][0] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][0] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][0] ),
    .S0(_09431_),
    .S1(_09386_),
    .X(_09432_));
 sky130_fd_sc_hd__clkbuf_4 _22267_ (.A(_09421_),
    .X(_09433_));
 sky130_fd_sc_hd__clkbuf_8 _22268_ (.A(_09392_),
    .X(_09434_));
 sky130_fd_sc_hd__mux4_1 _22269_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][0] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][0] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][0] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][0] ),
    .S0(_09434_),
    .S1(_09382_),
    .X(_09435_));
 sky130_fd_sc_hd__and2_1 _22270_ (.A(_09433_),
    .B(_09435_),
    .X(_09436_));
 sky130_fd_sc_hd__nand2_2 _22271_ (.A(_08589_),
    .B(_09404_),
    .Y(_09437_));
 sky130_fd_sc_hd__clkbuf_4 _22272_ (.A(_09437_),
    .X(_09438_));
 sky130_fd_sc_hd__a211o_1 _22273_ (.A1(_09429_),
    .A2(_09432_),
    .B1(_09436_),
    .C1(_09438_),
    .X(_09439_));
 sky130_fd_sc_hd__and4_1 _22274_ (.A(_09389_),
    .B(_09414_),
    .C(_09428_),
    .D(_09439_),
    .X(_09440_));
 sky130_fd_sc_hd__clkbuf_1 _22275_ (.A(_09440_),
    .X(_01124_));
 sky130_fd_sc_hd__buf_2 _22276_ (.A(_09413_),
    .X(_09441_));
 sky130_fd_sc_hd__buf_2 _22277_ (.A(_09411_),
    .X(_09442_));
 sky130_fd_sc_hd__clkbuf_8 _22278_ (.A(_09381_),
    .X(_09443_));
 sky130_fd_sc_hd__mux4_1 _22279_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][1] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][1] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][1] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][1] ),
    .S0(_09416_),
    .S1(_09443_),
    .X(_09444_));
 sky130_fd_sc_hd__buf_4 _22280_ (.A(_09401_),
    .X(_09445_));
 sky130_fd_sc_hd__clkbuf_8 _22281_ (.A(_08595_),
    .X(_09446_));
 sky130_fd_sc_hd__buf_4 _22282_ (.A(_09446_),
    .X(_09447_));
 sky130_fd_sc_hd__mux4_1 _22283_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][1] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][1] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][1] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][1] ),
    .S0(_09445_),
    .S1(_09447_),
    .X(_09448_));
 sky130_fd_sc_hd__buf_4 _22284_ (.A(_09421_),
    .X(_09449_));
 sky130_fd_sc_hd__mux2_1 _22285_ (.A0(_09444_),
    .A1(_09448_),
    .S(_09449_),
    .X(_09450_));
 sky130_fd_sc_hd__clkbuf_4 _22286_ (.A(_09398_),
    .X(_09451_));
 sky130_fd_sc_hd__buf_4 _22287_ (.A(_09451_),
    .X(_09452_));
 sky130_fd_sc_hd__buf_4 _22288_ (.A(_09423_),
    .X(_09453_));
 sky130_fd_sc_hd__mux4_1 _22289_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][1] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][1] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][1] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][1] ),
    .S0(_09443_),
    .S1(_09453_),
    .X(_09454_));
 sky130_fd_sc_hd__nor2_1 _22290_ (.A(_09452_),
    .B(_09454_),
    .Y(_09455_));
 sky130_fd_sc_hd__mux4_1 _22291_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][1] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][1] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][1] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][1] ),
    .S0(_09385_),
    .S1(_09431_),
    .X(_09456_));
 sky130_fd_sc_hd__buf_4 _22292_ (.A(_09404_),
    .X(_09457_));
 sky130_fd_sc_hd__o21ai_1 _22293_ (.A1(_09422_),
    .A2(_09456_),
    .B1(_09457_),
    .Y(_09458_));
 sky130_fd_sc_hd__o2bb2a_1 _22294_ (.A1_N(_09442_),
    .A2_N(_09450_),
    .B1(_09455_),
    .B2(_09458_),
    .X(_09459_));
 sky130_fd_sc_hd__nor2_1 _22295_ (.A(_09441_),
    .B(_09459_),
    .Y(_09460_));
 sky130_fd_sc_hd__buf_4 _22296_ (.A(_09452_),
    .X(_09461_));
 sky130_fd_sc_hd__buf_4 _22297_ (.A(_09392_),
    .X(_09462_));
 sky130_fd_sc_hd__clkbuf_8 _22298_ (.A(_09462_),
    .X(_09463_));
 sky130_fd_sc_hd__buf_6 _22299_ (.A(_09463_),
    .X(_09464_));
 sky130_fd_sc_hd__buf_4 _22300_ (.A(_09381_),
    .X(_09465_));
 sky130_fd_sc_hd__buf_4 _22301_ (.A(_09465_),
    .X(_09466_));
 sky130_fd_sc_hd__clkbuf_8 _22302_ (.A(_09466_),
    .X(_09467_));
 sky130_fd_sc_hd__mux4_1 _22303_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][1] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][1] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][1] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][1] ),
    .S0(_09464_),
    .S1(_09467_),
    .X(_09468_));
 sky130_fd_sc_hd__clkbuf_4 _22304_ (.A(_09391_),
    .X(_09469_));
 sky130_fd_sc_hd__mux4_1 _22305_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][1] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][1] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][1] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][1] ),
    .S0(_09463_),
    .S1(_09466_),
    .X(_09470_));
 sky130_fd_sc_hd__or2_1 _22306_ (.A(_09469_),
    .B(_09470_),
    .X(_09471_));
 sky130_fd_sc_hd__clkbuf_4 _22307_ (.A(\rvcpu.dp.plfd.InstrD[23] ),
    .X(_09472_));
 sky130_fd_sc_hd__nor2_1 _22308_ (.A(\rvcpu.dp.plfd.InstrD[24] ),
    .B(_09472_),
    .Y(_09473_));
 sky130_fd_sc_hd__clkbuf_4 _22309_ (.A(_09473_),
    .X(_09474_));
 sky130_fd_sc_hd__o211a_1 _22310_ (.A1(_09461_),
    .A2(_09468_),
    .B1(_09471_),
    .C1(_09474_),
    .X(_09475_));
 sky130_fd_sc_hd__clkbuf_8 _22311_ (.A(_09452_),
    .X(_09476_));
 sky130_fd_sc_hd__buf_4 _22312_ (.A(_09462_),
    .X(_09477_));
 sky130_fd_sc_hd__buf_6 _22313_ (.A(_09477_),
    .X(_09478_));
 sky130_fd_sc_hd__buf_6 _22314_ (.A(_09383_),
    .X(_09479_));
 sky130_fd_sc_hd__mux4_1 _22315_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][1] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][1] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][1] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][1] ),
    .S0(_09478_),
    .S1(_09479_),
    .X(_09480_));
 sky130_fd_sc_hd__buf_2 _22316_ (.A(_09390_),
    .X(_09481_));
 sky130_fd_sc_hd__buf_4 _22317_ (.A(_09481_),
    .X(_09482_));
 sky130_fd_sc_hd__buf_4 _22318_ (.A(_09400_),
    .X(_09483_));
 sky130_fd_sc_hd__clkbuf_8 _22319_ (.A(_09401_),
    .X(_09484_));
 sky130_fd_sc_hd__buf_4 _22320_ (.A(_09484_),
    .X(_09485_));
 sky130_fd_sc_hd__mux4_1 _22321_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][1] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][1] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][1] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][1] ),
    .S0(_09483_),
    .S1(_09485_),
    .X(_09486_));
 sky130_fd_sc_hd__or2_1 _22322_ (.A(_09482_),
    .B(_09486_),
    .X(_09487_));
 sky130_fd_sc_hd__nor2_2 _22323_ (.A(\rvcpu.dp.plfd.InstrD[24] ),
    .B(_09411_),
    .Y(_09488_));
 sky130_fd_sc_hd__buf_2 _22324_ (.A(_09488_),
    .X(_09489_));
 sky130_fd_sc_hd__o211a_1 _22325_ (.A1(_09476_),
    .A2(_09480_),
    .B1(_09487_),
    .C1(_09489_),
    .X(_09490_));
 sky130_fd_sc_hd__clkbuf_4 _22326_ (.A(_09389_),
    .X(_09491_));
 sky130_fd_sc_hd__o31a_1 _22327_ (.A1(_09460_),
    .A2(_09475_),
    .A3(_09490_),
    .B1(_09491_),
    .X(_01125_));
 sky130_fd_sc_hd__mux4_1 _22328_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][2] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][2] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][2] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][2] ),
    .S0(_09416_),
    .S1(_09443_),
    .X(_09492_));
 sky130_fd_sc_hd__mux4_1 _22329_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][2] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][2] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][2] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][2] ),
    .S0(_09445_),
    .S1(_09447_),
    .X(_09493_));
 sky130_fd_sc_hd__mux2_1 _22330_ (.A0(_09492_),
    .A1(_09493_),
    .S(_09449_),
    .X(_09494_));
 sky130_fd_sc_hd__clkbuf_4 _22331_ (.A(_09398_),
    .X(_09495_));
 sky130_fd_sc_hd__mux4_1 _22332_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][2] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][2] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][2] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][2] ),
    .S0(_09443_),
    .S1(_09453_),
    .X(_09496_));
 sky130_fd_sc_hd__nor2_1 _22333_ (.A(_09495_),
    .B(_09496_),
    .Y(_09497_));
 sky130_fd_sc_hd__mux4_1 _22334_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][2] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][2] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][2] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][2] ),
    .S0(_09385_),
    .S1(_09431_),
    .X(_09498_));
 sky130_fd_sc_hd__o21ai_1 _22335_ (.A1(_09422_),
    .A2(_09498_),
    .B1(_09457_),
    .Y(_09499_));
 sky130_fd_sc_hd__o2bb2a_1 _22336_ (.A1_N(_09442_),
    .A2_N(_09494_),
    .B1(_09497_),
    .B2(_09499_),
    .X(_09500_));
 sky130_fd_sc_hd__nor2_1 _22337_ (.A(_09441_),
    .B(_09500_),
    .Y(_09501_));
 sky130_fd_sc_hd__mux4_1 _22338_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][2] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][2] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][2] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][2] ),
    .S0(_09464_),
    .S1(_09467_),
    .X(_09502_));
 sky130_fd_sc_hd__mux4_1 _22339_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][2] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][2] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][2] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][2] ),
    .S0(_09463_),
    .S1(_09466_),
    .X(_09503_));
 sky130_fd_sc_hd__or2_1 _22340_ (.A(_09469_),
    .B(_09503_),
    .X(_09504_));
 sky130_fd_sc_hd__o211a_1 _22341_ (.A1(_09461_),
    .A2(_09502_),
    .B1(_09504_),
    .C1(_09474_),
    .X(_09505_));
 sky130_fd_sc_hd__mux4_1 _22342_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][2] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][2] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][2] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][2] ),
    .S0(_09478_),
    .S1(_09479_),
    .X(_09506_));
 sky130_fd_sc_hd__mux4_1 _22343_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][2] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][2] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][2] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][2] ),
    .S0(_09483_),
    .S1(_09485_),
    .X(_09507_));
 sky130_fd_sc_hd__or2_1 _22344_ (.A(_09482_),
    .B(_09507_),
    .X(_09508_));
 sky130_fd_sc_hd__o211a_1 _22345_ (.A1(_09476_),
    .A2(_09506_),
    .B1(_09508_),
    .C1(_09489_),
    .X(_09509_));
 sky130_fd_sc_hd__o31a_1 _22346_ (.A1(_09501_),
    .A2(_09505_),
    .A3(_09509_),
    .B1(_09491_),
    .X(_01126_));
 sky130_fd_sc_hd__buf_2 _22347_ (.A(_09411_),
    .X(_09510_));
 sky130_fd_sc_hd__clkbuf_4 _22348_ (.A(\rvcpu.dp.plfd.InstrD[22] ),
    .X(_09511_));
 sky130_fd_sc_hd__clkbuf_8 _22349_ (.A(_08592_),
    .X(_09512_));
 sky130_fd_sc_hd__buf_4 _22350_ (.A(_09394_),
    .X(_09513_));
 sky130_fd_sc_hd__mux4_1 _22351_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][3] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][3] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][3] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][3] ),
    .S0(_09512_),
    .S1(_09513_),
    .X(_09514_));
 sky130_fd_sc_hd__or2_1 _22352_ (.A(_09511_),
    .B(_09514_),
    .X(_09515_));
 sky130_fd_sc_hd__clkbuf_4 _22353_ (.A(_09398_),
    .X(_09516_));
 sky130_fd_sc_hd__clkbuf_8 _22354_ (.A(_08592_),
    .X(_09517_));
 sky130_fd_sc_hd__mux4_1 _22355_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][3] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][3] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][3] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][3] ),
    .S0(_09517_),
    .S1(_09513_),
    .X(_09518_));
 sky130_fd_sc_hd__or2_1 _22356_ (.A(_09516_),
    .B(_09518_),
    .X(_09519_));
 sky130_fd_sc_hd__mux4_1 _22357_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][3] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][3] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][3] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][3] ),
    .S0(_09446_),
    .S1(_09402_),
    .X(_09520_));
 sky130_fd_sc_hd__mux4_1 _22358_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][3] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][3] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][3] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][3] ),
    .S0(_09392_),
    .S1(_09394_),
    .X(_09521_));
 sky130_fd_sc_hd__or2_1 _22359_ (.A(_09390_),
    .B(_09521_),
    .X(_09522_));
 sky130_fd_sc_hd__clkbuf_4 _22360_ (.A(_09404_),
    .X(_09523_));
 sky130_fd_sc_hd__o211a_1 _22361_ (.A1(_09451_),
    .A2(_09520_),
    .B1(_09522_),
    .C1(_09523_),
    .X(_09524_));
 sky130_fd_sc_hd__clkbuf_4 _22362_ (.A(_08589_),
    .X(_09525_));
 sky130_fd_sc_hd__a311o_2 _22363_ (.A1(_09510_),
    .A2(_09515_),
    .A3(_09519_),
    .B1(_09524_),
    .C1(_09525_),
    .X(_09526_));
 sky130_fd_sc_hd__mux4_1 _22364_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][3] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][3] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][3] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][3] ),
    .S0(_09417_),
    .S1(_09419_),
    .X(_09527_));
 sky130_fd_sc_hd__clkbuf_4 _22365_ (.A(_09421_),
    .X(_09528_));
 sky130_fd_sc_hd__mux4_1 _22366_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][3] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][3] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][3] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][3] ),
    .S0(_09423_),
    .S1(_09424_),
    .X(_09529_));
 sky130_fd_sc_hd__a21o_1 _22367_ (.A1(_09528_),
    .A2(_09529_),
    .B1(_09426_),
    .X(_09530_));
 sky130_fd_sc_hd__a21o_1 _22368_ (.A1(_09415_),
    .A2(_09527_),
    .B1(_09530_),
    .X(_09531_));
 sky130_fd_sc_hd__clkbuf_4 _22369_ (.A(_09385_),
    .X(_09532_));
 sky130_fd_sc_hd__mux4_1 _22370_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][3] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][3] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][3] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][3] ),
    .S0(_09431_),
    .S1(_09532_),
    .X(_09533_));
 sky130_fd_sc_hd__clkbuf_2 _22371_ (.A(_09421_),
    .X(_09534_));
 sky130_fd_sc_hd__mux4_1 _22372_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][3] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][3] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][3] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][3] ),
    .S0(_09434_),
    .S1(_09382_),
    .X(_09535_));
 sky130_fd_sc_hd__and2_1 _22373_ (.A(_09534_),
    .B(_09535_),
    .X(_09536_));
 sky130_fd_sc_hd__a211o_1 _22374_ (.A1(_09429_),
    .A2(_09533_),
    .B1(_09536_),
    .C1(_09438_),
    .X(_09537_));
 sky130_fd_sc_hd__and4_1 _22375_ (.A(_09389_),
    .B(_09526_),
    .C(_09531_),
    .D(_09537_),
    .X(_09538_));
 sky130_fd_sc_hd__clkbuf_1 _22376_ (.A(_09538_),
    .X(_01127_));
 sky130_fd_sc_hd__mux4_1 _22377_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][4] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][4] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][4] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][4] ),
    .S0(_09393_),
    .S1(_09395_),
    .X(_09539_));
 sky130_fd_sc_hd__or2_1 _22378_ (.A(_09391_),
    .B(_09539_),
    .X(_09540_));
 sky130_fd_sc_hd__mux4_1 _22379_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][4] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][4] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][4] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][4] ),
    .S0(_09446_),
    .S1(_09402_),
    .X(_09541_));
 sky130_fd_sc_hd__o21a_1 _22380_ (.A1(_09451_),
    .A2(_09541_),
    .B1(_09404_),
    .X(_09542_));
 sky130_fd_sc_hd__mux4_1 _22381_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][4] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][4] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][4] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][4] ),
    .S0(_09406_),
    .S1(_09395_),
    .X(_09543_));
 sky130_fd_sc_hd__mux4_1 _22382_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][4] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][4] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][4] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][4] ),
    .S0(_09512_),
    .S1(_09408_),
    .X(_09544_));
 sky130_fd_sc_hd__mux2_2 _22383_ (.A0(_09543_),
    .A1(_09544_),
    .S(_09380_),
    .X(_09545_));
 sky130_fd_sc_hd__a221o_1 _22384_ (.A1(_09540_),
    .A2(_09542_),
    .B1(_09545_),
    .B2(_09412_),
    .C1(_09413_),
    .X(_09546_));
 sky130_fd_sc_hd__mux4_1 _22385_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][4] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][4] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][4] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][4] ),
    .S0(_09417_),
    .S1(_09419_),
    .X(_09547_));
 sky130_fd_sc_hd__mux4_1 _22386_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][4] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][4] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][4] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][4] ),
    .S0(_09423_),
    .S1(_09424_),
    .X(_09548_));
 sky130_fd_sc_hd__a21o_1 _22387_ (.A1(_09528_),
    .A2(_09548_),
    .B1(_09426_),
    .X(_09549_));
 sky130_fd_sc_hd__a21o_1 _22388_ (.A1(_09415_),
    .A2(_09547_),
    .B1(_09549_),
    .X(_09550_));
 sky130_fd_sc_hd__mux4_1 _22389_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][4] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][4] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][4] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][4] ),
    .S0(_09431_),
    .S1(_09532_),
    .X(_09551_));
 sky130_fd_sc_hd__buf_4 _22390_ (.A(_09392_),
    .X(_09552_));
 sky130_fd_sc_hd__mux4_1 _22391_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][4] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][4] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][4] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][4] ),
    .S0(_09552_),
    .S1(_09382_),
    .X(_09553_));
 sky130_fd_sc_hd__and2_1 _22392_ (.A(_09534_),
    .B(_09553_),
    .X(_09554_));
 sky130_fd_sc_hd__a211o_1 _22393_ (.A1(_09429_),
    .A2(_09551_),
    .B1(_09554_),
    .C1(_09438_),
    .X(_09555_));
 sky130_fd_sc_hd__and4_1 _22394_ (.A(_09389_),
    .B(_09546_),
    .C(_09550_),
    .D(_09555_),
    .X(_09556_));
 sky130_fd_sc_hd__clkbuf_1 _22395_ (.A(_09556_),
    .X(_01128_));
 sky130_fd_sc_hd__mux4_1 _22396_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][5] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][5] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][5] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][5] ),
    .S0(_09445_),
    .S1(_09447_),
    .X(_09557_));
 sky130_fd_sc_hd__buf_4 _22397_ (.A(_09381_),
    .X(_09558_));
 sky130_fd_sc_hd__mux4_1 _22398_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][5] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][5] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][5] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][5] ),
    .S0(_09434_),
    .S1(_09558_),
    .X(_09559_));
 sky130_fd_sc_hd__mux2_2 _22399_ (.A0(_09557_),
    .A1(_09559_),
    .S(_09449_),
    .X(_09560_));
 sky130_fd_sc_hd__mux4_1 _22400_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][5] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][5] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][5] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][5] ),
    .S0(_09443_),
    .S1(_09453_),
    .X(_09561_));
 sky130_fd_sc_hd__nor2_1 _22401_ (.A(_09495_),
    .B(_09561_),
    .Y(_09562_));
 sky130_fd_sc_hd__mux4_1 _22402_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][5] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][5] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][5] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][5] ),
    .S0(_09484_),
    .S1(_09431_),
    .X(_09563_));
 sky130_fd_sc_hd__o21ai_1 _22403_ (.A1(_09422_),
    .A2(_09563_),
    .B1(_09457_),
    .Y(_09564_));
 sky130_fd_sc_hd__o2bb2a_1 _22404_ (.A1_N(_09442_),
    .A2_N(_09560_),
    .B1(_09562_),
    .B2(_09564_),
    .X(_09565_));
 sky130_fd_sc_hd__nor2_1 _22405_ (.A(_09441_),
    .B(_09565_),
    .Y(_09566_));
 sky130_fd_sc_hd__mux4_1 _22406_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][5] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][5] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][5] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][5] ),
    .S0(_09464_),
    .S1(_09467_),
    .X(_09567_));
 sky130_fd_sc_hd__mux4_1 _22407_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][5] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][5] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][5] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][5] ),
    .S0(_09463_),
    .S1(_09466_),
    .X(_09568_));
 sky130_fd_sc_hd__or2_1 _22408_ (.A(_09469_),
    .B(_09568_),
    .X(_09569_));
 sky130_fd_sc_hd__o211a_1 _22409_ (.A1(_09461_),
    .A2(_09567_),
    .B1(_09569_),
    .C1(_09474_),
    .X(_09570_));
 sky130_fd_sc_hd__mux4_1 _22410_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][5] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][5] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][5] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][5] ),
    .S0(_09478_),
    .S1(_09479_),
    .X(_09571_));
 sky130_fd_sc_hd__mux4_1 _22411_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][5] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][5] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][5] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][5] ),
    .S0(_09483_),
    .S1(_09485_),
    .X(_09572_));
 sky130_fd_sc_hd__or2_1 _22412_ (.A(_09482_),
    .B(_09572_),
    .X(_09573_));
 sky130_fd_sc_hd__o211a_1 _22413_ (.A1(_09476_),
    .A2(_09571_),
    .B1(_09573_),
    .C1(_09489_),
    .X(_09574_));
 sky130_fd_sc_hd__o31a_1 _22414_ (.A1(_09566_),
    .A2(_09570_),
    .A3(_09574_),
    .B1(_09491_),
    .X(_01129_));
 sky130_fd_sc_hd__mux4_2 _22415_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][6] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][6] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][6] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][6] ),
    .S0(_09512_),
    .S1(_09513_),
    .X(_09575_));
 sky130_fd_sc_hd__or2_1 _22416_ (.A(_09511_),
    .B(_09575_),
    .X(_09576_));
 sky130_fd_sc_hd__buf_4 _22417_ (.A(_08595_),
    .X(_09577_));
 sky130_fd_sc_hd__mux4_2 _22418_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][6] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][6] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][6] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][6] ),
    .S0(_09517_),
    .S1(_09577_),
    .X(_09578_));
 sky130_fd_sc_hd__or2_1 _22419_ (.A(_09516_),
    .B(_09578_),
    .X(_09579_));
 sky130_fd_sc_hd__mux4_1 _22420_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][6] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][6] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][6] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][6] ),
    .S0(_09446_),
    .S1(_09402_),
    .X(_09580_));
 sky130_fd_sc_hd__mux4_1 _22421_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][6] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][6] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][6] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][6] ),
    .S0(_09392_),
    .S1(_09394_),
    .X(_09581_));
 sky130_fd_sc_hd__or2_1 _22422_ (.A(_09390_),
    .B(_09581_),
    .X(_09582_));
 sky130_fd_sc_hd__o211a_1 _22423_ (.A1(_09451_),
    .A2(_09580_),
    .B1(_09582_),
    .C1(_09523_),
    .X(_09583_));
 sky130_fd_sc_hd__a311o_2 _22424_ (.A1(_09510_),
    .A2(_09576_),
    .A3(_09579_),
    .B1(_09583_),
    .C1(_09525_),
    .X(_09584_));
 sky130_fd_sc_hd__clkbuf_4 _22425_ (.A(_09418_),
    .X(_09585_));
 sky130_fd_sc_hd__mux4_1 _22426_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][6] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][6] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][6] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][6] ),
    .S0(_09417_),
    .S1(_09585_),
    .X(_09586_));
 sky130_fd_sc_hd__mux4_1 _22427_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][6] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][6] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][6] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][6] ),
    .S0(_09423_),
    .S1(_09424_),
    .X(_09587_));
 sky130_fd_sc_hd__a21o_1 _22428_ (.A1(_09528_),
    .A2(_09587_),
    .B1(_09426_),
    .X(_09588_));
 sky130_fd_sc_hd__a21o_1 _22429_ (.A1(_09415_),
    .A2(_09586_),
    .B1(_09588_),
    .X(_09589_));
 sky130_fd_sc_hd__mux4_1 _22430_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][6] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][6] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][6] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][6] ),
    .S0(_09431_),
    .S1(_09532_),
    .X(_09590_));
 sky130_fd_sc_hd__mux4_1 _22431_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][6] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][6] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][6] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][6] ),
    .S0(_09552_),
    .S1(_09382_),
    .X(_09591_));
 sky130_fd_sc_hd__and2_1 _22432_ (.A(_09534_),
    .B(_09591_),
    .X(_09592_));
 sky130_fd_sc_hd__a211o_1 _22433_ (.A1(_09429_),
    .A2(_09590_),
    .B1(_09592_),
    .C1(_09438_),
    .X(_09593_));
 sky130_fd_sc_hd__and4_1 _22434_ (.A(_09389_),
    .B(_09584_),
    .C(_09589_),
    .D(_09593_),
    .X(_09594_));
 sky130_fd_sc_hd__clkbuf_1 _22435_ (.A(_09594_),
    .X(_01130_));
 sky130_fd_sc_hd__mux4_1 _22436_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][7] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][7] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][7] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][7] ),
    .S0(_09393_),
    .S1(_09395_),
    .X(_09595_));
 sky130_fd_sc_hd__or2_1 _22437_ (.A(_09511_),
    .B(_09595_),
    .X(_09596_));
 sky130_fd_sc_hd__mux4_1 _22438_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][7] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][7] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][7] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][7] ),
    .S0(_09446_),
    .S1(_09402_),
    .X(_09597_));
 sky130_fd_sc_hd__o21a_1 _22439_ (.A1(_09451_),
    .A2(_09597_),
    .B1(_09404_),
    .X(_09598_));
 sky130_fd_sc_hd__mux4_1 _22440_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][7] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][7] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][7] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][7] ),
    .S0(_09406_),
    .S1(_09408_),
    .X(_09599_));
 sky130_fd_sc_hd__mux4_1 _22441_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][7] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][7] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][7] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][7] ),
    .S0(_09512_),
    .S1(_09408_),
    .X(_09600_));
 sky130_fd_sc_hd__mux2_2 _22442_ (.A0(_09599_),
    .A1(_09600_),
    .S(_09380_),
    .X(_09601_));
 sky130_fd_sc_hd__a221o_1 _22443_ (.A1(_09596_),
    .A2(_09598_),
    .B1(_09601_),
    .B2(_09412_),
    .C1(_09413_),
    .X(_09602_));
 sky130_fd_sc_hd__mux4_1 _22444_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][7] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][7] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][7] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][7] ),
    .S0(_09417_),
    .S1(_09585_),
    .X(_09603_));
 sky130_fd_sc_hd__buf_4 _22445_ (.A(_09401_),
    .X(_09604_));
 sky130_fd_sc_hd__mux4_1 _22446_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][7] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][7] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][7] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][7] ),
    .S0(_09604_),
    .S1(_09424_),
    .X(_09605_));
 sky130_fd_sc_hd__a21o_1 _22447_ (.A1(_09528_),
    .A2(_09605_),
    .B1(_09426_),
    .X(_09606_));
 sky130_fd_sc_hd__a21o_1 _22448_ (.A1(_09415_),
    .A2(_09603_),
    .B1(_09606_),
    .X(_09607_));
 sky130_fd_sc_hd__clkbuf_8 _22449_ (.A(_09430_),
    .X(_09608_));
 sky130_fd_sc_hd__mux4_1 _22450_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][7] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][7] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][7] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][7] ),
    .S0(_09608_),
    .S1(_09532_),
    .X(_09609_));
 sky130_fd_sc_hd__mux4_1 _22451_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][7] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][7] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][7] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][7] ),
    .S0(_09552_),
    .S1(_09382_),
    .X(_09610_));
 sky130_fd_sc_hd__and2_1 _22452_ (.A(_09534_),
    .B(_09610_),
    .X(_09611_));
 sky130_fd_sc_hd__a211o_1 _22453_ (.A1(_09429_),
    .A2(_09609_),
    .B1(_09611_),
    .C1(_09438_),
    .X(_09612_));
 sky130_fd_sc_hd__and4_1 _22454_ (.A(_09389_),
    .B(_09602_),
    .C(_09607_),
    .D(_09612_),
    .X(_09613_));
 sky130_fd_sc_hd__clkbuf_1 _22455_ (.A(_09613_),
    .X(_01131_));
 sky130_fd_sc_hd__mux4_1 _22456_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][8] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][8] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][8] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][8] ),
    .S0(_09393_),
    .S1(_09395_),
    .X(_09614_));
 sky130_fd_sc_hd__or2_1 _22457_ (.A(_09511_),
    .B(_09614_),
    .X(_09615_));
 sky130_fd_sc_hd__mux4_1 _22458_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][8] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][8] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][8] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][8] ),
    .S0(_09446_),
    .S1(_09402_),
    .X(_09616_));
 sky130_fd_sc_hd__o21a_1 _22459_ (.A1(_09451_),
    .A2(_09616_),
    .B1(_09404_),
    .X(_09617_));
 sky130_fd_sc_hd__mux4_1 _22460_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][8] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][8] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][8] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][8] ),
    .S0(_09406_),
    .S1(_09408_),
    .X(_09618_));
 sky130_fd_sc_hd__mux4_1 _22461_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][8] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][8] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][8] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][8] ),
    .S0(_09512_),
    .S1(_09408_),
    .X(_09619_));
 sky130_fd_sc_hd__mux2_2 _22462_ (.A0(_09618_),
    .A1(_09619_),
    .S(_09380_),
    .X(_09620_));
 sky130_fd_sc_hd__a221o_1 _22463_ (.A1(_09615_),
    .A2(_09617_),
    .B1(_09620_),
    .B2(_09412_),
    .C1(_09413_),
    .X(_09621_));
 sky130_fd_sc_hd__clkbuf_4 _22464_ (.A(_09399_),
    .X(_09622_));
 sky130_fd_sc_hd__mux4_1 _22465_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][8] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][8] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][8] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][8] ),
    .S0(_09417_),
    .S1(_09585_),
    .X(_09623_));
 sky130_fd_sc_hd__mux4_1 _22466_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][8] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][8] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][8] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][8] ),
    .S0(_09604_),
    .S1(_09424_),
    .X(_09624_));
 sky130_fd_sc_hd__a21o_1 _22467_ (.A1(_09528_),
    .A2(_09624_),
    .B1(_09426_),
    .X(_09625_));
 sky130_fd_sc_hd__a21o_1 _22468_ (.A1(_09622_),
    .A2(_09623_),
    .B1(_09625_),
    .X(_09626_));
 sky130_fd_sc_hd__clkbuf_4 _22469_ (.A(_09399_),
    .X(_09627_));
 sky130_fd_sc_hd__mux4_1 _22470_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][8] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][8] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][8] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][8] ),
    .S0(_09608_),
    .S1(_09532_),
    .X(_09628_));
 sky130_fd_sc_hd__mux4_1 _22471_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][8] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][8] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][8] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][8] ),
    .S0(_09552_),
    .S1(_09382_),
    .X(_09629_));
 sky130_fd_sc_hd__and2_1 _22472_ (.A(_09534_),
    .B(_09629_),
    .X(_09630_));
 sky130_fd_sc_hd__a211o_1 _22473_ (.A1(_09627_),
    .A2(_09628_),
    .B1(_09630_),
    .C1(_09438_),
    .X(_09631_));
 sky130_fd_sc_hd__and4_1 _22474_ (.A(_09389_),
    .B(_09621_),
    .C(_09626_),
    .D(_09631_),
    .X(_09632_));
 sky130_fd_sc_hd__clkbuf_1 _22475_ (.A(_09632_),
    .X(_01132_));
 sky130_fd_sc_hd__mux4_1 _22476_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][9] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][9] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][9] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][9] ),
    .S0(_09445_),
    .S1(_09447_),
    .X(_09633_));
 sky130_fd_sc_hd__mux4_1 _22477_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][9] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][9] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][9] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][9] ),
    .S0(_09434_),
    .S1(_09558_),
    .X(_09634_));
 sky130_fd_sc_hd__mux2_2 _22478_ (.A0(_09633_),
    .A1(_09634_),
    .S(_09449_),
    .X(_09635_));
 sky130_fd_sc_hd__clkbuf_4 _22479_ (.A(_09391_),
    .X(_09636_));
 sky130_fd_sc_hd__clkbuf_8 _22480_ (.A(_09395_),
    .X(_09637_));
 sky130_fd_sc_hd__mux4_2 _22481_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][9] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][9] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][9] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][9] ),
    .S0(_09463_),
    .S1(_09637_),
    .X(_09638_));
 sky130_fd_sc_hd__nor2_1 _22482_ (.A(_09636_),
    .B(_09638_),
    .Y(_09639_));
 sky130_fd_sc_hd__mux4_1 _22483_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][9] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][9] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][9] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][9] ),
    .S0(_09558_),
    .S1(_09453_),
    .X(_09640_));
 sky130_fd_sc_hd__o21ai_1 _22484_ (.A1(_09495_),
    .A2(_09640_),
    .B1(_09457_),
    .Y(_09641_));
 sky130_fd_sc_hd__o2bb2a_1 _22485_ (.A1_N(_09442_),
    .A2_N(_09635_),
    .B1(_09639_),
    .B2(_09641_),
    .X(_09642_));
 sky130_fd_sc_hd__nor2_1 _22486_ (.A(_09441_),
    .B(_09642_),
    .Y(_09643_));
 sky130_fd_sc_hd__mux4_2 _22487_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][9] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][9] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][9] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][9] ),
    .S0(_09464_),
    .S1(_09467_),
    .X(_09644_));
 sky130_fd_sc_hd__mux4_1 _22488_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][9] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][9] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][9] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][9] ),
    .S0(_09418_),
    .S1(_09485_),
    .X(_09645_));
 sky130_fd_sc_hd__or2_1 _22489_ (.A(_09469_),
    .B(_09645_),
    .X(_09646_));
 sky130_fd_sc_hd__o211a_1 _22490_ (.A1(_09461_),
    .A2(_09644_),
    .B1(_09646_),
    .C1(_09489_),
    .X(_09647_));
 sky130_fd_sc_hd__mux4_1 _22491_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][9] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][9] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][9] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][9] ),
    .S0(_09478_),
    .S1(_09479_),
    .X(_09648_));
 sky130_fd_sc_hd__mux4_1 _22492_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][9] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][9] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][9] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][9] ),
    .S0(_09477_),
    .S1(_09383_),
    .X(_09649_));
 sky130_fd_sc_hd__or2_1 _22493_ (.A(_09482_),
    .B(_09649_),
    .X(_09650_));
 sky130_fd_sc_hd__o211a_1 _22494_ (.A1(_09476_),
    .A2(_09648_),
    .B1(_09650_),
    .C1(_09474_),
    .X(_09651_));
 sky130_fd_sc_hd__o31a_1 _22495_ (.A1(_09643_),
    .A2(_09647_),
    .A3(_09651_),
    .B1(_09491_),
    .X(_01133_));
 sky130_fd_sc_hd__mux4_2 _22496_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][10] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][10] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][10] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][10] ),
    .S0(_09385_),
    .S1(_09637_),
    .X(_09652_));
 sky130_fd_sc_hd__nor2_1 _22497_ (.A(_09422_),
    .B(_09652_),
    .Y(_09653_));
 sky130_fd_sc_hd__mux4_2 _22498_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][10] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][10] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][10] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][10] ),
    .S0(_09385_),
    .S1(_09637_),
    .X(_09654_));
 sky130_fd_sc_hd__nor2_1 _22499_ (.A(_09495_),
    .B(_09654_),
    .Y(_09655_));
 sky130_fd_sc_hd__buf_4 _22500_ (.A(_09385_),
    .X(_09656_));
 sky130_fd_sc_hd__mux4_1 _22501_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][10] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][10] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][10] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][10] ),
    .S0(_09483_),
    .S1(_09656_),
    .X(_09657_));
 sky130_fd_sc_hd__nor2_1 _22502_ (.A(_09452_),
    .B(_09657_),
    .Y(_09658_));
 sky130_fd_sc_hd__mux4_1 _22503_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][10] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][10] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][10] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][10] ),
    .S0(_09385_),
    .S1(_09637_),
    .X(_09659_));
 sky130_fd_sc_hd__o21ai_1 _22504_ (.A1(_09469_),
    .A2(_09659_),
    .B1(_09457_),
    .Y(_09660_));
 sky130_fd_sc_hd__o32a_1 _22505_ (.A1(_09457_),
    .A2(_09653_),
    .A3(_09655_),
    .B1(_09658_),
    .B2(_09660_),
    .X(_09661_));
 sky130_fd_sc_hd__nor2_1 _22506_ (.A(_09441_),
    .B(_09661_),
    .Y(_09662_));
 sky130_fd_sc_hd__mux4_2 _22507_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][10] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][10] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][10] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][10] ),
    .S0(_09386_),
    .S1(_09467_),
    .X(_09663_));
 sky130_fd_sc_hd__mux4_1 _22508_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][10] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][10] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][10] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][10] ),
    .S0(_09418_),
    .S1(_09485_),
    .X(_09664_));
 sky130_fd_sc_hd__or2_1 _22509_ (.A(_09469_),
    .B(_09664_),
    .X(_09665_));
 sky130_fd_sc_hd__o211a_1 _22510_ (.A1(_09461_),
    .A2(_09663_),
    .B1(_09665_),
    .C1(_09489_),
    .X(_09666_));
 sky130_fd_sc_hd__mux4_1 _22511_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][10] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][10] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][10] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][10] ),
    .S0(_09478_),
    .S1(_09479_),
    .X(_09667_));
 sky130_fd_sc_hd__mux4_1 _22512_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][10] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][10] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][10] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][10] ),
    .S0(_09477_),
    .S1(_09466_),
    .X(_09668_));
 sky130_fd_sc_hd__or2_1 _22513_ (.A(_09482_),
    .B(_09668_),
    .X(_09669_));
 sky130_fd_sc_hd__o211a_1 _22514_ (.A1(_09476_),
    .A2(_09667_),
    .B1(_09669_),
    .C1(_09474_),
    .X(_09670_));
 sky130_fd_sc_hd__o31a_1 _22515_ (.A1(_09662_),
    .A2(_09666_),
    .A3(_09670_),
    .B1(_09491_),
    .X(_01134_));
 sky130_fd_sc_hd__mux4_1 _22516_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][11] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][11] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][11] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][11] ),
    .S0(_09445_),
    .S1(_09447_),
    .X(_09671_));
 sky130_fd_sc_hd__mux4_1 _22517_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][11] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][11] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][11] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][11] ),
    .S0(_09434_),
    .S1(_09558_),
    .X(_09672_));
 sky130_fd_sc_hd__mux2_1 _22518_ (.A0(_09671_),
    .A1(_09672_),
    .S(_09449_),
    .X(_09673_));
 sky130_fd_sc_hd__mux4_1 _22519_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][11] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][11] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][11] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][11] ),
    .S0(_09463_),
    .S1(_09637_),
    .X(_09674_));
 sky130_fd_sc_hd__nor2_1 _22520_ (.A(_09636_),
    .B(_09674_),
    .Y(_09675_));
 sky130_fd_sc_hd__mux4_1 _22521_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][11] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][11] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][11] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][11] ),
    .S0(_09558_),
    .S1(_09417_),
    .X(_09676_));
 sky130_fd_sc_hd__o21ai_1 _22522_ (.A1(_09495_),
    .A2(_09676_),
    .B1(_09472_),
    .Y(_09677_));
 sky130_fd_sc_hd__o2bb2a_1 _22523_ (.A1_N(_09442_),
    .A2_N(_09673_),
    .B1(_09675_),
    .B2(_09677_),
    .X(_09678_));
 sky130_fd_sc_hd__nor2_1 _22524_ (.A(_09441_),
    .B(_09678_),
    .Y(_09679_));
 sky130_fd_sc_hd__mux4_1 _22525_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][11] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][11] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][11] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][11] ),
    .S0(_09386_),
    .S1(_09419_),
    .X(_09680_));
 sky130_fd_sc_hd__mux4_1 _22526_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][11] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][11] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][11] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][11] ),
    .S0(_09463_),
    .S1(_09466_),
    .X(_09681_));
 sky130_fd_sc_hd__or2_1 _22527_ (.A(_09636_),
    .B(_09681_),
    .X(_09682_));
 sky130_fd_sc_hd__o211a_1 _22528_ (.A1(_09461_),
    .A2(_09680_),
    .B1(_09682_),
    .C1(_09474_),
    .X(_09683_));
 sky130_fd_sc_hd__mux4_2 _22529_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][11] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][11] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][11] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][11] ),
    .S0(_09478_),
    .S1(_09479_),
    .X(_09684_));
 sky130_fd_sc_hd__mux4_1 _22530_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][11] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][11] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][11] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][11] ),
    .S0(_09424_),
    .S1(_09485_),
    .X(_09685_));
 sky130_fd_sc_hd__or2_1 _22531_ (.A(_09482_),
    .B(_09685_),
    .X(_09686_));
 sky130_fd_sc_hd__o211a_1 _22532_ (.A1(_09476_),
    .A2(_09684_),
    .B1(_09686_),
    .C1(_09489_),
    .X(_09687_));
 sky130_fd_sc_hd__o31a_1 _22533_ (.A1(_09679_),
    .A2(_09683_),
    .A3(_09687_),
    .B1(_09491_),
    .X(_01135_));
 sky130_fd_sc_hd__mux4_1 _22534_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][12] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][12] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][12] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][12] ),
    .S0(_09384_),
    .S1(_09577_),
    .X(_09688_));
 sky130_fd_sc_hd__mux4_1 _22535_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][12] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][12] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][12] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][12] ),
    .S0(_09384_),
    .S1(_09430_),
    .X(_09689_));
 sky130_fd_sc_hd__mux2_2 _22536_ (.A0(_09688_),
    .A1(_09689_),
    .S(_09421_),
    .X(_09690_));
 sky130_fd_sc_hd__mux4_1 _22537_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][12] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][12] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][12] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][12] ),
    .S0(_09393_),
    .S1(_09465_),
    .X(_09691_));
 sky130_fd_sc_hd__or2_1 _22538_ (.A(_09391_),
    .B(_09691_),
    .X(_09692_));
 sky130_fd_sc_hd__mux4_1 _22539_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][12] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][12] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][12] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][12] ),
    .S0(_09400_),
    .S1(_09484_),
    .X(_09693_));
 sky130_fd_sc_hd__o21a_1 _22540_ (.A1(_09399_),
    .A2(_09693_),
    .B1(_09472_),
    .X(_09694_));
 sky130_fd_sc_hd__a221o_1 _22541_ (.A1(_09412_),
    .A2(_09690_),
    .B1(_09692_),
    .B2(_09694_),
    .C1(_09413_),
    .X(_09695_));
 sky130_fd_sc_hd__mux4_1 _22542_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][12] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][12] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][12] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][12] ),
    .S0(_09417_),
    .S1(_09585_),
    .X(_09696_));
 sky130_fd_sc_hd__mux4_1 _22543_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][12] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][12] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][12] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][12] ),
    .S0(_09604_),
    .S1(_09424_),
    .X(_09697_));
 sky130_fd_sc_hd__a21o_1 _22544_ (.A1(_09528_),
    .A2(_09697_),
    .B1(_09426_),
    .X(_09698_));
 sky130_fd_sc_hd__a21o_1 _22545_ (.A1(_09622_),
    .A2(_09696_),
    .B1(_09698_),
    .X(_09699_));
 sky130_fd_sc_hd__mux4_1 _22546_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][12] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][12] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][12] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][12] ),
    .S0(_09608_),
    .S1(_09532_),
    .X(_09700_));
 sky130_fd_sc_hd__mux4_1 _22547_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][12] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][12] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][12] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][12] ),
    .S0(_09552_),
    .S1(_09382_),
    .X(_09701_));
 sky130_fd_sc_hd__and2_1 _22548_ (.A(_09534_),
    .B(_09701_),
    .X(_09702_));
 sky130_fd_sc_hd__a211o_1 _22549_ (.A1(_09627_),
    .A2(_09700_),
    .B1(_09702_),
    .C1(_09438_),
    .X(_09703_));
 sky130_fd_sc_hd__and4_1 _22550_ (.A(_09389_),
    .B(_09695_),
    .C(_09699_),
    .D(_09703_),
    .X(_09704_));
 sky130_fd_sc_hd__clkbuf_1 _22551_ (.A(_09704_),
    .X(_01136_));
 sky130_fd_sc_hd__buf_2 _22552_ (.A(_09388_),
    .X(_09705_));
 sky130_fd_sc_hd__mux4_1 _22553_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][13] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][13] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][13] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][13] ),
    .S0(_09384_),
    .S1(_09577_),
    .X(_09706_));
 sky130_fd_sc_hd__mux4_1 _22554_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][13] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][13] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][13] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][13] ),
    .S0(_09401_),
    .S1(_09430_),
    .X(_09707_));
 sky130_fd_sc_hd__mux2_1 _22555_ (.A0(_09706_),
    .A1(_09707_),
    .S(_09421_),
    .X(_09708_));
 sky130_fd_sc_hd__mux4_1 _22556_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][13] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][13] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][13] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][13] ),
    .S0(_09393_),
    .S1(_09465_),
    .X(_09709_));
 sky130_fd_sc_hd__or2_1 _22557_ (.A(_09391_),
    .B(_09709_),
    .X(_09710_));
 sky130_fd_sc_hd__mux4_1 _22558_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][13] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][13] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][13] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][13] ),
    .S0(_09400_),
    .S1(_09484_),
    .X(_09711_));
 sky130_fd_sc_hd__o21a_1 _22559_ (.A1(_09399_),
    .A2(_09711_),
    .B1(_09472_),
    .X(_09712_));
 sky130_fd_sc_hd__a221o_1 _22560_ (.A1(_09412_),
    .A2(_09708_),
    .B1(_09710_),
    .B2(_09712_),
    .C1(_09413_),
    .X(_09713_));
 sky130_fd_sc_hd__buf_4 _22561_ (.A(_09416_),
    .X(_09714_));
 sky130_fd_sc_hd__mux4_1 _22562_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][13] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][13] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][13] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][13] ),
    .S0(_09714_),
    .S1(_09585_),
    .X(_09715_));
 sky130_fd_sc_hd__buf_4 _22563_ (.A(_09400_),
    .X(_09716_));
 sky130_fd_sc_hd__mux4_1 _22564_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][13] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][13] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][13] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][13] ),
    .S0(_09604_),
    .S1(_09716_),
    .X(_09717_));
 sky130_fd_sc_hd__a21o_1 _22565_ (.A1(_09528_),
    .A2(_09717_),
    .B1(_09426_),
    .X(_09718_));
 sky130_fd_sc_hd__a21o_1 _22566_ (.A1(_09622_),
    .A2(_09715_),
    .B1(_09718_),
    .X(_09719_));
 sky130_fd_sc_hd__mux4_1 _22567_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][13] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][13] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][13] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][13] ),
    .S0(_09608_),
    .S1(_09532_),
    .X(_09720_));
 sky130_fd_sc_hd__buf_4 _22568_ (.A(_09381_),
    .X(_09721_));
 sky130_fd_sc_hd__mux4_1 _22569_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][13] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][13] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][13] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][13] ),
    .S0(_09552_),
    .S1(_09721_),
    .X(_09722_));
 sky130_fd_sc_hd__and2_1 _22570_ (.A(_09534_),
    .B(_09722_),
    .X(_09723_));
 sky130_fd_sc_hd__a211o_1 _22571_ (.A1(_09627_),
    .A2(_09720_),
    .B1(_09723_),
    .C1(_09438_),
    .X(_09724_));
 sky130_fd_sc_hd__and4_1 _22572_ (.A(_09705_),
    .B(_09713_),
    .C(_09719_),
    .D(_09724_),
    .X(_09725_));
 sky130_fd_sc_hd__clkbuf_1 _22573_ (.A(_09725_),
    .X(_01137_));
 sky130_fd_sc_hd__mux4_1 _22574_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][14] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][14] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][14] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][14] ),
    .S0(_09445_),
    .S1(_09447_),
    .X(_09726_));
 sky130_fd_sc_hd__mux4_1 _22575_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][14] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][14] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][14] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][14] ),
    .S0(_09434_),
    .S1(_09558_),
    .X(_09727_));
 sky130_fd_sc_hd__mux2_1 _22576_ (.A0(_09726_),
    .A1(_09727_),
    .S(_09449_),
    .X(_09728_));
 sky130_fd_sc_hd__mux4_1 _22577_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][14] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][14] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][14] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][14] ),
    .S0(_09443_),
    .S1(_09453_),
    .X(_09729_));
 sky130_fd_sc_hd__nor2_1 _22578_ (.A(_09495_),
    .B(_09729_),
    .Y(_09730_));
 sky130_fd_sc_hd__mux4_1 _22579_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][14] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][14] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][14] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][14] ),
    .S0(_09484_),
    .S1(_09431_),
    .X(_09731_));
 sky130_fd_sc_hd__o21ai_1 _22580_ (.A1(_09422_),
    .A2(_09731_),
    .B1(_09472_),
    .Y(_09732_));
 sky130_fd_sc_hd__o2bb2a_1 _22581_ (.A1_N(_09442_),
    .A2_N(_09728_),
    .B1(_09730_),
    .B2(_09732_),
    .X(_09733_));
 sky130_fd_sc_hd__nor2_1 _22582_ (.A(_09441_),
    .B(_09733_),
    .Y(_09734_));
 sky130_fd_sc_hd__mux4_2 _22583_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][14] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][14] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][14] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][14] ),
    .S0(_09386_),
    .S1(_09419_),
    .X(_09735_));
 sky130_fd_sc_hd__mux4_2 _22584_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][14] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][14] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][14] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][14] ),
    .S0(_09418_),
    .S1(_09485_),
    .X(_09736_));
 sky130_fd_sc_hd__or2_1 _22585_ (.A(_09636_),
    .B(_09736_),
    .X(_09737_));
 sky130_fd_sc_hd__o211a_1 _22586_ (.A1(_09461_),
    .A2(_09735_),
    .B1(_09737_),
    .C1(_09489_),
    .X(_09738_));
 sky130_fd_sc_hd__mux4_1 _22587_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][14] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][14] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][14] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][14] ),
    .S0(_09464_),
    .S1(_09479_),
    .X(_09739_));
 sky130_fd_sc_hd__mux4_1 _22588_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][14] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][14] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][14] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][14] ),
    .S0(_09477_),
    .S1(_09466_),
    .X(_09740_));
 sky130_fd_sc_hd__or2_1 _22589_ (.A(_09482_),
    .B(_09740_),
    .X(_09741_));
 sky130_fd_sc_hd__o211a_1 _22590_ (.A1(_09476_),
    .A2(_09739_),
    .B1(_09741_),
    .C1(_09474_),
    .X(_09742_));
 sky130_fd_sc_hd__o31a_1 _22591_ (.A1(_09734_),
    .A2(_09738_),
    .A3(_09742_),
    .B1(_09491_),
    .X(_01138_));
 sky130_fd_sc_hd__mux4_1 _22592_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][15] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][15] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][15] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][15] ),
    .S0(_09384_),
    .S1(_09430_),
    .X(_09743_));
 sky130_fd_sc_hd__mux4_1 _22593_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][15] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][15] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][15] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][15] ),
    .S0(_09401_),
    .S1(_09430_),
    .X(_09744_));
 sky130_fd_sc_hd__mux2_1 _22594_ (.A0(_09743_),
    .A1(_09744_),
    .S(_09421_),
    .X(_09745_));
 sky130_fd_sc_hd__mux4_1 _22595_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][15] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][15] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][15] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][15] ),
    .S0(_09393_),
    .S1(_09465_),
    .X(_09746_));
 sky130_fd_sc_hd__or2_1 _22596_ (.A(_09391_),
    .B(_09746_),
    .X(_09747_));
 sky130_fd_sc_hd__mux4_1 _22597_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][15] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][15] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][15] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][15] ),
    .S0(_09400_),
    .S1(_09484_),
    .X(_09748_));
 sky130_fd_sc_hd__o21a_1 _22598_ (.A1(_09399_),
    .A2(_09748_),
    .B1(_09472_),
    .X(_09749_));
 sky130_fd_sc_hd__a221o_1 _22599_ (.A1(_09412_),
    .A2(_09745_),
    .B1(_09747_),
    .B2(_09749_),
    .C1(_09413_),
    .X(_09750_));
 sky130_fd_sc_hd__mux4_1 _22600_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][15] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][15] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][15] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][15] ),
    .S0(_09714_),
    .S1(_09585_),
    .X(_09751_));
 sky130_fd_sc_hd__mux4_1 _22601_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][15] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][15] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][15] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][15] ),
    .S0(_09604_),
    .S1(_09716_),
    .X(_09752_));
 sky130_fd_sc_hd__a21o_1 _22602_ (.A1(_09528_),
    .A2(_09752_),
    .B1(_09426_),
    .X(_09753_));
 sky130_fd_sc_hd__a21o_1 _22603_ (.A1(_09622_),
    .A2(_09751_),
    .B1(_09753_),
    .X(_09754_));
 sky130_fd_sc_hd__mux4_1 _22604_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][15] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][15] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][15] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][15] ),
    .S0(_09608_),
    .S1(_09532_),
    .X(_09755_));
 sky130_fd_sc_hd__mux4_1 _22605_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][15] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][15] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][15] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][15] ),
    .S0(_09552_),
    .S1(_09721_),
    .X(_09756_));
 sky130_fd_sc_hd__and2_1 _22606_ (.A(_09534_),
    .B(_09756_),
    .X(_09757_));
 sky130_fd_sc_hd__a211o_1 _22607_ (.A1(_09627_),
    .A2(_09755_),
    .B1(_09757_),
    .C1(_09438_),
    .X(_09758_));
 sky130_fd_sc_hd__and4_1 _22608_ (.A(_09705_),
    .B(_09750_),
    .C(_09754_),
    .D(_09758_),
    .X(_09759_));
 sky130_fd_sc_hd__clkbuf_1 _22609_ (.A(_09759_),
    .X(_01139_));
 sky130_fd_sc_hd__mux4_1 _22610_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][16] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][16] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][16] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][16] ),
    .S0(_09512_),
    .S1(_09513_),
    .X(_09760_));
 sky130_fd_sc_hd__or2_1 _22611_ (.A(_09511_),
    .B(_09760_),
    .X(_09761_));
 sky130_fd_sc_hd__mux4_2 _22612_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][16] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][16] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][16] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][16] ),
    .S0(_09517_),
    .S1(_09577_),
    .X(_09762_));
 sky130_fd_sc_hd__or2_1 _22613_ (.A(_09516_),
    .B(_09762_),
    .X(_09763_));
 sky130_fd_sc_hd__mux4_1 _22614_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][16] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][16] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][16] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][16] ),
    .S0(_09446_),
    .S1(_09402_),
    .X(_09764_));
 sky130_fd_sc_hd__mux4_1 _22615_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][16] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][16] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][16] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][16] ),
    .S0(_09392_),
    .S1(_09394_),
    .X(_09765_));
 sky130_fd_sc_hd__or2_1 _22616_ (.A(_09390_),
    .B(_09765_),
    .X(_09766_));
 sky130_fd_sc_hd__o211a_1 _22617_ (.A1(_09451_),
    .A2(_09764_),
    .B1(_09766_),
    .C1(_09523_),
    .X(_09767_));
 sky130_fd_sc_hd__a311o_2 _22618_ (.A1(_09510_),
    .A2(_09761_),
    .A3(_09763_),
    .B1(_09767_),
    .C1(_09525_),
    .X(_09768_));
 sky130_fd_sc_hd__mux4_1 _22619_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][16] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][16] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][16] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][16] ),
    .S0(_09714_),
    .S1(_09585_),
    .X(_09769_));
 sky130_fd_sc_hd__mux4_1 _22620_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][16] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][16] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][16] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][16] ),
    .S0(_09604_),
    .S1(_09716_),
    .X(_09770_));
 sky130_fd_sc_hd__a21o_1 _22621_ (.A1(_09528_),
    .A2(_09770_),
    .B1(_09426_),
    .X(_09771_));
 sky130_fd_sc_hd__a21o_1 _22622_ (.A1(_09622_),
    .A2(_09769_),
    .B1(_09771_),
    .X(_09772_));
 sky130_fd_sc_hd__mux4_1 _22623_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][16] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][16] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][16] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][16] ),
    .S0(_09608_),
    .S1(_09532_),
    .X(_09773_));
 sky130_fd_sc_hd__mux4_1 _22624_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][16] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][16] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][16] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][16] ),
    .S0(_09552_),
    .S1(_09721_),
    .X(_09774_));
 sky130_fd_sc_hd__and2_1 _22625_ (.A(_09534_),
    .B(_09774_),
    .X(_09775_));
 sky130_fd_sc_hd__a211o_1 _22626_ (.A1(_09627_),
    .A2(_09773_),
    .B1(_09775_),
    .C1(_09438_),
    .X(_09776_));
 sky130_fd_sc_hd__and4_1 _22627_ (.A(_09705_),
    .B(_09768_),
    .C(_09772_),
    .D(_09776_),
    .X(_09777_));
 sky130_fd_sc_hd__clkbuf_1 _22628_ (.A(_09777_),
    .X(_01140_));
 sky130_fd_sc_hd__mux4_2 _22629_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][17] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][17] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][17] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][17] ),
    .S0(_09512_),
    .S1(_09513_),
    .X(_09778_));
 sky130_fd_sc_hd__or2_1 _22630_ (.A(_09511_),
    .B(_09778_),
    .X(_09779_));
 sky130_fd_sc_hd__mux4_2 _22631_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][17] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][17] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][17] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][17] ),
    .S0(_09517_),
    .S1(_09577_),
    .X(_09780_));
 sky130_fd_sc_hd__or2_1 _22632_ (.A(_09516_),
    .B(_09780_),
    .X(_09781_));
 sky130_fd_sc_hd__mux4_1 _22633_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][17] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][17] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][17] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][17] ),
    .S0(_09446_),
    .S1(_09402_),
    .X(_09782_));
 sky130_fd_sc_hd__mux4_1 _22634_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][17] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][17] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][17] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][17] ),
    .S0(_09392_),
    .S1(_09394_),
    .X(_09783_));
 sky130_fd_sc_hd__or2_1 _22635_ (.A(_09390_),
    .B(_09783_),
    .X(_09784_));
 sky130_fd_sc_hd__o211a_1 _22636_ (.A1(_09451_),
    .A2(_09782_),
    .B1(_09784_),
    .C1(_09523_),
    .X(_09785_));
 sky130_fd_sc_hd__a311o_1 _22637_ (.A1(_09510_),
    .A2(_09779_),
    .A3(_09781_),
    .B1(_09785_),
    .C1(_09525_),
    .X(_09786_));
 sky130_fd_sc_hd__mux4_1 _22638_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][17] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][17] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][17] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][17] ),
    .S0(_09714_),
    .S1(_09585_),
    .X(_09787_));
 sky130_fd_sc_hd__mux4_1 _22639_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][17] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][17] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][17] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][17] ),
    .S0(_09604_),
    .S1(_09716_),
    .X(_09788_));
 sky130_fd_sc_hd__clkbuf_4 _22640_ (.A(_09387_),
    .X(_09789_));
 sky130_fd_sc_hd__a21o_1 _22641_ (.A1(_09528_),
    .A2(_09788_),
    .B1(_09789_),
    .X(_09790_));
 sky130_fd_sc_hd__a21o_1 _22642_ (.A1(_09622_),
    .A2(_09787_),
    .B1(_09790_),
    .X(_09791_));
 sky130_fd_sc_hd__mux4_1 _22643_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][17] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][17] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][17] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][17] ),
    .S0(_09608_),
    .S1(_09532_),
    .X(_09792_));
 sky130_fd_sc_hd__mux4_1 _22644_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][17] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][17] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][17] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][17] ),
    .S0(_09552_),
    .S1(_09721_),
    .X(_09793_));
 sky130_fd_sc_hd__and2_1 _22645_ (.A(_09534_),
    .B(_09793_),
    .X(_09794_));
 sky130_fd_sc_hd__clkbuf_4 _22646_ (.A(_09437_),
    .X(_09795_));
 sky130_fd_sc_hd__a211o_1 _22647_ (.A1(_09627_),
    .A2(_09792_),
    .B1(_09794_),
    .C1(_09795_),
    .X(_09796_));
 sky130_fd_sc_hd__and4_1 _22648_ (.A(_09705_),
    .B(_09786_),
    .C(_09791_),
    .D(_09796_),
    .X(_09797_));
 sky130_fd_sc_hd__clkbuf_1 _22649_ (.A(_09797_),
    .X(_01141_));
 sky130_fd_sc_hd__mux4_1 _22650_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][18] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][18] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][18] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][18] ),
    .S0(_09384_),
    .S1(_09430_),
    .X(_09798_));
 sky130_fd_sc_hd__mux4_1 _22651_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][18] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][18] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][18] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][18] ),
    .S0(_09401_),
    .S1(_09430_),
    .X(_09799_));
 sky130_fd_sc_hd__mux2_2 _22652_ (.A0(_09798_),
    .A1(_09799_),
    .S(_09421_),
    .X(_09800_));
 sky130_fd_sc_hd__mux4_1 _22653_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][18] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][18] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][18] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][18] ),
    .S0(_09393_),
    .S1(_09465_),
    .X(_09801_));
 sky130_fd_sc_hd__or2_1 _22654_ (.A(_09391_),
    .B(_09801_),
    .X(_09802_));
 sky130_fd_sc_hd__mux4_1 _22655_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][18] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][18] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][18] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][18] ),
    .S0(_09400_),
    .S1(_09484_),
    .X(_09803_));
 sky130_fd_sc_hd__o21a_1 _22656_ (.A1(_09399_),
    .A2(_09803_),
    .B1(_09523_),
    .X(_09804_));
 sky130_fd_sc_hd__a221o_1 _22657_ (.A1(_09412_),
    .A2(_09800_),
    .B1(_09802_),
    .B2(_09804_),
    .C1(_09413_),
    .X(_09805_));
 sky130_fd_sc_hd__mux4_1 _22658_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][18] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][18] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][18] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][18] ),
    .S0(_09714_),
    .S1(_09585_),
    .X(_09806_));
 sky130_fd_sc_hd__mux4_1 _22659_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][18] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][18] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][18] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][18] ),
    .S0(_09604_),
    .S1(_09716_),
    .X(_09807_));
 sky130_fd_sc_hd__a21o_1 _22660_ (.A1(_09433_),
    .A2(_09807_),
    .B1(_09789_),
    .X(_09808_));
 sky130_fd_sc_hd__a21o_1 _22661_ (.A1(_09622_),
    .A2(_09806_),
    .B1(_09808_),
    .X(_09809_));
 sky130_fd_sc_hd__mux4_1 _22662_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][18] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][18] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][18] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][18] ),
    .S0(_09608_),
    .S1(_09656_),
    .X(_09810_));
 sky130_fd_sc_hd__mux4_1 _22663_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][18] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][18] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][18] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][18] ),
    .S0(_09552_),
    .S1(_09721_),
    .X(_09811_));
 sky130_fd_sc_hd__and2_1 _22664_ (.A(_09481_),
    .B(_09811_),
    .X(_09812_));
 sky130_fd_sc_hd__a211o_1 _22665_ (.A1(_09627_),
    .A2(_09810_),
    .B1(_09812_),
    .C1(_09795_),
    .X(_09813_));
 sky130_fd_sc_hd__and4_1 _22666_ (.A(_09705_),
    .B(_09805_),
    .C(_09809_),
    .D(_09813_),
    .X(_09814_));
 sky130_fd_sc_hd__clkbuf_1 _22667_ (.A(_09814_),
    .X(_01142_));
 sky130_fd_sc_hd__mux4_1 _22668_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][19] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][19] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][19] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][19] ),
    .S0(_09384_),
    .S1(_09430_),
    .X(_09815_));
 sky130_fd_sc_hd__mux4_1 _22669_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][19] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][19] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][19] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][19] ),
    .S0(_09401_),
    .S1(_09430_),
    .X(_09816_));
 sky130_fd_sc_hd__mux2_1 _22670_ (.A0(_09815_),
    .A1(_09816_),
    .S(_09421_),
    .X(_09817_));
 sky130_fd_sc_hd__mux4_1 _22671_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][19] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][19] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][19] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][19] ),
    .S0(_09393_),
    .S1(_09465_),
    .X(_09818_));
 sky130_fd_sc_hd__or2_1 _22672_ (.A(_09391_),
    .B(_09818_),
    .X(_09819_));
 sky130_fd_sc_hd__mux4_1 _22673_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][19] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][19] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][19] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][19] ),
    .S0(_09400_),
    .S1(_09484_),
    .X(_09820_));
 sky130_fd_sc_hd__o21a_1 _22674_ (.A1(_09399_),
    .A2(_09820_),
    .B1(_09523_),
    .X(_09821_));
 sky130_fd_sc_hd__a221o_1 _22675_ (.A1(_09412_),
    .A2(_09817_),
    .B1(_09819_),
    .B2(_09821_),
    .C1(_09525_),
    .X(_09822_));
 sky130_fd_sc_hd__mux4_1 _22676_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][19] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][19] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][19] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][19] ),
    .S0(_09714_),
    .S1(_09585_),
    .X(_09823_));
 sky130_fd_sc_hd__mux4_1 _22677_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][19] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][19] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][19] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][19] ),
    .S0(_09604_),
    .S1(_09716_),
    .X(_09824_));
 sky130_fd_sc_hd__a21o_1 _22678_ (.A1(_09433_),
    .A2(_09824_),
    .B1(_09789_),
    .X(_09825_));
 sky130_fd_sc_hd__a21o_1 _22679_ (.A1(_09622_),
    .A2(_09823_),
    .B1(_09825_),
    .X(_09826_));
 sky130_fd_sc_hd__mux4_1 _22680_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][19] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][19] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][19] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][19] ),
    .S0(_09608_),
    .S1(_09656_),
    .X(_09827_));
 sky130_fd_sc_hd__mux4_1 _22681_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][19] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][19] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][19] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][19] ),
    .S0(_09462_),
    .S1(_09721_),
    .X(_09828_));
 sky130_fd_sc_hd__and2_1 _22682_ (.A(_09481_),
    .B(_09828_),
    .X(_09829_));
 sky130_fd_sc_hd__a211o_1 _22683_ (.A1(_09627_),
    .A2(_09827_),
    .B1(_09829_),
    .C1(_09795_),
    .X(_09830_));
 sky130_fd_sc_hd__and4_1 _22684_ (.A(_09705_),
    .B(_09822_),
    .C(_09826_),
    .D(_09830_),
    .X(_09831_));
 sky130_fd_sc_hd__clkbuf_1 _22685_ (.A(_09831_),
    .X(_01143_));
 sky130_fd_sc_hd__mux4_1 _22686_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][20] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][20] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][20] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][20] ),
    .S0(_09512_),
    .S1(_09513_),
    .X(_09832_));
 sky130_fd_sc_hd__or2_1 _22687_ (.A(_09511_),
    .B(_09832_),
    .X(_09833_));
 sky130_fd_sc_hd__mux4_2 _22688_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][20] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][20] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][20] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][20] ),
    .S0(_09517_),
    .S1(_09577_),
    .X(_09834_));
 sky130_fd_sc_hd__or2_1 _22689_ (.A(_09398_),
    .B(_09834_),
    .X(_09835_));
 sky130_fd_sc_hd__mux4_1 _22690_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][20] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][20] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][20] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][20] ),
    .S0(_09381_),
    .S1(_09423_),
    .X(_09836_));
 sky130_fd_sc_hd__mux4_1 _22691_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][20] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][20] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][20] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][20] ),
    .S0(_09392_),
    .S1(_09394_),
    .X(_09837_));
 sky130_fd_sc_hd__or2_1 _22692_ (.A(_09390_),
    .B(_09837_),
    .X(_09838_));
 sky130_fd_sc_hd__o211a_1 _22693_ (.A1(_09516_),
    .A2(_09836_),
    .B1(_09838_),
    .C1(_09523_),
    .X(_09839_));
 sky130_fd_sc_hd__a311o_1 _22694_ (.A1(_09510_),
    .A2(_09833_),
    .A3(_09835_),
    .B1(_09839_),
    .C1(_09525_),
    .X(_09840_));
 sky130_fd_sc_hd__mux4_1 _22695_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][20] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][20] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][20] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][20] ),
    .S0(_09714_),
    .S1(_09383_),
    .X(_09841_));
 sky130_fd_sc_hd__mux4_1 _22696_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][20] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][20] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][20] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][20] ),
    .S0(_09604_),
    .S1(_09716_),
    .X(_09842_));
 sky130_fd_sc_hd__a21o_1 _22697_ (.A1(_09433_),
    .A2(_09842_),
    .B1(_09789_),
    .X(_09843_));
 sky130_fd_sc_hd__a21o_1 _22698_ (.A1(_09622_),
    .A2(_09841_),
    .B1(_09843_),
    .X(_09844_));
 sky130_fd_sc_hd__mux4_1 _22699_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][20] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][20] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][20] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][20] ),
    .S0(_09608_),
    .S1(_09656_),
    .X(_09845_));
 sky130_fd_sc_hd__mux4_1 _22700_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][20] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][20] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][20] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][20] ),
    .S0(_09462_),
    .S1(_09721_),
    .X(_09846_));
 sky130_fd_sc_hd__and2_1 _22701_ (.A(_09481_),
    .B(_09846_),
    .X(_09847_));
 sky130_fd_sc_hd__a211o_1 _22702_ (.A1(_09627_),
    .A2(_09845_),
    .B1(_09847_),
    .C1(_09795_),
    .X(_09848_));
 sky130_fd_sc_hd__and4_1 _22703_ (.A(_09705_),
    .B(_09840_),
    .C(_09844_),
    .D(_09848_),
    .X(_09849_));
 sky130_fd_sc_hd__clkbuf_1 _22704_ (.A(_09849_),
    .X(_01144_));
 sky130_fd_sc_hd__mux4_1 _22705_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][21] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][21] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][21] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][21] ),
    .S0(_09445_),
    .S1(_09447_),
    .X(_09850_));
 sky130_fd_sc_hd__mux4_1 _22706_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][21] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][21] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][21] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][21] ),
    .S0(_09434_),
    .S1(_09558_),
    .X(_09851_));
 sky130_fd_sc_hd__mux2_1 _22707_ (.A0(_09850_),
    .A1(_09851_),
    .S(_09449_),
    .X(_09852_));
 sky130_fd_sc_hd__mux4_1 _22708_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][21] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][21] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][21] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][21] ),
    .S0(_09443_),
    .S1(_09453_),
    .X(_09853_));
 sky130_fd_sc_hd__nor2_1 _22709_ (.A(_09495_),
    .B(_09853_),
    .Y(_09854_));
 sky130_fd_sc_hd__mux4_1 _22710_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][21] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][21] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][21] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][21] ),
    .S0(_09484_),
    .S1(_09431_),
    .X(_09855_));
 sky130_fd_sc_hd__o21ai_1 _22711_ (.A1(_09422_),
    .A2(_09855_),
    .B1(_09472_),
    .Y(_09856_));
 sky130_fd_sc_hd__o2bb2a_1 _22712_ (.A1_N(_09442_),
    .A2_N(_09852_),
    .B1(_09854_),
    .B2(_09856_),
    .X(_09857_));
 sky130_fd_sc_hd__nor2_1 _22713_ (.A(_09441_),
    .B(_09857_),
    .Y(_09858_));
 sky130_fd_sc_hd__mux4_1 _22714_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][21] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][21] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][21] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][21] ),
    .S0(_09386_),
    .S1(_09419_),
    .X(_09859_));
 sky130_fd_sc_hd__mux4_1 _22715_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][21] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][21] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][21] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][21] ),
    .S0(_09418_),
    .S1(_09485_),
    .X(_09860_));
 sky130_fd_sc_hd__or2_1 _22716_ (.A(_09636_),
    .B(_09860_),
    .X(_09861_));
 sky130_fd_sc_hd__o211a_1 _22717_ (.A1(_09415_),
    .A2(_09859_),
    .B1(_09861_),
    .C1(_09489_),
    .X(_09862_));
 sky130_fd_sc_hd__mux4_1 _22718_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][21] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][21] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][21] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][21] ),
    .S0(_09464_),
    .S1(_09467_),
    .X(_09863_));
 sky130_fd_sc_hd__mux4_1 _22719_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][21] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][21] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][21] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][21] ),
    .S0(_09477_),
    .S1(_09466_),
    .X(_09864_));
 sky130_fd_sc_hd__or2_1 _22720_ (.A(_09482_),
    .B(_09864_),
    .X(_09865_));
 sky130_fd_sc_hd__o211a_1 _22721_ (.A1(_09476_),
    .A2(_09863_),
    .B1(_09865_),
    .C1(_09474_),
    .X(_09866_));
 sky130_fd_sc_hd__o31a_1 _22722_ (.A1(_09858_),
    .A2(_09862_),
    .A3(_09866_),
    .B1(_09491_),
    .X(_01145_));
 sky130_fd_sc_hd__mux4_1 _22723_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][22] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][22] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][22] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][22] ),
    .S0(_09385_),
    .S1(_09637_),
    .X(_09867_));
 sky130_fd_sc_hd__mux4_1 _22724_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][22] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][22] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][22] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][22] ),
    .S0(_09406_),
    .S1(_09395_),
    .X(_09868_));
 sky130_fd_sc_hd__or2_1 _22725_ (.A(_09516_),
    .B(_09868_),
    .X(_09869_));
 sky130_fd_sc_hd__o211a_1 _22726_ (.A1(_09636_),
    .A2(_09867_),
    .B1(_09869_),
    .C1(_09510_),
    .X(_09870_));
 sky130_fd_sc_hd__mux4_1 _22727_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][22] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][22] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][22] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][22] ),
    .S0(_09443_),
    .S1(_09453_),
    .X(_09871_));
 sky130_fd_sc_hd__mux4_1 _22728_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][22] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][22] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][22] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][22] ),
    .S0(_09393_),
    .S1(_09465_),
    .X(_09872_));
 sky130_fd_sc_hd__or2_1 _22729_ (.A(_09391_),
    .B(_09872_),
    .X(_09873_));
 sky130_fd_sc_hd__o211a_1 _22730_ (.A1(_09452_),
    .A2(_09871_),
    .B1(_09873_),
    .C1(_09457_),
    .X(_09874_));
 sky130_fd_sc_hd__o21a_1 _22731_ (.A1(_09870_),
    .A2(_09874_),
    .B1(\rvcpu.dp.plfd.InstrD[24] ),
    .X(_09875_));
 sky130_fd_sc_hd__mux4_1 _22732_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][22] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][22] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][22] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][22] ),
    .S0(_09386_),
    .S1(_09419_),
    .X(_09876_));
 sky130_fd_sc_hd__mux4_1 _22733_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][22] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][22] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][22] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][22] ),
    .S0(_09418_),
    .S1(_09453_),
    .X(_09877_));
 sky130_fd_sc_hd__or2_1 _22734_ (.A(_09636_),
    .B(_09877_),
    .X(_09878_));
 sky130_fd_sc_hd__o211a_1 _22735_ (.A1(_09415_),
    .A2(_09876_),
    .B1(_09878_),
    .C1(_09488_),
    .X(_09879_));
 sky130_fd_sc_hd__mux4_1 _22736_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][22] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][22] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][22] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][22] ),
    .S0(_09464_),
    .S1(_09467_),
    .X(_09880_));
 sky130_fd_sc_hd__mux4_1 _22737_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][22] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][22] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][22] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][22] ),
    .S0(_09477_),
    .S1(_09466_),
    .X(_09881_));
 sky130_fd_sc_hd__or2_1 _22738_ (.A(_09469_),
    .B(_09881_),
    .X(_09882_));
 sky130_fd_sc_hd__o211a_1 _22739_ (.A1(_09476_),
    .A2(_09880_),
    .B1(_09882_),
    .C1(_09474_),
    .X(_09883_));
 sky130_fd_sc_hd__o31a_1 _22740_ (.A1(_09875_),
    .A2(_09879_),
    .A3(_09883_),
    .B1(_09491_),
    .X(_01146_));
 sky130_fd_sc_hd__mux4_1 _22741_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][23] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][23] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][23] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][23] ),
    .S0(_09517_),
    .S1(_09513_),
    .X(_09884_));
 sky130_fd_sc_hd__or2_1 _22742_ (.A(_09511_),
    .B(_09884_),
    .X(_09885_));
 sky130_fd_sc_hd__mux4_2 _22743_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][23] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][23] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][23] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][23] ),
    .S0(_09517_),
    .S1(_09577_),
    .X(_09886_));
 sky130_fd_sc_hd__or2_1 _22744_ (.A(_09398_),
    .B(_09886_),
    .X(_09887_));
 sky130_fd_sc_hd__mux4_1 _22745_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][23] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][23] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][23] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][23] ),
    .S0(_09381_),
    .S1(_09423_),
    .X(_09888_));
 sky130_fd_sc_hd__mux4_1 _22746_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][23] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][23] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][23] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][23] ),
    .S0(_09392_),
    .S1(_09394_),
    .X(_09889_));
 sky130_fd_sc_hd__or2_1 _22747_ (.A(_09390_),
    .B(_09889_),
    .X(_09890_));
 sky130_fd_sc_hd__o211a_1 _22748_ (.A1(_09516_),
    .A2(_09888_),
    .B1(_09890_),
    .C1(_09523_),
    .X(_09891_));
 sky130_fd_sc_hd__a311o_1 _22749_ (.A1(_09510_),
    .A2(_09885_),
    .A3(_09887_),
    .B1(_09891_),
    .C1(_09525_),
    .X(_09892_));
 sky130_fd_sc_hd__mux4_1 _22750_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][23] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][23] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][23] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][23] ),
    .S0(_09714_),
    .S1(_09383_),
    .X(_09893_));
 sky130_fd_sc_hd__mux4_1 _22751_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][23] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][23] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][23] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][23] ),
    .S0(_09416_),
    .S1(_09716_),
    .X(_09894_));
 sky130_fd_sc_hd__a21o_1 _22752_ (.A1(_09433_),
    .A2(_09894_),
    .B1(_09789_),
    .X(_09895_));
 sky130_fd_sc_hd__a21o_1 _22753_ (.A1(_09622_),
    .A2(_09893_),
    .B1(_09895_),
    .X(_09896_));
 sky130_fd_sc_hd__mux4_1 _22754_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][23] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][23] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][23] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][23] ),
    .S0(_09483_),
    .S1(_09656_),
    .X(_09897_));
 sky130_fd_sc_hd__mux4_1 _22755_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][23] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][23] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][23] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][23] ),
    .S0(_09462_),
    .S1(_09721_),
    .X(_09898_));
 sky130_fd_sc_hd__and2_1 _22756_ (.A(_09481_),
    .B(_09898_),
    .X(_09899_));
 sky130_fd_sc_hd__a211o_1 _22757_ (.A1(_09627_),
    .A2(_09897_),
    .B1(_09899_),
    .C1(_09795_),
    .X(_09900_));
 sky130_fd_sc_hd__and4_1 _22758_ (.A(_09705_),
    .B(_09892_),
    .C(_09896_),
    .D(_09900_),
    .X(_09901_));
 sky130_fd_sc_hd__clkbuf_1 _22759_ (.A(_09901_),
    .X(_01147_));
 sky130_fd_sc_hd__mux4_2 _22760_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][24] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][24] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][24] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][24] ),
    .S0(_09406_),
    .S1(_09395_),
    .X(_09902_));
 sky130_fd_sc_hd__or2_1 _22761_ (.A(_09511_),
    .B(_09902_),
    .X(_09903_));
 sky130_fd_sc_hd__mux4_1 _22762_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][24] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][24] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][24] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][24] ),
    .S0(_09446_),
    .S1(_09402_),
    .X(_09904_));
 sky130_fd_sc_hd__o21a_1 _22763_ (.A1(_09451_),
    .A2(_09904_),
    .B1(_09404_),
    .X(_09905_));
 sky130_fd_sc_hd__mux4_1 _22764_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][24] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][24] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][24] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][24] ),
    .S0(_09406_),
    .S1(_09408_),
    .X(_09906_));
 sky130_fd_sc_hd__mux4_1 _22765_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][24] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][24] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][24] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][24] ),
    .S0(_09512_),
    .S1(_09408_),
    .X(_09907_));
 sky130_fd_sc_hd__mux2_1 _22766_ (.A0(_09906_),
    .A1(_09907_),
    .S(_09380_),
    .X(_09908_));
 sky130_fd_sc_hd__a221o_1 _22767_ (.A1(_09903_),
    .A2(_09905_),
    .B1(_09908_),
    .B2(_09412_),
    .C1(_09525_),
    .X(_09909_));
 sky130_fd_sc_hd__mux4_1 _22768_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][24] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][24] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][24] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][24] ),
    .S0(_09714_),
    .S1(_09383_),
    .X(_09910_));
 sky130_fd_sc_hd__mux4_1 _22769_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][24] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][24] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][24] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][24] ),
    .S0(_09416_),
    .S1(_09716_),
    .X(_09911_));
 sky130_fd_sc_hd__a21o_1 _22770_ (.A1(_09433_),
    .A2(_09911_),
    .B1(_09789_),
    .X(_09912_));
 sky130_fd_sc_hd__a21o_1 _22771_ (.A1(_09429_),
    .A2(_09910_),
    .B1(_09912_),
    .X(_09913_));
 sky130_fd_sc_hd__mux4_1 _22772_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][24] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][24] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][24] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][24] ),
    .S0(_09483_),
    .S1(_09656_),
    .X(_09914_));
 sky130_fd_sc_hd__mux4_1 _22773_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][24] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][24] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][24] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][24] ),
    .S0(_09462_),
    .S1(_09721_),
    .X(_09915_));
 sky130_fd_sc_hd__and2_1 _22774_ (.A(_09481_),
    .B(_09915_),
    .X(_09916_));
 sky130_fd_sc_hd__a211o_1 _22775_ (.A1(_09452_),
    .A2(_09914_),
    .B1(_09916_),
    .C1(_09795_),
    .X(_09917_));
 sky130_fd_sc_hd__and4_1 _22776_ (.A(_09705_),
    .B(_09909_),
    .C(_09913_),
    .D(_09917_),
    .X(_09918_));
 sky130_fd_sc_hd__clkbuf_1 _22777_ (.A(_09918_),
    .X(_01148_));
 sky130_fd_sc_hd__mux4_1 _22778_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][25] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][25] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][25] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][25] ),
    .S0(_09445_),
    .S1(_09447_),
    .X(_09919_));
 sky130_fd_sc_hd__mux4_1 _22779_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][25] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][25] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][25] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][25] ),
    .S0(_09434_),
    .S1(_09558_),
    .X(_09920_));
 sky130_fd_sc_hd__mux2_2 _22780_ (.A0(_09919_),
    .A1(_09920_),
    .S(_09449_),
    .X(_09921_));
 sky130_fd_sc_hd__mux4_1 _22781_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][25] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][25] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][25] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][25] ),
    .S0(_09463_),
    .S1(_09637_),
    .X(_09922_));
 sky130_fd_sc_hd__nor2_1 _22782_ (.A(_09422_),
    .B(_09922_),
    .Y(_09923_));
 sky130_fd_sc_hd__mux4_1 _22783_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][25] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][25] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][25] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][25] ),
    .S0(_09382_),
    .S1(_09417_),
    .X(_09924_));
 sky130_fd_sc_hd__o21ai_1 _22784_ (.A1(_09495_),
    .A2(_09924_),
    .B1(_09472_),
    .Y(_09925_));
 sky130_fd_sc_hd__o2bb2a_1 _22785_ (.A1_N(_09442_),
    .A2_N(_09921_),
    .B1(_09923_),
    .B2(_09925_),
    .X(_09926_));
 sky130_fd_sc_hd__nor2_1 _22786_ (.A(_09441_),
    .B(_09926_),
    .Y(_09927_));
 sky130_fd_sc_hd__mux4_1 _22787_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][25] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][25] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][25] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][25] ),
    .S0(_09386_),
    .S1(_09419_),
    .X(_09928_));
 sky130_fd_sc_hd__mux4_1 _22788_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][25] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][25] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][25] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][25] ),
    .S0(_09443_),
    .S1(_09453_),
    .X(_09929_));
 sky130_fd_sc_hd__or2_1 _22789_ (.A(_09636_),
    .B(_09929_),
    .X(_09930_));
 sky130_fd_sc_hd__o211a_1 _22790_ (.A1(_09415_),
    .A2(_09928_),
    .B1(_09930_),
    .C1(_09488_),
    .X(_09931_));
 sky130_fd_sc_hd__mux4_1 _22791_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][25] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][25] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][25] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][25] ),
    .S0(_09464_),
    .S1(_09467_),
    .X(_09932_));
 sky130_fd_sc_hd__mux4_1 _22792_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][25] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][25] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][25] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][25] ),
    .S0(_09477_),
    .S1(_09466_),
    .X(_09933_));
 sky130_fd_sc_hd__or2_1 _22793_ (.A(_09469_),
    .B(_09933_),
    .X(_09934_));
 sky130_fd_sc_hd__o211a_1 _22794_ (.A1(_09461_),
    .A2(_09932_),
    .B1(_09934_),
    .C1(_09474_),
    .X(_09935_));
 sky130_fd_sc_hd__o31a_1 _22795_ (.A1(_09927_),
    .A2(_09931_),
    .A3(_09935_),
    .B1(_09491_),
    .X(_01149_));
 sky130_fd_sc_hd__mux4_1 _22796_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][26] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][26] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][26] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][26] ),
    .S0(_09445_),
    .S1(_09447_),
    .X(_09936_));
 sky130_fd_sc_hd__mux4_1 _22797_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][26] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][26] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][26] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][26] ),
    .S0(_09434_),
    .S1(_09558_),
    .X(_09937_));
 sky130_fd_sc_hd__mux2_2 _22798_ (.A0(_09936_),
    .A1(_09937_),
    .S(_09449_),
    .X(_09938_));
 sky130_fd_sc_hd__mux4_1 _22799_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][26] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][26] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][26] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][26] ),
    .S0(_09443_),
    .S1(_09453_),
    .X(_09939_));
 sky130_fd_sc_hd__nor2_1 _22800_ (.A(_09495_),
    .B(_09939_),
    .Y(_09940_));
 sky130_fd_sc_hd__mux4_1 _22801_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][26] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][26] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][26] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][26] ),
    .S0(_09484_),
    .S1(_09431_),
    .X(_09941_));
 sky130_fd_sc_hd__o21ai_1 _22802_ (.A1(_09422_),
    .A2(_09941_),
    .B1(_09472_),
    .Y(_09942_));
 sky130_fd_sc_hd__o2bb2a_1 _22803_ (.A1_N(_09442_),
    .A2_N(_09938_),
    .B1(_09940_),
    .B2(_09942_),
    .X(_09943_));
 sky130_fd_sc_hd__nor2_1 _22804_ (.A(_09441_),
    .B(_09943_),
    .Y(_09944_));
 sky130_fd_sc_hd__mux4_1 _22805_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][26] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][26] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][26] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][26] ),
    .S0(_09386_),
    .S1(_09419_),
    .X(_09945_));
 sky130_fd_sc_hd__mux4_1 _22806_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][26] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][26] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][26] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][26] ),
    .S0(_09463_),
    .S1(_09637_),
    .X(_09946_));
 sky130_fd_sc_hd__or2_1 _22807_ (.A(_09636_),
    .B(_09946_),
    .X(_09947_));
 sky130_fd_sc_hd__o211a_1 _22808_ (.A1(_09415_),
    .A2(_09945_),
    .B1(_09947_),
    .C1(_09473_),
    .X(_09948_));
 sky130_fd_sc_hd__mux4_1 _22809_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][26] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][26] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][26] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][26] ),
    .S0(_09464_),
    .S1(_09467_),
    .X(_09949_));
 sky130_fd_sc_hd__mux4_1 _22810_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][26] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][26] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][26] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][26] ),
    .S0(_09424_),
    .S1(_09485_),
    .X(_09950_));
 sky130_fd_sc_hd__or2_1 _22811_ (.A(_09469_),
    .B(_09950_),
    .X(_09951_));
 sky130_fd_sc_hd__o211a_1 _22812_ (.A1(_09461_),
    .A2(_09949_),
    .B1(_09951_),
    .C1(_09489_),
    .X(_09952_));
 sky130_fd_sc_hd__o31a_1 _22813_ (.A1(_09944_),
    .A2(_09948_),
    .A3(_09952_),
    .B1(_09389_),
    .X(_01150_));
 sky130_fd_sc_hd__mux4_2 _22814_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][27] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][27] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][27] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][27] ),
    .S0(_09406_),
    .S1(_09395_),
    .X(_09953_));
 sky130_fd_sc_hd__or2_1 _22815_ (.A(_09511_),
    .B(_09953_),
    .X(_09954_));
 sky130_fd_sc_hd__mux4_1 _22816_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][27] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][27] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][27] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][27] ),
    .S0(_09446_),
    .S1(_09402_),
    .X(_09955_));
 sky130_fd_sc_hd__o21a_1 _22817_ (.A1(_09451_),
    .A2(_09955_),
    .B1(_09404_),
    .X(_09956_));
 sky130_fd_sc_hd__mux4_1 _22818_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][27] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][27] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][27] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][27] ),
    .S0(_09406_),
    .S1(_09408_),
    .X(_09957_));
 sky130_fd_sc_hd__mux4_1 _22819_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][27] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][27] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][27] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][27] ),
    .S0(_09512_),
    .S1(_09408_),
    .X(_09958_));
 sky130_fd_sc_hd__mux2_1 _22820_ (.A0(_09957_),
    .A1(_09958_),
    .S(_09380_),
    .X(_09959_));
 sky130_fd_sc_hd__a221o_1 _22821_ (.A1(_09954_),
    .A2(_09956_),
    .B1(_09959_),
    .B2(_09411_),
    .C1(_09525_),
    .X(_09960_));
 sky130_fd_sc_hd__mux4_1 _22822_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][27] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][27] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][27] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][27] ),
    .S0(_09714_),
    .S1(_09383_),
    .X(_09961_));
 sky130_fd_sc_hd__mux4_1 _22823_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][27] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][27] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][27] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][27] ),
    .S0(_09416_),
    .S1(_09716_),
    .X(_09962_));
 sky130_fd_sc_hd__a21o_1 _22824_ (.A1(_09433_),
    .A2(_09962_),
    .B1(_09789_),
    .X(_09963_));
 sky130_fd_sc_hd__a21o_1 _22825_ (.A1(_09429_),
    .A2(_09961_),
    .B1(_09963_),
    .X(_09964_));
 sky130_fd_sc_hd__mux4_1 _22826_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][27] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][27] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][27] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][27] ),
    .S0(_09483_),
    .S1(_09656_),
    .X(_09965_));
 sky130_fd_sc_hd__mux4_1 _22827_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][27] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][27] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][27] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][27] ),
    .S0(_09462_),
    .S1(_09721_),
    .X(_09966_));
 sky130_fd_sc_hd__and2_1 _22828_ (.A(_09481_),
    .B(_09966_),
    .X(_09967_));
 sky130_fd_sc_hd__a211o_1 _22829_ (.A1(_09452_),
    .A2(_09965_),
    .B1(_09967_),
    .C1(_09795_),
    .X(_09968_));
 sky130_fd_sc_hd__and4_1 _22830_ (.A(_09705_),
    .B(_09960_),
    .C(_09964_),
    .D(_09968_),
    .X(_09969_));
 sky130_fd_sc_hd__clkbuf_1 _22831_ (.A(_09969_),
    .X(_01151_));
 sky130_fd_sc_hd__mux4_1 _22832_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][28] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][28] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][28] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][28] ),
    .S0(_09445_),
    .S1(_09447_),
    .X(_09970_));
 sky130_fd_sc_hd__mux4_1 _22833_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][28] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][28] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][28] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][28] ),
    .S0(_09434_),
    .S1(_09558_),
    .X(_09971_));
 sky130_fd_sc_hd__mux2_1 _22834_ (.A0(_09970_),
    .A1(_09971_),
    .S(_09449_),
    .X(_09972_));
 sky130_fd_sc_hd__mux4_1 _22835_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][28] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][28] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][28] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][28] ),
    .S0(_09385_),
    .S1(_09637_),
    .X(_09973_));
 sky130_fd_sc_hd__nor2_1 _22836_ (.A(_09422_),
    .B(_09973_),
    .Y(_09974_));
 sky130_fd_sc_hd__mux4_1 _22837_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][28] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][28] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][28] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][28] ),
    .S0(_09382_),
    .S1(_09417_),
    .X(_09975_));
 sky130_fd_sc_hd__o21ai_1 _22838_ (.A1(_09495_),
    .A2(_09975_),
    .B1(_09472_),
    .Y(_09976_));
 sky130_fd_sc_hd__o2bb2a_1 _22839_ (.A1_N(_09442_),
    .A2_N(_09972_),
    .B1(_09974_),
    .B2(_09976_),
    .X(_09977_));
 sky130_fd_sc_hd__nor2_1 _22840_ (.A(_09413_),
    .B(_09977_),
    .Y(_09978_));
 sky130_fd_sc_hd__mux4_1 _22841_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][28] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][28] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][28] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][28] ),
    .S0(_09386_),
    .S1(_09419_),
    .X(_09979_));
 sky130_fd_sc_hd__mux4_1 _22842_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][28] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][28] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][28] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][28] ),
    .S0(_09463_),
    .S1(_09637_),
    .X(_09980_));
 sky130_fd_sc_hd__or2_1 _22843_ (.A(_09636_),
    .B(_09980_),
    .X(_09981_));
 sky130_fd_sc_hd__o211a_1 _22844_ (.A1(_09415_),
    .A2(_09979_),
    .B1(_09981_),
    .C1(_09473_),
    .X(_09982_));
 sky130_fd_sc_hd__mux4_1 _22845_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][28] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][28] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][28] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][28] ),
    .S0(_09464_),
    .S1(_09467_),
    .X(_09983_));
 sky130_fd_sc_hd__mux4_1 _22846_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][28] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][28] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][28] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][28] ),
    .S0(_09424_),
    .S1(_09485_),
    .X(_09984_));
 sky130_fd_sc_hd__or2_1 _22847_ (.A(_09469_),
    .B(_09984_),
    .X(_09985_));
 sky130_fd_sc_hd__o211a_1 _22848_ (.A1(_09461_),
    .A2(_09983_),
    .B1(_09985_),
    .C1(_09489_),
    .X(_09986_));
 sky130_fd_sc_hd__o31a_1 _22849_ (.A1(_09978_),
    .A2(_09982_),
    .A3(_09986_),
    .B1(_09389_),
    .X(_01152_));
 sky130_fd_sc_hd__mux4_1 _22850_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][29] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][29] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][29] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][29] ),
    .S0(_09517_),
    .S1(_09513_),
    .X(_09987_));
 sky130_fd_sc_hd__or2_1 _22851_ (.A(_09380_),
    .B(_09987_),
    .X(_09988_));
 sky130_fd_sc_hd__mux4_1 _22852_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][29] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][29] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][29] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][29] ),
    .S0(_09384_),
    .S1(_09577_),
    .X(_09989_));
 sky130_fd_sc_hd__or2_1 _22853_ (.A(_09398_),
    .B(_09989_),
    .X(_09990_));
 sky130_fd_sc_hd__mux4_1 _22854_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][29] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][29] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][29] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][29] ),
    .S0(_09381_),
    .S1(_09423_),
    .X(_09991_));
 sky130_fd_sc_hd__mux4_1 _22855_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][29] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][29] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][29] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][29] ),
    .S0(_08592_),
    .S1(_09394_),
    .X(_09992_));
 sky130_fd_sc_hd__or2_1 _22856_ (.A(_09390_),
    .B(_09992_),
    .X(_09993_));
 sky130_fd_sc_hd__o211a_1 _22857_ (.A1(_09516_),
    .A2(_09991_),
    .B1(_09993_),
    .C1(_09523_),
    .X(_09994_));
 sky130_fd_sc_hd__a311o_1 _22858_ (.A1(_09510_),
    .A2(_09988_),
    .A3(_09990_),
    .B1(_09994_),
    .C1(_09525_),
    .X(_09995_));
 sky130_fd_sc_hd__mux4_1 _22859_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][29] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][29] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][29] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][29] ),
    .S0(_09477_),
    .S1(_09383_),
    .X(_09996_));
 sky130_fd_sc_hd__mux4_1 _22860_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][29] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][29] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][29] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][29] ),
    .S0(_09416_),
    .S1(_09418_),
    .X(_09997_));
 sky130_fd_sc_hd__a21o_1 _22861_ (.A1(_09433_),
    .A2(_09997_),
    .B1(_09789_),
    .X(_09998_));
 sky130_fd_sc_hd__a21o_1 _22862_ (.A1(_09429_),
    .A2(_09996_),
    .B1(_09998_),
    .X(_09999_));
 sky130_fd_sc_hd__mux4_1 _22863_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][29] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][29] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][29] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][29] ),
    .S0(_09483_),
    .S1(_09656_),
    .X(_10000_));
 sky130_fd_sc_hd__mux4_1 _22864_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][29] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][29] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][29] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][29] ),
    .S0(_09462_),
    .S1(_09465_),
    .X(_10001_));
 sky130_fd_sc_hd__and2_1 _22865_ (.A(_09481_),
    .B(_10001_),
    .X(_10002_));
 sky130_fd_sc_hd__a211o_1 _22866_ (.A1(_09452_),
    .A2(_10000_),
    .B1(_10002_),
    .C1(_09795_),
    .X(_10003_));
 sky130_fd_sc_hd__and4_1 _22867_ (.A(_09388_),
    .B(_09995_),
    .C(_09999_),
    .D(_10003_),
    .X(_10004_));
 sky130_fd_sc_hd__clkbuf_1 _22868_ (.A(_10004_),
    .X(_01153_));
 sky130_fd_sc_hd__mux4_1 _22869_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][30] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][30] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][30] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][30] ),
    .S0(_09517_),
    .S1(_09513_),
    .X(_10005_));
 sky130_fd_sc_hd__or2_1 _22870_ (.A(_09380_),
    .B(_10005_),
    .X(_10006_));
 sky130_fd_sc_hd__mux4_1 _22871_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][30] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][30] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][30] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][30] ),
    .S0(_09384_),
    .S1(_09577_),
    .X(_10007_));
 sky130_fd_sc_hd__or2_1 _22872_ (.A(_09398_),
    .B(_10007_),
    .X(_10008_));
 sky130_fd_sc_hd__mux4_1 _22873_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][30] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][30] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][30] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][30] ),
    .S0(_09381_),
    .S1(_09423_),
    .X(_10009_));
 sky130_fd_sc_hd__mux4_1 _22874_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][30] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][30] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][30] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][30] ),
    .S0(_08592_),
    .S1(_08595_),
    .X(_10010_));
 sky130_fd_sc_hd__or2_1 _22875_ (.A(_09390_),
    .B(_10010_),
    .X(_10011_));
 sky130_fd_sc_hd__o211a_1 _22876_ (.A1(_09516_),
    .A2(_10009_),
    .B1(_10011_),
    .C1(_09523_),
    .X(_10012_));
 sky130_fd_sc_hd__a311o_1 _22877_ (.A1(_09510_),
    .A2(_10006_),
    .A3(_10008_),
    .B1(_10012_),
    .C1(_08589_),
    .X(_10013_));
 sky130_fd_sc_hd__mux4_1 _22878_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][30] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][30] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][30] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][30] ),
    .S0(_09477_),
    .S1(_09383_),
    .X(_10014_));
 sky130_fd_sc_hd__mux4_1 _22879_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][30] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][30] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][30] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][30] ),
    .S0(_09416_),
    .S1(_09418_),
    .X(_10015_));
 sky130_fd_sc_hd__a21o_1 _22880_ (.A1(_09433_),
    .A2(_10015_),
    .B1(_09789_),
    .X(_10016_));
 sky130_fd_sc_hd__a21o_1 _22881_ (.A1(_09429_),
    .A2(_10014_),
    .B1(_10016_),
    .X(_10017_));
 sky130_fd_sc_hd__mux4_1 _22882_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][30] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][30] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][30] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][30] ),
    .S0(_09483_),
    .S1(_09656_),
    .X(_10018_));
 sky130_fd_sc_hd__mux4_1 _22883_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][30] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][30] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][30] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][30] ),
    .S0(_09462_),
    .S1(_09465_),
    .X(_10019_));
 sky130_fd_sc_hd__and2_1 _22884_ (.A(_09481_),
    .B(_10019_),
    .X(_10020_));
 sky130_fd_sc_hd__a211o_1 _22885_ (.A1(_09452_),
    .A2(_10018_),
    .B1(_10020_),
    .C1(_09795_),
    .X(_10021_));
 sky130_fd_sc_hd__and4_1 _22886_ (.A(_09388_),
    .B(_10013_),
    .C(_10017_),
    .D(_10021_),
    .X(_10022_));
 sky130_fd_sc_hd__clkbuf_1 _22887_ (.A(_10022_),
    .X(_01154_));
 sky130_fd_sc_hd__mux4_1 _22888_ (.A0(\rvcpu.dp.rf.reg_file_arr[16][31] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[17][31] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[18][31] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[19][31] ),
    .S0(_09517_),
    .S1(_09513_),
    .X(_10023_));
 sky130_fd_sc_hd__or2_1 _22889_ (.A(_09380_),
    .B(_10023_),
    .X(_10024_));
 sky130_fd_sc_hd__mux4_1 _22890_ (.A0(\rvcpu.dp.rf.reg_file_arr[20][31] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[21][31] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[22][31] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[23][31] ),
    .S0(_09384_),
    .S1(_09577_),
    .X(_10025_));
 sky130_fd_sc_hd__or2_1 _22891_ (.A(_09398_),
    .B(_10025_),
    .X(_10026_));
 sky130_fd_sc_hd__mux4_1 _22892_ (.A0(\rvcpu.dp.rf.reg_file_arr[28][31] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[30][31] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[29][31] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[31][31] ),
    .S0(_09381_),
    .S1(_09423_),
    .X(_10027_));
 sky130_fd_sc_hd__mux4_1 _22893_ (.A0(\rvcpu.dp.rf.reg_file_arr[24][31] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[25][31] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[26][31] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[27][31] ),
    .S0(_08592_),
    .S1(_08595_),
    .X(_10028_));
 sky130_fd_sc_hd__or2_1 _22894_ (.A(\rvcpu.dp.plfd.InstrD[22] ),
    .B(_10028_),
    .X(_10029_));
 sky130_fd_sc_hd__o211a_1 _22895_ (.A1(_09516_),
    .A2(_10027_),
    .B1(_10029_),
    .C1(_09404_),
    .X(_10030_));
 sky130_fd_sc_hd__a311o_1 _22896_ (.A1(_09510_),
    .A2(_10024_),
    .A3(_10026_),
    .B1(_10030_),
    .C1(_08589_),
    .X(_10031_));
 sky130_fd_sc_hd__mux4_1 _22897_ (.A0(\rvcpu.dp.rf.reg_file_arr[0][31] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[1][31] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[2][31] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[3][31] ),
    .S0(_09477_),
    .S1(_09383_),
    .X(_10032_));
 sky130_fd_sc_hd__mux4_1 _22898_ (.A0(\rvcpu.dp.rf.reg_file_arr[4][31] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[5][31] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[6][31] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[7][31] ),
    .S0(_09416_),
    .S1(_09418_),
    .X(_10033_));
 sky130_fd_sc_hd__a21o_1 _22899_ (.A1(_09433_),
    .A2(_10033_),
    .B1(_09789_),
    .X(_10034_));
 sky130_fd_sc_hd__a21o_1 _22900_ (.A1(_09429_),
    .A2(_10032_),
    .B1(_10034_),
    .X(_10035_));
 sky130_fd_sc_hd__mux4_1 _22901_ (.A0(\rvcpu.dp.rf.reg_file_arr[8][31] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[10][31] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[9][31] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[11][31] ),
    .S0(_09483_),
    .S1(_09656_),
    .X(_10036_));
 sky130_fd_sc_hd__mux4_1 _22902_ (.A0(\rvcpu.dp.rf.reg_file_arr[12][31] ),
    .A1(\rvcpu.dp.rf.reg_file_arr[13][31] ),
    .A2(\rvcpu.dp.rf.reg_file_arr[14][31] ),
    .A3(\rvcpu.dp.rf.reg_file_arr[15][31] ),
    .S0(_09462_),
    .S1(_09465_),
    .X(_10037_));
 sky130_fd_sc_hd__and2_1 _22903_ (.A(_09481_),
    .B(_10037_),
    .X(_10038_));
 sky130_fd_sc_hd__a211o_1 _22904_ (.A1(_09452_),
    .A2(_10036_),
    .B1(_10038_),
    .C1(_09795_),
    .X(_10039_));
 sky130_fd_sc_hd__and4_1 _22905_ (.A(_09388_),
    .B(_10031_),
    .C(_10035_),
    .D(_10039_),
    .X(_10040_));
 sky130_fd_sc_hd__clkbuf_1 _22906_ (.A(_10040_),
    .X(_01155_));
 sky130_fd_sc_hd__buf_4 _22907_ (.A(_06587_),
    .X(_10041_));
 sky130_fd_sc_hd__buf_4 _22908_ (.A(_08144_),
    .X(_10042_));
 sky130_fd_sc_hd__a21oi_4 _22909_ (.A1(_09217_),
    .A2(_09262_),
    .B1(_09220_),
    .Y(_10043_));
 sky130_fd_sc_hd__clkbuf_4 _22910_ (.A(_10043_),
    .X(_10044_));
 sky130_fd_sc_hd__or3_1 _22911_ (.A(_07019_),
    .B(_10042_),
    .C(_10044_),
    .X(_10045_));
 sky130_fd_sc_hd__buf_2 _22912_ (.A(_10045_),
    .X(_10046_));
 sky130_fd_sc_hd__clkbuf_4 _22913_ (.A(\rvcpu.dp.plem.WriteDataM[0] ),
    .X(_10047_));
 sky130_fd_sc_hd__buf_2 _22914_ (.A(_10047_),
    .X(_10048_));
 sky130_fd_sc_hd__nor2_1 _22915_ (.A(_06604_),
    .B(_07154_),
    .Y(_10049_));
 sky130_fd_sc_hd__a21o_2 _22916_ (.A1(_09217_),
    .A2(_09262_),
    .B1(_09220_),
    .X(_10050_));
 sky130_fd_sc_hd__buf_6 _22917_ (.A(_10050_),
    .X(_10051_));
 sky130_fd_sc_hd__buf_2 _22918_ (.A(_10051_),
    .X(_10052_));
 sky130_fd_sc_hd__and3_2 _22919_ (.A(_09299_),
    .B(_10049_),
    .C(_10052_),
    .X(_10053_));
 sky130_fd_sc_hd__and2_1 _22920_ (.A(_10048_),
    .B(_10053_),
    .X(_10054_));
 sky130_fd_sc_hd__a31o_1 _22921_ (.A1(_10041_),
    .A2(\datamem.data_ram[5][0] ),
    .A3(_10046_),
    .B1(_10054_),
    .X(_01156_));
 sky130_fd_sc_hd__buf_2 _22922_ (.A(_06587_),
    .X(_10055_));
 sky130_fd_sc_hd__clkbuf_4 _22923_ (.A(_10055_),
    .X(_10056_));
 sky130_fd_sc_hd__buf_4 _22924_ (.A(\rvcpu.dp.plem.WriteDataM[1] ),
    .X(_10057_));
 sky130_fd_sc_hd__buf_2 _22925_ (.A(_10057_),
    .X(_10058_));
 sky130_fd_sc_hd__and2_1 _22926_ (.A(_10058_),
    .B(_10053_),
    .X(_10059_));
 sky130_fd_sc_hd__a31o_1 _22927_ (.A1(_10056_),
    .A2(\datamem.data_ram[5][1] ),
    .A3(_10046_),
    .B1(_10059_),
    .X(_01157_));
 sky130_fd_sc_hd__clkbuf_4 _22928_ (.A(\rvcpu.dp.plem.WriteDataM[2] ),
    .X(_10060_));
 sky130_fd_sc_hd__buf_2 _22929_ (.A(_10060_),
    .X(_10061_));
 sky130_fd_sc_hd__and2_1 _22930_ (.A(_10061_),
    .B(_10053_),
    .X(_10062_));
 sky130_fd_sc_hd__a31o_1 _22931_ (.A1(_10056_),
    .A2(\datamem.data_ram[5][2] ),
    .A3(_10046_),
    .B1(_10062_),
    .X(_01158_));
 sky130_fd_sc_hd__buf_4 _22932_ (.A(\rvcpu.dp.plem.WriteDataM[3] ),
    .X(_10063_));
 sky130_fd_sc_hd__buf_2 _22933_ (.A(_10063_),
    .X(_10064_));
 sky130_fd_sc_hd__and2_1 _22934_ (.A(_10064_),
    .B(_10053_),
    .X(_10065_));
 sky130_fd_sc_hd__a31o_1 _22935_ (.A1(_10056_),
    .A2(\datamem.data_ram[5][3] ),
    .A3(_10046_),
    .B1(_10065_),
    .X(_01159_));
 sky130_fd_sc_hd__buf_4 _22936_ (.A(\rvcpu.dp.plem.WriteDataM[4] ),
    .X(_10066_));
 sky130_fd_sc_hd__buf_2 _22937_ (.A(_10066_),
    .X(_10067_));
 sky130_fd_sc_hd__and2_1 _22938_ (.A(_10067_),
    .B(_10053_),
    .X(_10068_));
 sky130_fd_sc_hd__a31o_1 _22939_ (.A1(_10056_),
    .A2(\datamem.data_ram[5][4] ),
    .A3(_10046_),
    .B1(_10068_),
    .X(_01160_));
 sky130_fd_sc_hd__buf_4 _22940_ (.A(\rvcpu.dp.plem.WriteDataM[5] ),
    .X(_10069_));
 sky130_fd_sc_hd__buf_2 _22941_ (.A(_10069_),
    .X(_10070_));
 sky130_fd_sc_hd__and2_1 _22942_ (.A(_10070_),
    .B(_10053_),
    .X(_10071_));
 sky130_fd_sc_hd__a31o_1 _22943_ (.A1(_10056_),
    .A2(\datamem.data_ram[5][5] ),
    .A3(_10046_),
    .B1(_10071_),
    .X(_01161_));
 sky130_fd_sc_hd__buf_4 _22944_ (.A(\rvcpu.dp.plem.WriteDataM[6] ),
    .X(_10072_));
 sky130_fd_sc_hd__clkbuf_4 _22945_ (.A(_10072_),
    .X(_10073_));
 sky130_fd_sc_hd__and2_1 _22946_ (.A(_10073_),
    .B(_10053_),
    .X(_10074_));
 sky130_fd_sc_hd__a31o_1 _22947_ (.A1(_10056_),
    .A2(\datamem.data_ram[5][6] ),
    .A3(_10046_),
    .B1(_10074_),
    .X(_01162_));
 sky130_fd_sc_hd__clkbuf_4 _22948_ (.A(\rvcpu.dp.plem.WriteDataM[7] ),
    .X(_10075_));
 sky130_fd_sc_hd__buf_2 _22949_ (.A(_10075_),
    .X(_10076_));
 sky130_fd_sc_hd__and2_1 _22950_ (.A(_10076_),
    .B(_10053_),
    .X(_10077_));
 sky130_fd_sc_hd__a31o_1 _22951_ (.A1(_10056_),
    .A2(\datamem.data_ram[5][7] ),
    .A3(_10046_),
    .B1(_10077_),
    .X(_01163_));
 sky130_fd_sc_hd__buf_1 _22952_ (.A(clk),
    .X(_10078_));
 sky130_fd_sc_hd__buf_1 _22953_ (.A(_10078_),
    .X(_10079_));
 sky130_fd_sc_hd__buf_1 _22954_ (.A(_10079_),
    .X(_10080_));
 sky130_fd_sc_hd__buf_1 _22955_ (.A(_10080_),
    .X(_10081_));
 sky130_fd_sc_hd__inv_2 _22956_ (.A(_10081_),
    .Y(_00004_));
 sky130_fd_sc_hd__inv_2 _22957_ (.A(_10081_),
    .Y(_00005_));
 sky130_fd_sc_hd__inv_2 _22958_ (.A(_10081_),
    .Y(_00006_));
 sky130_fd_sc_hd__inv_2 _22959_ (.A(_10081_),
    .Y(_00007_));
 sky130_fd_sc_hd__inv_2 _22960_ (.A(_10081_),
    .Y(_00008_));
 sky130_fd_sc_hd__inv_2 _22961_ (.A(_10081_),
    .Y(_00009_));
 sky130_fd_sc_hd__inv_2 _22962_ (.A(_10081_),
    .Y(_00010_));
 sky130_fd_sc_hd__inv_2 _22963_ (.A(_10081_),
    .Y(_00011_));
 sky130_fd_sc_hd__inv_2 _22964_ (.A(_10081_),
    .Y(_00012_));
 sky130_fd_sc_hd__inv_2 _22965_ (.A(_10081_),
    .Y(_00013_));
 sky130_fd_sc_hd__buf_1 _22966_ (.A(_10080_),
    .X(_10082_));
 sky130_fd_sc_hd__inv_2 _22967_ (.A(_10082_),
    .Y(_00014_));
 sky130_fd_sc_hd__inv_2 _22968_ (.A(_10082_),
    .Y(_00015_));
 sky130_fd_sc_hd__inv_2 _22969_ (.A(_10082_),
    .Y(_00016_));
 sky130_fd_sc_hd__inv_2 _22970_ (.A(_10082_),
    .Y(_00017_));
 sky130_fd_sc_hd__inv_2 _22971_ (.A(_10082_),
    .Y(_00018_));
 sky130_fd_sc_hd__inv_2 _22972_ (.A(_10082_),
    .Y(_00019_));
 sky130_fd_sc_hd__inv_2 _22973_ (.A(_10082_),
    .Y(_00020_));
 sky130_fd_sc_hd__inv_2 _22974_ (.A(_10082_),
    .Y(_00021_));
 sky130_fd_sc_hd__inv_2 _22975_ (.A(_10082_),
    .Y(_00022_));
 sky130_fd_sc_hd__inv_2 _22976_ (.A(_10082_),
    .Y(_00023_));
 sky130_fd_sc_hd__buf_1 _22977_ (.A(_10080_),
    .X(_10083_));
 sky130_fd_sc_hd__inv_2 _22978_ (.A(_10083_),
    .Y(_00024_));
 sky130_fd_sc_hd__inv_2 _22979_ (.A(_10083_),
    .Y(_00025_));
 sky130_fd_sc_hd__inv_2 _22980_ (.A(_10083_),
    .Y(_00026_));
 sky130_fd_sc_hd__inv_2 _22981_ (.A(_10083_),
    .Y(_00027_));
 sky130_fd_sc_hd__inv_2 _22982_ (.A(_10083_),
    .Y(_00028_));
 sky130_fd_sc_hd__inv_2 _22983_ (.A(_10083_),
    .Y(_00029_));
 sky130_fd_sc_hd__inv_2 _22984_ (.A(_10083_),
    .Y(_00030_));
 sky130_fd_sc_hd__inv_2 _22985_ (.A(_10083_),
    .Y(_00031_));
 sky130_fd_sc_hd__inv_2 _22986_ (.A(_10083_),
    .Y(_00032_));
 sky130_fd_sc_hd__inv_2 _22987_ (.A(_10083_),
    .Y(_00033_));
 sky130_fd_sc_hd__buf_1 _22988_ (.A(_10080_),
    .X(_10084_));
 sky130_fd_sc_hd__inv_2 _22989_ (.A(_10084_),
    .Y(_00034_));
 sky130_fd_sc_hd__inv_2 _22990_ (.A(_10084_),
    .Y(_00035_));
 sky130_fd_sc_hd__inv_2 _22991_ (.A(_10084_),
    .Y(_00036_));
 sky130_fd_sc_hd__inv_2 _22992_ (.A(_10084_),
    .Y(_00037_));
 sky130_fd_sc_hd__inv_2 _22993_ (.A(_10084_),
    .Y(_00038_));
 sky130_fd_sc_hd__inv_2 _22994_ (.A(_10084_),
    .Y(_00039_));
 sky130_fd_sc_hd__inv_2 _22995_ (.A(_10084_),
    .Y(_00040_));
 sky130_fd_sc_hd__inv_2 _22996_ (.A(_10084_),
    .Y(_00041_));
 sky130_fd_sc_hd__inv_2 _22997_ (.A(_10084_),
    .Y(_00042_));
 sky130_fd_sc_hd__inv_2 _22998_ (.A(_10084_),
    .Y(_00043_));
 sky130_fd_sc_hd__buf_1 _22999_ (.A(_10080_),
    .X(_10085_));
 sky130_fd_sc_hd__inv_2 _23000_ (.A(_10085_),
    .Y(_00044_));
 sky130_fd_sc_hd__inv_2 _23001_ (.A(_10085_),
    .Y(_00045_));
 sky130_fd_sc_hd__inv_2 _23002_ (.A(_10085_),
    .Y(_00046_));
 sky130_fd_sc_hd__inv_2 _23003_ (.A(_10085_),
    .Y(_00047_));
 sky130_fd_sc_hd__inv_2 _23004_ (.A(_10085_),
    .Y(_00048_));
 sky130_fd_sc_hd__inv_2 _23005_ (.A(_10085_),
    .Y(_00049_));
 sky130_fd_sc_hd__inv_2 _23006_ (.A(_10085_),
    .Y(_00050_));
 sky130_fd_sc_hd__inv_2 _23007_ (.A(_10085_),
    .Y(_00051_));
 sky130_fd_sc_hd__inv_2 _23008_ (.A(_10085_),
    .Y(_00052_));
 sky130_fd_sc_hd__inv_2 _23009_ (.A(_10085_),
    .Y(_00053_));
 sky130_fd_sc_hd__buf_1 _23010_ (.A(_10080_),
    .X(_10086_));
 sky130_fd_sc_hd__inv_2 _23011_ (.A(_10086_),
    .Y(_00054_));
 sky130_fd_sc_hd__inv_2 _23012_ (.A(_10086_),
    .Y(_00055_));
 sky130_fd_sc_hd__inv_2 _23013_ (.A(_10086_),
    .Y(_00056_));
 sky130_fd_sc_hd__inv_2 _23014_ (.A(_10086_),
    .Y(_00057_));
 sky130_fd_sc_hd__inv_2 _23015_ (.A(_10086_),
    .Y(_00058_));
 sky130_fd_sc_hd__inv_2 _23016_ (.A(_10086_),
    .Y(_00059_));
 sky130_fd_sc_hd__inv_2 _23017_ (.A(_10086_),
    .Y(_00060_));
 sky130_fd_sc_hd__inv_2 _23018_ (.A(_10086_),
    .Y(_00061_));
 sky130_fd_sc_hd__inv_2 _23019_ (.A(_10086_),
    .Y(_00062_));
 sky130_fd_sc_hd__inv_2 _23020_ (.A(_10086_),
    .Y(_00063_));
 sky130_fd_sc_hd__buf_1 _23021_ (.A(_10079_),
    .X(_10087_));
 sky130_fd_sc_hd__buf_1 _23022_ (.A(_10087_),
    .X(_10088_));
 sky130_fd_sc_hd__inv_2 _23023_ (.A(_10088_),
    .Y(_00064_));
 sky130_fd_sc_hd__inv_2 _23024_ (.A(_10088_),
    .Y(_00065_));
 sky130_fd_sc_hd__inv_2 _23025_ (.A(_10088_),
    .Y(_00066_));
 sky130_fd_sc_hd__inv_2 _23026_ (.A(_10088_),
    .Y(_00067_));
 sky130_fd_sc_hd__inv_2 _23027_ (.A(_10088_),
    .Y(_00068_));
 sky130_fd_sc_hd__inv_2 _23028_ (.A(_10088_),
    .Y(_00069_));
 sky130_fd_sc_hd__inv_2 _23029_ (.A(_10088_),
    .Y(_00070_));
 sky130_fd_sc_hd__inv_2 _23030_ (.A(_10088_),
    .Y(_00071_));
 sky130_fd_sc_hd__inv_2 _23031_ (.A(_10088_),
    .Y(_00072_));
 sky130_fd_sc_hd__inv_2 _23032_ (.A(_10088_),
    .Y(_00073_));
 sky130_fd_sc_hd__buf_1 _23033_ (.A(_10087_),
    .X(_10089_));
 sky130_fd_sc_hd__inv_2 _23034_ (.A(_10089_),
    .Y(_00074_));
 sky130_fd_sc_hd__inv_2 _23035_ (.A(_10089_),
    .Y(_00075_));
 sky130_fd_sc_hd__inv_2 _23036_ (.A(_10089_),
    .Y(_00076_));
 sky130_fd_sc_hd__inv_2 _23037_ (.A(_10089_),
    .Y(_00077_));
 sky130_fd_sc_hd__inv_2 _23038_ (.A(_10089_),
    .Y(_00078_));
 sky130_fd_sc_hd__inv_2 _23039_ (.A(_10089_),
    .Y(_00079_));
 sky130_fd_sc_hd__inv_2 _23040_ (.A(_10089_),
    .Y(_00080_));
 sky130_fd_sc_hd__inv_2 _23041_ (.A(_10089_),
    .Y(_00081_));
 sky130_fd_sc_hd__inv_2 _23042_ (.A(_10089_),
    .Y(_00082_));
 sky130_fd_sc_hd__inv_2 _23043_ (.A(_10089_),
    .Y(_00083_));
 sky130_fd_sc_hd__buf_1 _23044_ (.A(_10087_),
    .X(_10090_));
 sky130_fd_sc_hd__inv_2 _23045_ (.A(_10090_),
    .Y(_00084_));
 sky130_fd_sc_hd__inv_2 _23046_ (.A(_10090_),
    .Y(_00085_));
 sky130_fd_sc_hd__inv_2 _23047_ (.A(_10090_),
    .Y(_00086_));
 sky130_fd_sc_hd__inv_2 _23048_ (.A(_10090_),
    .Y(_00087_));
 sky130_fd_sc_hd__inv_2 _23049_ (.A(_10090_),
    .Y(_00088_));
 sky130_fd_sc_hd__inv_2 _23050_ (.A(_10090_),
    .Y(_00089_));
 sky130_fd_sc_hd__inv_2 _23051_ (.A(_10090_),
    .Y(_00090_));
 sky130_fd_sc_hd__inv_2 _23052_ (.A(_10090_),
    .Y(_00091_));
 sky130_fd_sc_hd__inv_2 _23053_ (.A(_10090_),
    .Y(_00092_));
 sky130_fd_sc_hd__inv_2 _23054_ (.A(_10090_),
    .Y(_00093_));
 sky130_fd_sc_hd__buf_1 _23055_ (.A(_10087_),
    .X(_10091_));
 sky130_fd_sc_hd__inv_2 _23056_ (.A(_10091_),
    .Y(_00094_));
 sky130_fd_sc_hd__inv_2 _23057_ (.A(_10091_),
    .Y(_00095_));
 sky130_fd_sc_hd__inv_2 _23058_ (.A(_10091_),
    .Y(_00096_));
 sky130_fd_sc_hd__inv_2 _23059_ (.A(_10091_),
    .Y(_00097_));
 sky130_fd_sc_hd__inv_2 _23060_ (.A(_10091_),
    .Y(_00098_));
 sky130_fd_sc_hd__inv_2 _23061_ (.A(_10091_),
    .Y(_00099_));
 sky130_fd_sc_hd__nor2_8 _23062_ (.A(_10042_),
    .B(_09268_),
    .Y(_10092_));
 sky130_fd_sc_hd__a21oi_4 _23063_ (.A1(_09299_),
    .A2(_10092_),
    .B1(_09361_),
    .Y(_10093_));
 sky130_fd_sc_hd__mux2_1 _23064_ (.A0(_09267_),
    .A1(\datamem.data_ram[5][8] ),
    .S(_10093_),
    .X(_10094_));
 sky130_fd_sc_hd__clkbuf_1 _23065_ (.A(_10094_),
    .X(_01260_));
 sky130_fd_sc_hd__mux2_1 _23066_ (.A0(_09273_),
    .A1(\datamem.data_ram[5][9] ),
    .S(_10093_),
    .X(_10095_));
 sky130_fd_sc_hd__clkbuf_1 _23067_ (.A(_10095_),
    .X(_01261_));
 sky130_fd_sc_hd__mux2_1 _23068_ (.A0(_09276_),
    .A1(\datamem.data_ram[5][10] ),
    .S(_10093_),
    .X(_10096_));
 sky130_fd_sc_hd__clkbuf_1 _23069_ (.A(_10096_),
    .X(_01262_));
 sky130_fd_sc_hd__mux2_1 _23070_ (.A0(_09279_),
    .A1(\datamem.data_ram[5][11] ),
    .S(_10093_),
    .X(_10097_));
 sky130_fd_sc_hd__clkbuf_1 _23071_ (.A(_10097_),
    .X(_01263_));
 sky130_fd_sc_hd__mux2_1 _23072_ (.A0(_09282_),
    .A1(\datamem.data_ram[5][12] ),
    .S(_10093_),
    .X(_10098_));
 sky130_fd_sc_hd__clkbuf_1 _23073_ (.A(_10098_),
    .X(_01264_));
 sky130_fd_sc_hd__mux2_1 _23074_ (.A0(_09285_),
    .A1(\datamem.data_ram[5][13] ),
    .S(_10093_),
    .X(_10099_));
 sky130_fd_sc_hd__clkbuf_1 _23075_ (.A(_10099_),
    .X(_01265_));
 sky130_fd_sc_hd__mux2_1 _23076_ (.A0(_09288_),
    .A1(\datamem.data_ram[5][14] ),
    .S(_10093_),
    .X(_10100_));
 sky130_fd_sc_hd__clkbuf_1 _23077_ (.A(_10100_),
    .X(_01266_));
 sky130_fd_sc_hd__mux2_1 _23078_ (.A0(_09291_),
    .A1(\datamem.data_ram[5][15] ),
    .S(_10093_),
    .X(_10101_));
 sky130_fd_sc_hd__clkbuf_1 _23079_ (.A(_10101_),
    .X(_01267_));
 sky130_fd_sc_hd__inv_2 _23080_ (.A(_10091_),
    .Y(_00100_));
 sky130_fd_sc_hd__inv_2 _23081_ (.A(_10091_),
    .Y(_00101_));
 sky130_fd_sc_hd__inv_2 _23082_ (.A(_10091_),
    .Y(_00102_));
 sky130_fd_sc_hd__inv_2 _23083_ (.A(_10091_),
    .Y(_00103_));
 sky130_fd_sc_hd__buf_1 _23084_ (.A(_10087_),
    .X(_10102_));
 sky130_fd_sc_hd__inv_2 _23085_ (.A(_10102_),
    .Y(_00104_));
 sky130_fd_sc_hd__inv_2 _23086_ (.A(_10102_),
    .Y(_00105_));
 sky130_fd_sc_hd__inv_2 _23087_ (.A(_10102_),
    .Y(_00106_));
 sky130_fd_sc_hd__inv_2 _23088_ (.A(_10102_),
    .Y(_00107_));
 sky130_fd_sc_hd__inv_2 _23089_ (.A(_10102_),
    .Y(_00108_));
 sky130_fd_sc_hd__inv_2 _23090_ (.A(_10102_),
    .Y(_00109_));
 sky130_fd_sc_hd__inv_2 _23091_ (.A(_10102_),
    .Y(_00110_));
 sky130_fd_sc_hd__inv_2 _23092_ (.A(_10102_),
    .Y(_00111_));
 sky130_fd_sc_hd__inv_2 _23093_ (.A(_10102_),
    .Y(_00112_));
 sky130_fd_sc_hd__inv_2 _23094_ (.A(_10102_),
    .Y(_00113_));
 sky130_fd_sc_hd__buf_1 _23095_ (.A(_10087_),
    .X(_10103_));
 sky130_fd_sc_hd__inv_2 _23096_ (.A(_10103_),
    .Y(_00114_));
 sky130_fd_sc_hd__inv_2 _23097_ (.A(_10103_),
    .Y(_00115_));
 sky130_fd_sc_hd__inv_2 _23098_ (.A(_10103_),
    .Y(_00116_));
 sky130_fd_sc_hd__inv_2 _23099_ (.A(_10103_),
    .Y(_00117_));
 sky130_fd_sc_hd__inv_2 _23100_ (.A(_10103_),
    .Y(_00118_));
 sky130_fd_sc_hd__inv_2 _23101_ (.A(_10103_),
    .Y(_00119_));
 sky130_fd_sc_hd__inv_2 _23102_ (.A(_10103_),
    .Y(_00120_));
 sky130_fd_sc_hd__inv_2 _23103_ (.A(_10103_),
    .Y(_00121_));
 sky130_fd_sc_hd__inv_2 _23104_ (.A(_10103_),
    .Y(_00122_));
 sky130_fd_sc_hd__inv_2 _23105_ (.A(_10103_),
    .Y(_00123_));
 sky130_fd_sc_hd__buf_1 _23106_ (.A(_10087_),
    .X(_10104_));
 sky130_fd_sc_hd__inv_2 _23107_ (.A(_10104_),
    .Y(_00124_));
 sky130_fd_sc_hd__inv_2 _23108_ (.A(_10104_),
    .Y(_00125_));
 sky130_fd_sc_hd__inv_2 _23109_ (.A(_10104_),
    .Y(_00126_));
 sky130_fd_sc_hd__inv_2 _23110_ (.A(_10104_),
    .Y(_00127_));
 sky130_fd_sc_hd__inv_2 _23111_ (.A(_10104_),
    .Y(_00128_));
 sky130_fd_sc_hd__inv_2 _23112_ (.A(_10104_),
    .Y(_00129_));
 sky130_fd_sc_hd__inv_2 _23113_ (.A(_10104_),
    .Y(_00130_));
 sky130_fd_sc_hd__inv_2 _23114_ (.A(_10104_),
    .Y(_00131_));
 sky130_fd_sc_hd__inv_2 _23115_ (.A(_10104_),
    .Y(_00132_));
 sky130_fd_sc_hd__inv_2 _23116_ (.A(_10104_),
    .Y(_00133_));
 sky130_fd_sc_hd__buf_1 _23117_ (.A(_10087_),
    .X(_10105_));
 sky130_fd_sc_hd__inv_2 _23118_ (.A(_10105_),
    .Y(_00134_));
 sky130_fd_sc_hd__inv_2 _23119_ (.A(_10105_),
    .Y(_00135_));
 sky130_fd_sc_hd__inv_2 _23120_ (.A(_10105_),
    .Y(_00136_));
 sky130_fd_sc_hd__inv_2 _23121_ (.A(_10105_),
    .Y(_00137_));
 sky130_fd_sc_hd__inv_2 _23122_ (.A(_10105_),
    .Y(_00138_));
 sky130_fd_sc_hd__inv_2 _23123_ (.A(_10105_),
    .Y(_00139_));
 sky130_fd_sc_hd__inv_2 _23124_ (.A(_10105_),
    .Y(_00140_));
 sky130_fd_sc_hd__inv_2 _23125_ (.A(_10105_),
    .Y(_00141_));
 sky130_fd_sc_hd__inv_2 _23126_ (.A(_10105_),
    .Y(_00142_));
 sky130_fd_sc_hd__inv_2 _23127_ (.A(_10105_),
    .Y(_00143_));
 sky130_fd_sc_hd__buf_1 _23128_ (.A(_10087_),
    .X(_10106_));
 sky130_fd_sc_hd__inv_2 _23129_ (.A(_10106_),
    .Y(_00144_));
 sky130_fd_sc_hd__inv_2 _23130_ (.A(_10106_),
    .Y(_00145_));
 sky130_fd_sc_hd__inv_2 _23131_ (.A(_10106_),
    .Y(_00146_));
 sky130_fd_sc_hd__inv_2 _23132_ (.A(_10106_),
    .Y(_00147_));
 sky130_fd_sc_hd__inv_2 _23133_ (.A(_10106_),
    .Y(_00148_));
 sky130_fd_sc_hd__inv_2 _23134_ (.A(_10106_),
    .Y(_00149_));
 sky130_fd_sc_hd__inv_2 _23135_ (.A(_10106_),
    .Y(_00150_));
 sky130_fd_sc_hd__inv_2 _23136_ (.A(_10106_),
    .Y(_00151_));
 sky130_fd_sc_hd__inv_2 _23137_ (.A(_10106_),
    .Y(_00152_));
 sky130_fd_sc_hd__inv_2 _23138_ (.A(_10106_),
    .Y(_00153_));
 sky130_fd_sc_hd__buf_1 _23139_ (.A(_10087_),
    .X(_10107_));
 sky130_fd_sc_hd__inv_2 _23140_ (.A(_10107_),
    .Y(_00154_));
 sky130_fd_sc_hd__inv_2 _23141_ (.A(_10107_),
    .Y(_00155_));
 sky130_fd_sc_hd__inv_2 _23142_ (.A(_10107_),
    .Y(_00156_));
 sky130_fd_sc_hd__inv_2 _23143_ (.A(_10107_),
    .Y(_00157_));
 sky130_fd_sc_hd__inv_2 _23144_ (.A(_10107_),
    .Y(_00158_));
 sky130_fd_sc_hd__inv_2 _23145_ (.A(_10107_),
    .Y(_00159_));
 sky130_fd_sc_hd__inv_2 _23146_ (.A(_10107_),
    .Y(_00160_));
 sky130_fd_sc_hd__inv_2 _23147_ (.A(_10107_),
    .Y(_00161_));
 sky130_fd_sc_hd__inv_2 _23148_ (.A(_10107_),
    .Y(_00162_));
 sky130_fd_sc_hd__inv_2 _23149_ (.A(_10107_),
    .Y(_00163_));
 sky130_fd_sc_hd__buf_1 _23150_ (.A(_10079_),
    .X(_10108_));
 sky130_fd_sc_hd__buf_1 _23151_ (.A(_10108_),
    .X(_10109_));
 sky130_fd_sc_hd__inv_2 _23152_ (.A(_10109_),
    .Y(_00164_));
 sky130_fd_sc_hd__inv_2 _23153_ (.A(_10109_),
    .Y(_00165_));
 sky130_fd_sc_hd__inv_2 _23154_ (.A(_10109_),
    .Y(_00166_));
 sky130_fd_sc_hd__inv_2 _23155_ (.A(_10109_),
    .Y(_00167_));
 sky130_fd_sc_hd__inv_2 _23156_ (.A(_10109_),
    .Y(_00168_));
 sky130_fd_sc_hd__inv_2 _23157_ (.A(_10109_),
    .Y(_00169_));
 sky130_fd_sc_hd__inv_2 _23158_ (.A(_10109_),
    .Y(_00170_));
 sky130_fd_sc_hd__inv_2 _23159_ (.A(_10109_),
    .Y(_00171_));
 sky130_fd_sc_hd__inv_2 _23160_ (.A(_10109_),
    .Y(_00172_));
 sky130_fd_sc_hd__inv_2 _23161_ (.A(_10109_),
    .Y(_00173_));
 sky130_fd_sc_hd__buf_1 _23162_ (.A(_10108_),
    .X(_10110_));
 sky130_fd_sc_hd__inv_2 _23163_ (.A(_10110_),
    .Y(_00174_));
 sky130_fd_sc_hd__inv_2 _23164_ (.A(_10110_),
    .Y(_00175_));
 sky130_fd_sc_hd__inv_2 _23165_ (.A(_10110_),
    .Y(_00176_));
 sky130_fd_sc_hd__inv_2 _23166_ (.A(_10110_),
    .Y(_00177_));
 sky130_fd_sc_hd__inv_2 _23167_ (.A(_10110_),
    .Y(_00178_));
 sky130_fd_sc_hd__inv_2 _23168_ (.A(_10110_),
    .Y(_00179_));
 sky130_fd_sc_hd__inv_2 _23169_ (.A(_10110_),
    .Y(_00180_));
 sky130_fd_sc_hd__inv_2 _23170_ (.A(_10110_),
    .Y(_00181_));
 sky130_fd_sc_hd__inv_2 _23171_ (.A(_10110_),
    .Y(_00182_));
 sky130_fd_sc_hd__inv_2 _23172_ (.A(_10110_),
    .Y(_00183_));
 sky130_fd_sc_hd__buf_1 _23173_ (.A(_10108_),
    .X(_10111_));
 sky130_fd_sc_hd__inv_2 _23174_ (.A(_10111_),
    .Y(_00184_));
 sky130_fd_sc_hd__inv_2 _23175_ (.A(_10111_),
    .Y(_00185_));
 sky130_fd_sc_hd__inv_2 _23176_ (.A(_10111_),
    .Y(_00186_));
 sky130_fd_sc_hd__inv_2 _23177_ (.A(_10111_),
    .Y(_00187_));
 sky130_fd_sc_hd__inv_2 _23178_ (.A(_10111_),
    .Y(_00188_));
 sky130_fd_sc_hd__inv_2 _23179_ (.A(_10111_),
    .Y(_00189_));
 sky130_fd_sc_hd__inv_2 _23180_ (.A(_10111_),
    .Y(_00190_));
 sky130_fd_sc_hd__inv_2 _23181_ (.A(_10111_),
    .Y(_00191_));
 sky130_fd_sc_hd__inv_2 _23182_ (.A(_10111_),
    .Y(_00192_));
 sky130_fd_sc_hd__inv_2 _23183_ (.A(_10111_),
    .Y(_00193_));
 sky130_fd_sc_hd__buf_1 _23184_ (.A(_10108_),
    .X(_10112_));
 sky130_fd_sc_hd__inv_2 _23185_ (.A(_10112_),
    .Y(_00194_));
 sky130_fd_sc_hd__inv_2 _23186_ (.A(_10112_),
    .Y(_00195_));
 sky130_fd_sc_hd__buf_8 _23187_ (.A(_07132_),
    .X(_10113_));
 sky130_fd_sc_hd__nor2_8 _23188_ (.A(_08144_),
    .B(net104),
    .Y(_10114_));
 sky130_fd_sc_hd__a21oi_4 _23189_ (.A1(_10113_),
    .A2(_10114_),
    .B1(_09361_),
    .Y(_10115_));
 sky130_fd_sc_hd__mux2_1 _23190_ (.A0(_09224_),
    .A1(\datamem.data_ram[5][16] ),
    .S(_10115_),
    .X(_10116_));
 sky130_fd_sc_hd__clkbuf_1 _23191_ (.A(_10116_),
    .X(_01364_));
 sky130_fd_sc_hd__mux2_1 _23192_ (.A0(_09236_),
    .A1(\datamem.data_ram[5][17] ),
    .S(_10115_),
    .X(_10117_));
 sky130_fd_sc_hd__clkbuf_1 _23193_ (.A(_10117_),
    .X(_01365_));
 sky130_fd_sc_hd__mux2_1 _23194_ (.A0(_09240_),
    .A1(\datamem.data_ram[5][18] ),
    .S(_10115_),
    .X(_10118_));
 sky130_fd_sc_hd__clkbuf_1 _23195_ (.A(_10118_),
    .X(_01366_));
 sky130_fd_sc_hd__mux2_1 _23196_ (.A0(_09244_),
    .A1(\datamem.data_ram[5][19] ),
    .S(_10115_),
    .X(_10119_));
 sky130_fd_sc_hd__clkbuf_1 _23197_ (.A(_10119_),
    .X(_01367_));
 sky130_fd_sc_hd__mux2_1 _23198_ (.A0(_09248_),
    .A1(\datamem.data_ram[5][20] ),
    .S(_10115_),
    .X(_10120_));
 sky130_fd_sc_hd__clkbuf_1 _23199_ (.A(_10120_),
    .X(_01368_));
 sky130_fd_sc_hd__mux2_1 _23200_ (.A0(_09252_),
    .A1(\datamem.data_ram[5][21] ),
    .S(_10115_),
    .X(_10121_));
 sky130_fd_sc_hd__clkbuf_1 _23201_ (.A(_10121_),
    .X(_01369_));
 sky130_fd_sc_hd__mux2_1 _23202_ (.A0(_09256_),
    .A1(\datamem.data_ram[5][22] ),
    .S(_10115_),
    .X(_10122_));
 sky130_fd_sc_hd__clkbuf_1 _23203_ (.A(_10122_),
    .X(_01370_));
 sky130_fd_sc_hd__mux2_1 _23204_ (.A0(_09260_),
    .A1(\datamem.data_ram[5][23] ),
    .S(_10115_),
    .X(_10123_));
 sky130_fd_sc_hd__clkbuf_1 _23205_ (.A(_10123_),
    .X(_01371_));
 sky130_fd_sc_hd__inv_2 _23206_ (.A(_10112_),
    .Y(_00196_));
 sky130_fd_sc_hd__inv_2 _23207_ (.A(_10112_),
    .Y(_00197_));
 sky130_fd_sc_hd__inv_2 _23208_ (.A(_10112_),
    .Y(_00198_));
 sky130_fd_sc_hd__inv_2 _23209_ (.A(_10112_),
    .Y(_00199_));
 sky130_fd_sc_hd__inv_2 _23210_ (.A(_10112_),
    .Y(_00200_));
 sky130_fd_sc_hd__inv_2 _23211_ (.A(_10112_),
    .Y(_00201_));
 sky130_fd_sc_hd__inv_2 _23212_ (.A(_10112_),
    .Y(_00202_));
 sky130_fd_sc_hd__inv_2 _23213_ (.A(_10112_),
    .Y(_00203_));
 sky130_fd_sc_hd__buf_1 _23214_ (.A(_10108_),
    .X(_10124_));
 sky130_fd_sc_hd__inv_2 _23215_ (.A(_10124_),
    .Y(_00204_));
 sky130_fd_sc_hd__inv_2 _23216_ (.A(_10124_),
    .Y(_00205_));
 sky130_fd_sc_hd__inv_2 _23217_ (.A(_10124_),
    .Y(_00206_));
 sky130_fd_sc_hd__inv_2 _23218_ (.A(_10124_),
    .Y(_00207_));
 sky130_fd_sc_hd__inv_2 _23219_ (.A(_10124_),
    .Y(_00208_));
 sky130_fd_sc_hd__inv_2 _23220_ (.A(_10124_),
    .Y(_00209_));
 sky130_fd_sc_hd__inv_2 _23221_ (.A(_10124_),
    .Y(_00210_));
 sky130_fd_sc_hd__inv_2 _23222_ (.A(_10124_),
    .Y(_00211_));
 sky130_fd_sc_hd__inv_2 _23223_ (.A(_10124_),
    .Y(_00212_));
 sky130_fd_sc_hd__inv_2 _23224_ (.A(_10124_),
    .Y(_00213_));
 sky130_fd_sc_hd__buf_1 _23225_ (.A(_10108_),
    .X(_10125_));
 sky130_fd_sc_hd__inv_2 _23226_ (.A(_10125_),
    .Y(_00214_));
 sky130_fd_sc_hd__inv_2 _23227_ (.A(_10125_),
    .Y(_00215_));
 sky130_fd_sc_hd__inv_2 _23228_ (.A(_10125_),
    .Y(_00216_));
 sky130_fd_sc_hd__inv_2 _23229_ (.A(_10125_),
    .Y(_00217_));
 sky130_fd_sc_hd__inv_2 _23230_ (.A(_10125_),
    .Y(_00218_));
 sky130_fd_sc_hd__inv_2 _23231_ (.A(_10125_),
    .Y(_00219_));
 sky130_fd_sc_hd__inv_2 _23232_ (.A(_10125_),
    .Y(_00220_));
 sky130_fd_sc_hd__inv_2 _23233_ (.A(_10125_),
    .Y(_00221_));
 sky130_fd_sc_hd__inv_2 _23234_ (.A(_10125_),
    .Y(_00222_));
 sky130_fd_sc_hd__inv_2 _23235_ (.A(_10125_),
    .Y(_00223_));
 sky130_fd_sc_hd__buf_1 _23236_ (.A(_10108_),
    .X(_10126_));
 sky130_fd_sc_hd__inv_2 _23237_ (.A(_10126_),
    .Y(_00224_));
 sky130_fd_sc_hd__inv_2 _23238_ (.A(_10126_),
    .Y(_00225_));
 sky130_fd_sc_hd__inv_2 _23239_ (.A(_10126_),
    .Y(_00226_));
 sky130_fd_sc_hd__inv_2 _23240_ (.A(_10126_),
    .Y(_00227_));
 sky130_fd_sc_hd__inv_2 _23241_ (.A(_10126_),
    .Y(_00228_));
 sky130_fd_sc_hd__inv_2 _23242_ (.A(_10126_),
    .Y(_00229_));
 sky130_fd_sc_hd__inv_2 _23243_ (.A(_10126_),
    .Y(_00230_));
 sky130_fd_sc_hd__inv_2 _23244_ (.A(_10126_),
    .Y(_00231_));
 sky130_fd_sc_hd__inv_2 _23245_ (.A(_10126_),
    .Y(_00232_));
 sky130_fd_sc_hd__inv_2 _23246_ (.A(_10126_),
    .Y(_00233_));
 sky130_fd_sc_hd__buf_1 _23247_ (.A(_10108_),
    .X(_10127_));
 sky130_fd_sc_hd__inv_2 _23248_ (.A(_10127_),
    .Y(_00234_));
 sky130_fd_sc_hd__inv_2 _23249_ (.A(_10127_),
    .Y(_00235_));
 sky130_fd_sc_hd__inv_2 _23250_ (.A(_10127_),
    .Y(_00236_));
 sky130_fd_sc_hd__inv_2 _23251_ (.A(_10127_),
    .Y(_00237_));
 sky130_fd_sc_hd__inv_2 _23252_ (.A(_10127_),
    .Y(_00238_));
 sky130_fd_sc_hd__inv_2 _23253_ (.A(_10127_),
    .Y(_00239_));
 sky130_fd_sc_hd__inv_2 _23254_ (.A(_10127_),
    .Y(_00240_));
 sky130_fd_sc_hd__inv_2 _23255_ (.A(_10127_),
    .Y(_00241_));
 sky130_fd_sc_hd__inv_2 _23256_ (.A(_10127_),
    .Y(_00242_));
 sky130_fd_sc_hd__inv_2 _23257_ (.A(_10127_),
    .Y(_00243_));
 sky130_fd_sc_hd__buf_1 _23258_ (.A(_10108_),
    .X(_10128_));
 sky130_fd_sc_hd__inv_2 _23259_ (.A(_10128_),
    .Y(_00244_));
 sky130_fd_sc_hd__inv_2 _23260_ (.A(_10128_),
    .Y(_00245_));
 sky130_fd_sc_hd__inv_2 _23261_ (.A(_10128_),
    .Y(_00246_));
 sky130_fd_sc_hd__inv_2 _23262_ (.A(_10128_),
    .Y(_00247_));
 sky130_fd_sc_hd__inv_2 _23263_ (.A(_10128_),
    .Y(_00248_));
 sky130_fd_sc_hd__inv_2 _23264_ (.A(_10128_),
    .Y(_00249_));
 sky130_fd_sc_hd__inv_2 _23265_ (.A(_10128_),
    .Y(_00250_));
 sky130_fd_sc_hd__inv_2 _23266_ (.A(_10128_),
    .Y(_00251_));
 sky130_fd_sc_hd__inv_2 _23267_ (.A(_10128_),
    .Y(_00252_));
 sky130_fd_sc_hd__inv_2 _23268_ (.A(_10128_),
    .Y(_00253_));
 sky130_fd_sc_hd__buf_1 _23269_ (.A(_10108_),
    .X(_10129_));
 sky130_fd_sc_hd__inv_2 _23270_ (.A(_10129_),
    .Y(_00254_));
 sky130_fd_sc_hd__inv_2 _23271_ (.A(_10129_),
    .Y(_00255_));
 sky130_fd_sc_hd__inv_2 _23272_ (.A(_10129_),
    .Y(_00256_));
 sky130_fd_sc_hd__inv_2 _23273_ (.A(_10129_),
    .Y(_00257_));
 sky130_fd_sc_hd__inv_2 _23274_ (.A(_10129_),
    .Y(_00258_));
 sky130_fd_sc_hd__inv_2 _23275_ (.A(_10129_),
    .Y(_00259_));
 sky130_fd_sc_hd__inv_2 _23276_ (.A(_10129_),
    .Y(_00260_));
 sky130_fd_sc_hd__inv_2 _23277_ (.A(_10129_),
    .Y(_00261_));
 sky130_fd_sc_hd__inv_2 _23278_ (.A(_10129_),
    .Y(_00262_));
 sky130_fd_sc_hd__inv_2 _23279_ (.A(_10129_),
    .Y(_00263_));
 sky130_fd_sc_hd__buf_1 _23280_ (.A(_10079_),
    .X(_10130_));
 sky130_fd_sc_hd__buf_1 _23281_ (.A(_10130_),
    .X(_10131_));
 sky130_fd_sc_hd__inv_2 _23282_ (.A(_10131_),
    .Y(_00264_));
 sky130_fd_sc_hd__inv_2 _23283_ (.A(_10131_),
    .Y(_00265_));
 sky130_fd_sc_hd__inv_2 _23284_ (.A(_10131_),
    .Y(_00266_));
 sky130_fd_sc_hd__inv_2 _23285_ (.A(_10131_),
    .Y(_00267_));
 sky130_fd_sc_hd__inv_2 _23286_ (.A(_10131_),
    .Y(_00268_));
 sky130_fd_sc_hd__inv_2 _23287_ (.A(_10131_),
    .Y(_00269_));
 sky130_fd_sc_hd__inv_2 _23288_ (.A(_10131_),
    .Y(_00270_));
 sky130_fd_sc_hd__inv_2 _23289_ (.A(_10131_),
    .Y(_00271_));
 sky130_fd_sc_hd__inv_2 _23290_ (.A(_10131_),
    .Y(_00272_));
 sky130_fd_sc_hd__inv_2 _23291_ (.A(_10131_),
    .Y(_00273_));
 sky130_fd_sc_hd__buf_1 _23292_ (.A(_10130_),
    .X(_10132_));
 sky130_fd_sc_hd__inv_2 _23293_ (.A(_10132_),
    .Y(_00274_));
 sky130_fd_sc_hd__inv_2 _23294_ (.A(_10132_),
    .Y(_00275_));
 sky130_fd_sc_hd__inv_2 _23295_ (.A(_10132_),
    .Y(_00276_));
 sky130_fd_sc_hd__inv_2 _23296_ (.A(_10132_),
    .Y(_00277_));
 sky130_fd_sc_hd__inv_2 _23297_ (.A(_10132_),
    .Y(_00278_));
 sky130_fd_sc_hd__inv_2 _23298_ (.A(_10132_),
    .Y(_00279_));
 sky130_fd_sc_hd__inv_2 _23299_ (.A(_10132_),
    .Y(_00280_));
 sky130_fd_sc_hd__inv_2 _23300_ (.A(_10132_),
    .Y(_00281_));
 sky130_fd_sc_hd__inv_2 _23301_ (.A(_10132_),
    .Y(_00282_));
 sky130_fd_sc_hd__inv_2 _23302_ (.A(_10132_),
    .Y(_00283_));
 sky130_fd_sc_hd__buf_1 _23303_ (.A(_10130_),
    .X(_10133_));
 sky130_fd_sc_hd__inv_2 _23304_ (.A(_10133_),
    .Y(_00284_));
 sky130_fd_sc_hd__inv_2 _23305_ (.A(_10133_),
    .Y(_00285_));
 sky130_fd_sc_hd__inv_2 _23306_ (.A(_10133_),
    .Y(_00286_));
 sky130_fd_sc_hd__inv_2 _23307_ (.A(_10133_),
    .Y(_00287_));
 sky130_fd_sc_hd__inv_2 _23308_ (.A(_10133_),
    .Y(_00288_));
 sky130_fd_sc_hd__inv_2 _23309_ (.A(_10133_),
    .Y(_00289_));
 sky130_fd_sc_hd__inv_2 _23310_ (.A(_10133_),
    .Y(_00290_));
 sky130_fd_sc_hd__inv_2 _23311_ (.A(_10133_),
    .Y(_00291_));
 sky130_fd_sc_hd__inv_2 _23312_ (.A(_10133_),
    .Y(_00292_));
 sky130_fd_sc_hd__inv_2 _23313_ (.A(_10133_),
    .Y(_00293_));
 sky130_fd_sc_hd__buf_1 _23314_ (.A(_10130_),
    .X(_10134_));
 sky130_fd_sc_hd__inv_2 _23315_ (.A(_10134_),
    .Y(_00294_));
 sky130_fd_sc_hd__inv_2 _23316_ (.A(_10134_),
    .Y(_00295_));
 sky130_fd_sc_hd__inv_2 _23317_ (.A(_10134_),
    .Y(_00296_));
 sky130_fd_sc_hd__inv_2 _23318_ (.A(_10134_),
    .Y(_00297_));
 sky130_fd_sc_hd__inv_2 _23319_ (.A(_10134_),
    .Y(_00298_));
 sky130_fd_sc_hd__inv_2 _23320_ (.A(_10134_),
    .Y(_00299_));
 sky130_fd_sc_hd__inv_2 _23321_ (.A(_10134_),
    .Y(_00300_));
 sky130_fd_sc_hd__inv_2 _23322_ (.A(_10134_),
    .Y(_00301_));
 sky130_fd_sc_hd__inv_2 _23323_ (.A(_10134_),
    .Y(_00302_));
 sky130_fd_sc_hd__inv_2 _23324_ (.A(_10134_),
    .Y(_00303_));
 sky130_fd_sc_hd__buf_1 _23325_ (.A(_10130_),
    .X(_10135_));
 sky130_fd_sc_hd__inv_2 _23326_ (.A(_10135_),
    .Y(_00304_));
 sky130_fd_sc_hd__inv_2 _23327_ (.A(_10135_),
    .Y(_00305_));
 sky130_fd_sc_hd__inv_2 _23328_ (.A(_10135_),
    .Y(_00306_));
 sky130_fd_sc_hd__inv_2 _23329_ (.A(_10135_),
    .Y(_00307_));
 sky130_fd_sc_hd__inv_2 _23330_ (.A(_10135_),
    .Y(_00308_));
 sky130_fd_sc_hd__inv_2 _23331_ (.A(_10135_),
    .Y(_00309_));
 sky130_fd_sc_hd__inv_2 _23332_ (.A(_10135_),
    .Y(_00310_));
 sky130_fd_sc_hd__inv_2 _23333_ (.A(_10135_),
    .Y(_00311_));
 sky130_fd_sc_hd__inv_2 _23334_ (.A(_10135_),
    .Y(_00312_));
 sky130_fd_sc_hd__inv_2 _23335_ (.A(_10135_),
    .Y(_00313_));
 sky130_fd_sc_hd__buf_1 _23336_ (.A(_10130_),
    .X(_10136_));
 sky130_fd_sc_hd__inv_2 _23337_ (.A(_10136_),
    .Y(_00314_));
 sky130_fd_sc_hd__inv_2 _23338_ (.A(_10136_),
    .Y(_00315_));
 sky130_fd_sc_hd__inv_2 _23339_ (.A(_10136_),
    .Y(_00316_));
 sky130_fd_sc_hd__inv_2 _23340_ (.A(_10136_),
    .Y(_00317_));
 sky130_fd_sc_hd__inv_2 _23341_ (.A(_10136_),
    .Y(_00318_));
 sky130_fd_sc_hd__inv_2 _23342_ (.A(_10136_),
    .Y(_00319_));
 sky130_fd_sc_hd__inv_2 _23343_ (.A(_10136_),
    .Y(_00320_));
 sky130_fd_sc_hd__inv_2 _23344_ (.A(_10136_),
    .Y(_00321_));
 sky130_fd_sc_hd__inv_2 _23345_ (.A(_10136_),
    .Y(_00322_));
 sky130_fd_sc_hd__inv_2 _23346_ (.A(_10136_),
    .Y(_00323_));
 sky130_fd_sc_hd__buf_1 _23347_ (.A(_10130_),
    .X(_10137_));
 sky130_fd_sc_hd__inv_2 _23348_ (.A(_10137_),
    .Y(_00324_));
 sky130_fd_sc_hd__inv_2 _23349_ (.A(_10137_),
    .Y(_00325_));
 sky130_fd_sc_hd__inv_2 _23350_ (.A(_10137_),
    .Y(_00326_));
 sky130_fd_sc_hd__inv_2 _23351_ (.A(_10137_),
    .Y(_00327_));
 sky130_fd_sc_hd__inv_2 _23352_ (.A(_10137_),
    .Y(_00328_));
 sky130_fd_sc_hd__inv_2 _23353_ (.A(_10137_),
    .Y(_00329_));
 sky130_fd_sc_hd__inv_2 _23354_ (.A(_10137_),
    .Y(_00330_));
 sky130_fd_sc_hd__inv_2 _23355_ (.A(_10137_),
    .Y(_00331_));
 sky130_fd_sc_hd__inv_2 _23356_ (.A(_10137_),
    .Y(_00332_));
 sky130_fd_sc_hd__inv_2 _23357_ (.A(_10137_),
    .Y(_00333_));
 sky130_fd_sc_hd__buf_1 _23358_ (.A(_10130_),
    .X(_10138_));
 sky130_fd_sc_hd__inv_2 _23359_ (.A(_10138_),
    .Y(_00334_));
 sky130_fd_sc_hd__inv_2 _23360_ (.A(_10138_),
    .Y(_00335_));
 sky130_fd_sc_hd__inv_2 _23361_ (.A(_10138_),
    .Y(_00336_));
 sky130_fd_sc_hd__inv_2 _23362_ (.A(_10138_),
    .Y(_00337_));
 sky130_fd_sc_hd__inv_2 _23363_ (.A(_10138_),
    .Y(_00338_));
 sky130_fd_sc_hd__inv_2 _23364_ (.A(_10138_),
    .Y(_00339_));
 sky130_fd_sc_hd__inv_2 _23365_ (.A(_10138_),
    .Y(_00340_));
 sky130_fd_sc_hd__inv_2 _23366_ (.A(_10138_),
    .Y(_00341_));
 sky130_fd_sc_hd__inv_2 _23367_ (.A(_10138_),
    .Y(_00342_));
 sky130_fd_sc_hd__inv_2 _23368_ (.A(_10138_),
    .Y(_00343_));
 sky130_fd_sc_hd__buf_1 _23369_ (.A(_10130_),
    .X(_10139_));
 sky130_fd_sc_hd__inv_2 _23370_ (.A(_10139_),
    .Y(_00344_));
 sky130_fd_sc_hd__inv_2 _23371_ (.A(_10139_),
    .Y(_00345_));
 sky130_fd_sc_hd__inv_2 _23372_ (.A(_10139_),
    .Y(_00346_));
 sky130_fd_sc_hd__inv_2 _23373_ (.A(_10139_),
    .Y(_00347_));
 sky130_fd_sc_hd__inv_2 _23374_ (.A(_10139_),
    .Y(_00348_));
 sky130_fd_sc_hd__inv_2 _23375_ (.A(_10139_),
    .Y(_00349_));
 sky130_fd_sc_hd__inv_2 _23376_ (.A(_10139_),
    .Y(_00350_));
 sky130_fd_sc_hd__inv_2 _23377_ (.A(_10139_),
    .Y(_00351_));
 sky130_fd_sc_hd__inv_2 _23378_ (.A(_10139_),
    .Y(_00352_));
 sky130_fd_sc_hd__inv_2 _23379_ (.A(_10139_),
    .Y(_00353_));
 sky130_fd_sc_hd__buf_1 _23380_ (.A(_10130_),
    .X(_10140_));
 sky130_fd_sc_hd__inv_2 _23381_ (.A(_10140_),
    .Y(_00354_));
 sky130_fd_sc_hd__inv_2 _23382_ (.A(_10140_),
    .Y(_00355_));
 sky130_fd_sc_hd__buf_12 _23383_ (.A(_07137_),
    .X(_10141_));
 sky130_fd_sc_hd__buf_8 _23384_ (.A(_10141_),
    .X(_10142_));
 sky130_fd_sc_hd__a21oi_4 _23385_ (.A1(_10142_),
    .A2(_09301_),
    .B1(_09361_),
    .Y(_10143_));
 sky130_fd_sc_hd__mux2_1 _23386_ (.A0(_09298_),
    .A1(\datamem.data_ram[59][24] ),
    .S(_10143_),
    .X(_10144_));
 sky130_fd_sc_hd__clkbuf_1 _23387_ (.A(_10144_),
    .X(_01532_));
 sky130_fd_sc_hd__mux2_1 _23388_ (.A0(_09306_),
    .A1(\datamem.data_ram[59][25] ),
    .S(_10143_),
    .X(_10145_));
 sky130_fd_sc_hd__clkbuf_1 _23389_ (.A(_10145_),
    .X(_01533_));
 sky130_fd_sc_hd__mux2_1 _23390_ (.A0(_09310_),
    .A1(\datamem.data_ram[59][26] ),
    .S(_10143_),
    .X(_10146_));
 sky130_fd_sc_hd__clkbuf_1 _23391_ (.A(_10146_),
    .X(_01534_));
 sky130_fd_sc_hd__mux2_1 _23392_ (.A0(_09314_),
    .A1(\datamem.data_ram[59][27] ),
    .S(_10143_),
    .X(_10147_));
 sky130_fd_sc_hd__clkbuf_1 _23393_ (.A(_10147_),
    .X(_01535_));
 sky130_fd_sc_hd__mux2_1 _23394_ (.A0(_09318_),
    .A1(\datamem.data_ram[59][28] ),
    .S(_10143_),
    .X(_10148_));
 sky130_fd_sc_hd__clkbuf_1 _23395_ (.A(_10148_),
    .X(_01536_));
 sky130_fd_sc_hd__mux2_1 _23396_ (.A0(_09322_),
    .A1(\datamem.data_ram[59][29] ),
    .S(_10143_),
    .X(_10149_));
 sky130_fd_sc_hd__clkbuf_1 _23397_ (.A(_10149_),
    .X(_01537_));
 sky130_fd_sc_hd__mux2_1 _23398_ (.A0(_09326_),
    .A1(\datamem.data_ram[59][30] ),
    .S(_10143_),
    .X(_10150_));
 sky130_fd_sc_hd__clkbuf_1 _23399_ (.A(_10150_),
    .X(_01538_));
 sky130_fd_sc_hd__mux2_1 _23400_ (.A0(_09330_),
    .A1(\datamem.data_ram[59][31] ),
    .S(_10143_),
    .X(_10151_));
 sky130_fd_sc_hd__clkbuf_1 _23401_ (.A(_10151_),
    .X(_01539_));
 sky130_fd_sc_hd__inv_2 _23402_ (.A(_10140_),
    .Y(_00356_));
 sky130_fd_sc_hd__inv_2 _23403_ (.A(_10140_),
    .Y(_00357_));
 sky130_fd_sc_hd__inv_2 _23404_ (.A(_10140_),
    .Y(_00358_));
 sky130_fd_sc_hd__inv_2 _23405_ (.A(_10140_),
    .Y(_00359_));
 sky130_fd_sc_hd__inv_2 _23406_ (.A(_10140_),
    .Y(_00360_));
 sky130_fd_sc_hd__inv_2 _23407_ (.A(_10140_),
    .Y(_00361_));
 sky130_fd_sc_hd__inv_2 _23408_ (.A(_10140_),
    .Y(_00362_));
 sky130_fd_sc_hd__inv_2 _23409_ (.A(_10140_),
    .Y(_00363_));
 sky130_fd_sc_hd__buf_1 _23410_ (.A(_10078_),
    .X(_10152_));
 sky130_fd_sc_hd__buf_1 _23411_ (.A(_10152_),
    .X(_10153_));
 sky130_fd_sc_hd__inv_2 _23412_ (.A(_10153_),
    .Y(_00364_));
 sky130_fd_sc_hd__inv_2 _23413_ (.A(_10153_),
    .Y(_00365_));
 sky130_fd_sc_hd__inv_2 _23414_ (.A(_10153_),
    .Y(_00366_));
 sky130_fd_sc_hd__inv_2 _23415_ (.A(_10153_),
    .Y(_00367_));
 sky130_fd_sc_hd__inv_2 _23416_ (.A(_10153_),
    .Y(_00368_));
 sky130_fd_sc_hd__inv_2 _23417_ (.A(_10153_),
    .Y(_00369_));
 sky130_fd_sc_hd__inv_2 _23418_ (.A(_10153_),
    .Y(_00370_));
 sky130_fd_sc_hd__inv_2 _23419_ (.A(_10153_),
    .Y(_00371_));
 sky130_fd_sc_hd__inv_2 _23420_ (.A(_10153_),
    .Y(_00372_));
 sky130_fd_sc_hd__inv_2 _23421_ (.A(_10153_),
    .Y(_00373_));
 sky130_fd_sc_hd__buf_1 _23422_ (.A(_10152_),
    .X(_10154_));
 sky130_fd_sc_hd__inv_2 _23423_ (.A(_10154_),
    .Y(_00374_));
 sky130_fd_sc_hd__inv_2 _23424_ (.A(_10154_),
    .Y(_00375_));
 sky130_fd_sc_hd__inv_2 _23425_ (.A(_10154_),
    .Y(_00376_));
 sky130_fd_sc_hd__inv_2 _23426_ (.A(_10154_),
    .Y(_00377_));
 sky130_fd_sc_hd__inv_2 _23427_ (.A(_10154_),
    .Y(_00378_));
 sky130_fd_sc_hd__inv_2 _23428_ (.A(_10154_),
    .Y(_00379_));
 sky130_fd_sc_hd__inv_2 _23429_ (.A(_10154_),
    .Y(_00380_));
 sky130_fd_sc_hd__inv_2 _23430_ (.A(_10154_),
    .Y(_00381_));
 sky130_fd_sc_hd__inv_2 _23431_ (.A(_10154_),
    .Y(_00382_));
 sky130_fd_sc_hd__inv_2 _23432_ (.A(_10154_),
    .Y(_00383_));
 sky130_fd_sc_hd__buf_1 _23433_ (.A(_10152_),
    .X(_10155_));
 sky130_fd_sc_hd__inv_2 _23434_ (.A(_10155_),
    .Y(_00384_));
 sky130_fd_sc_hd__inv_2 _23435_ (.A(_10155_),
    .Y(_00385_));
 sky130_fd_sc_hd__inv_2 _23436_ (.A(_10155_),
    .Y(_00386_));
 sky130_fd_sc_hd__inv_2 _23437_ (.A(_10155_),
    .Y(_00387_));
 sky130_fd_sc_hd__inv_2 _23438_ (.A(_10155_),
    .Y(_00388_));
 sky130_fd_sc_hd__inv_2 _23439_ (.A(_10155_),
    .Y(_00389_));
 sky130_fd_sc_hd__inv_2 _23440_ (.A(_10155_),
    .Y(_00390_));
 sky130_fd_sc_hd__inv_2 _23441_ (.A(_10155_),
    .Y(_00391_));
 sky130_fd_sc_hd__inv_2 _23442_ (.A(_10155_),
    .Y(_00392_));
 sky130_fd_sc_hd__inv_2 _23443_ (.A(_10155_),
    .Y(_00393_));
 sky130_fd_sc_hd__buf_1 _23444_ (.A(_10152_),
    .X(_10156_));
 sky130_fd_sc_hd__inv_2 _23445_ (.A(_10156_),
    .Y(_00394_));
 sky130_fd_sc_hd__inv_2 _23446_ (.A(_10156_),
    .Y(_00395_));
 sky130_fd_sc_hd__inv_2 _23447_ (.A(_10156_),
    .Y(_00396_));
 sky130_fd_sc_hd__inv_2 _23448_ (.A(_10156_),
    .Y(_00397_));
 sky130_fd_sc_hd__inv_2 _23449_ (.A(_10156_),
    .Y(_00398_));
 sky130_fd_sc_hd__inv_2 _23450_ (.A(_10156_),
    .Y(_00399_));
 sky130_fd_sc_hd__inv_2 _23451_ (.A(_10156_),
    .Y(_00400_));
 sky130_fd_sc_hd__inv_2 _23452_ (.A(_10156_),
    .Y(_00401_));
 sky130_fd_sc_hd__inv_2 _23453_ (.A(_10156_),
    .Y(_00402_));
 sky130_fd_sc_hd__inv_2 _23454_ (.A(_10156_),
    .Y(_00403_));
 sky130_fd_sc_hd__buf_1 _23455_ (.A(_10152_),
    .X(_10157_));
 sky130_fd_sc_hd__inv_2 _23456_ (.A(_10157_),
    .Y(_00404_));
 sky130_fd_sc_hd__inv_2 _23457_ (.A(_10157_),
    .Y(_00405_));
 sky130_fd_sc_hd__inv_2 _23458_ (.A(_10157_),
    .Y(_00406_));
 sky130_fd_sc_hd__inv_2 _23459_ (.A(_10157_),
    .Y(_00407_));
 sky130_fd_sc_hd__inv_2 _23460_ (.A(_10157_),
    .Y(_00408_));
 sky130_fd_sc_hd__inv_2 _23461_ (.A(_10157_),
    .Y(_00409_));
 sky130_fd_sc_hd__inv_2 _23462_ (.A(_10157_),
    .Y(_00410_));
 sky130_fd_sc_hd__inv_2 _23463_ (.A(_10157_),
    .Y(_00411_));
 sky130_fd_sc_hd__inv_2 _23464_ (.A(_10157_),
    .Y(_00412_));
 sky130_fd_sc_hd__inv_2 _23465_ (.A(_10157_),
    .Y(_00413_));
 sky130_fd_sc_hd__buf_1 _23466_ (.A(_10152_),
    .X(_10158_));
 sky130_fd_sc_hd__inv_2 _23467_ (.A(_10158_),
    .Y(_00414_));
 sky130_fd_sc_hd__inv_2 _23468_ (.A(_10158_),
    .Y(_00415_));
 sky130_fd_sc_hd__inv_2 _23469_ (.A(_10158_),
    .Y(_00416_));
 sky130_fd_sc_hd__inv_2 _23470_ (.A(_10158_),
    .Y(_00417_));
 sky130_fd_sc_hd__inv_2 _23471_ (.A(_10158_),
    .Y(_00418_));
 sky130_fd_sc_hd__inv_2 _23472_ (.A(_10158_),
    .Y(_00419_));
 sky130_fd_sc_hd__inv_2 _23473_ (.A(_10158_),
    .Y(_00420_));
 sky130_fd_sc_hd__inv_2 _23474_ (.A(_10158_),
    .Y(_00421_));
 sky130_fd_sc_hd__inv_2 _23475_ (.A(_10158_),
    .Y(_00422_));
 sky130_fd_sc_hd__inv_2 _23476_ (.A(_10158_),
    .Y(_00423_));
 sky130_fd_sc_hd__buf_1 _23477_ (.A(_10152_),
    .X(_10159_));
 sky130_fd_sc_hd__inv_2 _23478_ (.A(_10159_),
    .Y(_00424_));
 sky130_fd_sc_hd__inv_2 _23479_ (.A(_10159_),
    .Y(_00425_));
 sky130_fd_sc_hd__inv_2 _23480_ (.A(_10159_),
    .Y(_00426_));
 sky130_fd_sc_hd__inv_2 _23481_ (.A(_10159_),
    .Y(_00427_));
 sky130_fd_sc_hd__inv_2 _23482_ (.A(_10159_),
    .Y(_00428_));
 sky130_fd_sc_hd__inv_2 _23483_ (.A(_10159_),
    .Y(_00429_));
 sky130_fd_sc_hd__inv_2 _23484_ (.A(_10159_),
    .Y(_00430_));
 sky130_fd_sc_hd__inv_2 _23485_ (.A(_10159_),
    .Y(_00431_));
 sky130_fd_sc_hd__inv_2 _23486_ (.A(_10159_),
    .Y(_00432_));
 sky130_fd_sc_hd__inv_2 _23487_ (.A(_10159_),
    .Y(_00433_));
 sky130_fd_sc_hd__buf_1 _23488_ (.A(_10152_),
    .X(_10160_));
 sky130_fd_sc_hd__inv_2 _23489_ (.A(_10160_),
    .Y(_00434_));
 sky130_fd_sc_hd__inv_2 _23490_ (.A(_10160_),
    .Y(_00435_));
 sky130_fd_sc_hd__inv_2 _23491_ (.A(_10160_),
    .Y(_00436_));
 sky130_fd_sc_hd__inv_2 _23492_ (.A(_10160_),
    .Y(_00437_));
 sky130_fd_sc_hd__inv_2 _23493_ (.A(_10160_),
    .Y(_00438_));
 sky130_fd_sc_hd__inv_2 _23494_ (.A(_10160_),
    .Y(_00439_));
 sky130_fd_sc_hd__inv_2 _23495_ (.A(_10160_),
    .Y(_00440_));
 sky130_fd_sc_hd__inv_2 _23496_ (.A(_10160_),
    .Y(_00441_));
 sky130_fd_sc_hd__inv_2 _23497_ (.A(_10160_),
    .Y(_00442_));
 sky130_fd_sc_hd__inv_2 _23498_ (.A(_10160_),
    .Y(_00443_));
 sky130_fd_sc_hd__buf_1 _23499_ (.A(_10152_),
    .X(_10161_));
 sky130_fd_sc_hd__inv_2 _23500_ (.A(_10161_),
    .Y(_00444_));
 sky130_fd_sc_hd__inv_2 _23501_ (.A(_10161_),
    .Y(_00445_));
 sky130_fd_sc_hd__inv_2 _23502_ (.A(_10161_),
    .Y(_00446_));
 sky130_fd_sc_hd__inv_2 _23503_ (.A(_10161_),
    .Y(_00447_));
 sky130_fd_sc_hd__inv_2 _23504_ (.A(_10161_),
    .Y(_00448_));
 sky130_fd_sc_hd__inv_2 _23505_ (.A(_10161_),
    .Y(_00449_));
 sky130_fd_sc_hd__inv_2 _23506_ (.A(_10161_),
    .Y(_00450_));
 sky130_fd_sc_hd__inv_2 _23507_ (.A(_10161_),
    .Y(_00451_));
 sky130_fd_sc_hd__a21oi_4 _23508_ (.A1(_10142_),
    .A2(_09229_),
    .B1(_09361_),
    .Y(_10162_));
 sky130_fd_sc_hd__mux2_1 _23509_ (.A0(_09224_),
    .A1(\datamem.data_ram[59][16] ),
    .S(_10162_),
    .X(_10163_));
 sky130_fd_sc_hd__clkbuf_1 _23510_ (.A(_10163_),
    .X(_01636_));
 sky130_fd_sc_hd__mux2_1 _23511_ (.A0(_09236_),
    .A1(\datamem.data_ram[59][17] ),
    .S(_10162_),
    .X(_10164_));
 sky130_fd_sc_hd__clkbuf_1 _23512_ (.A(_10164_),
    .X(_01637_));
 sky130_fd_sc_hd__mux2_1 _23513_ (.A0(_09240_),
    .A1(\datamem.data_ram[59][18] ),
    .S(_10162_),
    .X(_10165_));
 sky130_fd_sc_hd__clkbuf_1 _23514_ (.A(_10165_),
    .X(_01638_));
 sky130_fd_sc_hd__mux2_1 _23515_ (.A0(_09244_),
    .A1(\datamem.data_ram[59][19] ),
    .S(_10162_),
    .X(_10166_));
 sky130_fd_sc_hd__clkbuf_1 _23516_ (.A(_10166_),
    .X(_01639_));
 sky130_fd_sc_hd__mux2_1 _23517_ (.A0(_09248_),
    .A1(\datamem.data_ram[59][20] ),
    .S(_10162_),
    .X(_10167_));
 sky130_fd_sc_hd__clkbuf_1 _23518_ (.A(_10167_),
    .X(_01640_));
 sky130_fd_sc_hd__mux2_1 _23519_ (.A0(_09252_),
    .A1(\datamem.data_ram[59][21] ),
    .S(_10162_),
    .X(_10168_));
 sky130_fd_sc_hd__clkbuf_1 _23520_ (.A(_10168_),
    .X(_01641_));
 sky130_fd_sc_hd__mux2_1 _23521_ (.A0(_09256_),
    .A1(\datamem.data_ram[59][22] ),
    .S(_10162_),
    .X(_10169_));
 sky130_fd_sc_hd__clkbuf_1 _23522_ (.A(_10169_),
    .X(_01642_));
 sky130_fd_sc_hd__mux2_1 _23523_ (.A0(_09260_),
    .A1(\datamem.data_ram[59][23] ),
    .S(_10162_),
    .X(_10170_));
 sky130_fd_sc_hd__clkbuf_1 _23524_ (.A(_10170_),
    .X(_01643_));
 sky130_fd_sc_hd__inv_2 _23525_ (.A(_10161_),
    .Y(_00452_));
 sky130_fd_sc_hd__inv_2 _23526_ (.A(_10161_),
    .Y(_00453_));
 sky130_fd_sc_hd__buf_1 _23527_ (.A(_10152_),
    .X(_10171_));
 sky130_fd_sc_hd__inv_2 _23528_ (.A(_10171_),
    .Y(_00454_));
 sky130_fd_sc_hd__inv_2 _23529_ (.A(_10171_),
    .Y(_00455_));
 sky130_fd_sc_hd__inv_2 _23530_ (.A(_10171_),
    .Y(_00456_));
 sky130_fd_sc_hd__inv_2 _23531_ (.A(_10171_),
    .Y(_00457_));
 sky130_fd_sc_hd__inv_2 _23532_ (.A(_10171_),
    .Y(_00458_));
 sky130_fd_sc_hd__inv_2 _23533_ (.A(_10171_),
    .Y(_00459_));
 sky130_fd_sc_hd__inv_2 _23534_ (.A(_10171_),
    .Y(_00460_));
 sky130_fd_sc_hd__inv_2 _23535_ (.A(_10171_),
    .Y(_00461_));
 sky130_fd_sc_hd__inv_2 _23536_ (.A(_10171_),
    .Y(_00462_));
 sky130_fd_sc_hd__inv_2 _23537_ (.A(_10171_),
    .Y(_00463_));
 sky130_fd_sc_hd__buf_1 _23538_ (.A(_10078_),
    .X(_10172_));
 sky130_fd_sc_hd__buf_1 _23539_ (.A(_10172_),
    .X(_10173_));
 sky130_fd_sc_hd__inv_2 _23540_ (.A(_10173_),
    .Y(_00464_));
 sky130_fd_sc_hd__inv_2 _23541_ (.A(_10173_),
    .Y(_00465_));
 sky130_fd_sc_hd__inv_2 _23542_ (.A(_10173_),
    .Y(_00466_));
 sky130_fd_sc_hd__inv_2 _23543_ (.A(_10173_),
    .Y(_00467_));
 sky130_fd_sc_hd__inv_2 _23544_ (.A(_10173_),
    .Y(_00468_));
 sky130_fd_sc_hd__inv_2 _23545_ (.A(_10173_),
    .Y(_00469_));
 sky130_fd_sc_hd__inv_2 _23546_ (.A(_10173_),
    .Y(_00470_));
 sky130_fd_sc_hd__inv_2 _23547_ (.A(_10173_),
    .Y(_00471_));
 sky130_fd_sc_hd__inv_2 _23548_ (.A(_10173_),
    .Y(_00472_));
 sky130_fd_sc_hd__inv_2 _23549_ (.A(_10173_),
    .Y(_00473_));
 sky130_fd_sc_hd__buf_1 _23550_ (.A(_10172_),
    .X(_10174_));
 sky130_fd_sc_hd__inv_2 _23551_ (.A(_10174_),
    .Y(_00474_));
 sky130_fd_sc_hd__inv_2 _23552_ (.A(_10174_),
    .Y(_00475_));
 sky130_fd_sc_hd__inv_2 _23553_ (.A(_10174_),
    .Y(_00476_));
 sky130_fd_sc_hd__inv_2 _23554_ (.A(_10174_),
    .Y(_00477_));
 sky130_fd_sc_hd__inv_2 _23555_ (.A(_10174_),
    .Y(_00478_));
 sky130_fd_sc_hd__inv_2 _23556_ (.A(_10174_),
    .Y(_00479_));
 sky130_fd_sc_hd__inv_2 _23557_ (.A(_10174_),
    .Y(_00480_));
 sky130_fd_sc_hd__inv_2 _23558_ (.A(_10174_),
    .Y(_00481_));
 sky130_fd_sc_hd__inv_2 _23559_ (.A(_10174_),
    .Y(_00482_));
 sky130_fd_sc_hd__inv_2 _23560_ (.A(_10174_),
    .Y(_00483_));
 sky130_fd_sc_hd__buf_1 _23561_ (.A(_10172_),
    .X(_10175_));
 sky130_fd_sc_hd__inv_2 _23562_ (.A(_10175_),
    .Y(_00484_));
 sky130_fd_sc_hd__inv_2 _23563_ (.A(_10175_),
    .Y(_00485_));
 sky130_fd_sc_hd__inv_2 _23564_ (.A(_10175_),
    .Y(_00486_));
 sky130_fd_sc_hd__inv_2 _23565_ (.A(_10175_),
    .Y(_00487_));
 sky130_fd_sc_hd__inv_2 _23566_ (.A(_10175_),
    .Y(_00488_));
 sky130_fd_sc_hd__inv_2 _23567_ (.A(_10175_),
    .Y(_00489_));
 sky130_fd_sc_hd__inv_2 _23568_ (.A(_10175_),
    .Y(_00490_));
 sky130_fd_sc_hd__inv_2 _23569_ (.A(_10175_),
    .Y(_00491_));
 sky130_fd_sc_hd__inv_2 _23570_ (.A(_10175_),
    .Y(_00492_));
 sky130_fd_sc_hd__inv_2 _23571_ (.A(_10175_),
    .Y(_00493_));
 sky130_fd_sc_hd__buf_1 _23572_ (.A(_10172_),
    .X(_10176_));
 sky130_fd_sc_hd__inv_2 _23573_ (.A(_10176_),
    .Y(_00494_));
 sky130_fd_sc_hd__inv_2 _23574_ (.A(_10176_),
    .Y(_00495_));
 sky130_fd_sc_hd__inv_2 _23575_ (.A(_10176_),
    .Y(_00496_));
 sky130_fd_sc_hd__inv_2 _23576_ (.A(_10176_),
    .Y(_00497_));
 sky130_fd_sc_hd__inv_2 _23577_ (.A(_10176_),
    .Y(_00498_));
 sky130_fd_sc_hd__inv_2 _23578_ (.A(_10176_),
    .Y(_00499_));
 sky130_fd_sc_hd__inv_2 _23579_ (.A(_10176_),
    .Y(_00500_));
 sky130_fd_sc_hd__inv_2 _23580_ (.A(_10176_),
    .Y(_00501_));
 sky130_fd_sc_hd__inv_2 _23581_ (.A(_10176_),
    .Y(_00502_));
 sky130_fd_sc_hd__inv_2 _23582_ (.A(_10176_),
    .Y(_00503_));
 sky130_fd_sc_hd__buf_1 _23583_ (.A(_10172_),
    .X(_10177_));
 sky130_fd_sc_hd__inv_2 _23584_ (.A(_10177_),
    .Y(_00504_));
 sky130_fd_sc_hd__inv_2 _23585_ (.A(_10177_),
    .Y(_00505_));
 sky130_fd_sc_hd__inv_2 _23586_ (.A(_10177_),
    .Y(_00506_));
 sky130_fd_sc_hd__inv_2 _23587_ (.A(_10177_),
    .Y(_00507_));
 sky130_fd_sc_hd__inv_2 _23588_ (.A(_10177_),
    .Y(_00508_));
 sky130_fd_sc_hd__inv_2 _23589_ (.A(_10177_),
    .Y(_00509_));
 sky130_fd_sc_hd__inv_2 _23590_ (.A(_10177_),
    .Y(_00510_));
 sky130_fd_sc_hd__inv_2 _23591_ (.A(_10177_),
    .Y(_00511_));
 sky130_fd_sc_hd__inv_2 _23592_ (.A(_10177_),
    .Y(_00512_));
 sky130_fd_sc_hd__inv_2 _23593_ (.A(_10177_),
    .Y(_00513_));
 sky130_fd_sc_hd__buf_1 _23594_ (.A(_10172_),
    .X(_10178_));
 sky130_fd_sc_hd__inv_2 _23595_ (.A(_10178_),
    .Y(_00514_));
 sky130_fd_sc_hd__inv_2 _23596_ (.A(_10178_),
    .Y(_00515_));
 sky130_fd_sc_hd__inv_2 _23597_ (.A(_10178_),
    .Y(_00516_));
 sky130_fd_sc_hd__inv_2 _23598_ (.A(_10178_),
    .Y(_00517_));
 sky130_fd_sc_hd__inv_2 _23599_ (.A(_10178_),
    .Y(_00518_));
 sky130_fd_sc_hd__inv_2 _23600_ (.A(_10178_),
    .Y(_00519_));
 sky130_fd_sc_hd__inv_2 _23601_ (.A(_10178_),
    .Y(_00520_));
 sky130_fd_sc_hd__inv_2 _23602_ (.A(_10178_),
    .Y(_00521_));
 sky130_fd_sc_hd__inv_2 _23603_ (.A(_10178_),
    .Y(_00522_));
 sky130_fd_sc_hd__inv_2 _23604_ (.A(_10178_),
    .Y(_00523_));
 sky130_fd_sc_hd__buf_1 _23605_ (.A(_10172_),
    .X(_10179_));
 sky130_fd_sc_hd__inv_2 _23606_ (.A(_10179_),
    .Y(_00524_));
 sky130_fd_sc_hd__inv_2 _23607_ (.A(_10179_),
    .Y(_00525_));
 sky130_fd_sc_hd__inv_2 _23608_ (.A(_10179_),
    .Y(_00526_));
 sky130_fd_sc_hd__inv_2 _23609_ (.A(_10179_),
    .Y(_00527_));
 sky130_fd_sc_hd__inv_2 _23610_ (.A(_10179_),
    .Y(_00528_));
 sky130_fd_sc_hd__inv_2 _23611_ (.A(_10179_),
    .Y(_00529_));
 sky130_fd_sc_hd__inv_2 _23612_ (.A(_10179_),
    .Y(_00530_));
 sky130_fd_sc_hd__inv_2 _23613_ (.A(_10179_),
    .Y(_00531_));
 sky130_fd_sc_hd__inv_2 _23614_ (.A(_10179_),
    .Y(_00532_));
 sky130_fd_sc_hd__inv_2 _23615_ (.A(_10179_),
    .Y(_00533_));
 sky130_fd_sc_hd__buf_1 _23616_ (.A(_10172_),
    .X(_10180_));
 sky130_fd_sc_hd__inv_2 _23617_ (.A(_10180_),
    .Y(_00534_));
 sky130_fd_sc_hd__inv_2 _23618_ (.A(_10180_),
    .Y(_00535_));
 sky130_fd_sc_hd__inv_2 _23619_ (.A(_10180_),
    .Y(_00536_));
 sky130_fd_sc_hd__inv_2 _23620_ (.A(_10180_),
    .Y(_00537_));
 sky130_fd_sc_hd__inv_2 _23621_ (.A(_10180_),
    .Y(_00538_));
 sky130_fd_sc_hd__inv_2 _23622_ (.A(_10180_),
    .Y(_00539_));
 sky130_fd_sc_hd__inv_2 _23623_ (.A(_10180_),
    .Y(_00540_));
 sky130_fd_sc_hd__inv_2 _23624_ (.A(_10180_),
    .Y(_00541_));
 sky130_fd_sc_hd__inv_2 _23625_ (.A(_10180_),
    .Y(_00542_));
 sky130_fd_sc_hd__inv_2 _23626_ (.A(_10180_),
    .Y(_00543_));
 sky130_fd_sc_hd__buf_1 _23627_ (.A(_10172_),
    .X(_10181_));
 sky130_fd_sc_hd__inv_2 _23628_ (.A(_10181_),
    .Y(_00544_));
 sky130_fd_sc_hd__inv_2 _23629_ (.A(_10181_),
    .Y(_00545_));
 sky130_fd_sc_hd__inv_2 _23630_ (.A(_10181_),
    .Y(_00546_));
 sky130_fd_sc_hd__inv_2 _23631_ (.A(_10181_),
    .Y(_00547_));
 sky130_fd_sc_hd__a21oi_4 _23632_ (.A1(_10142_),
    .A2(_09269_),
    .B1(_09361_),
    .Y(_10182_));
 sky130_fd_sc_hd__mux2_1 _23633_ (.A0(_09267_),
    .A1(\datamem.data_ram[59][8] ),
    .S(_10182_),
    .X(_10183_));
 sky130_fd_sc_hd__clkbuf_1 _23634_ (.A(_10183_),
    .X(_01740_));
 sky130_fd_sc_hd__mux2_1 _23635_ (.A0(_09273_),
    .A1(\datamem.data_ram[59][9] ),
    .S(_10182_),
    .X(_10184_));
 sky130_fd_sc_hd__clkbuf_1 _23636_ (.A(_10184_),
    .X(_01741_));
 sky130_fd_sc_hd__mux2_1 _23637_ (.A0(_09276_),
    .A1(\datamem.data_ram[59][10] ),
    .S(_10182_),
    .X(_10185_));
 sky130_fd_sc_hd__clkbuf_1 _23638_ (.A(_10185_),
    .X(_01742_));
 sky130_fd_sc_hd__mux2_1 _23639_ (.A0(_09279_),
    .A1(\datamem.data_ram[59][11] ),
    .S(_10182_),
    .X(_10186_));
 sky130_fd_sc_hd__clkbuf_1 _23640_ (.A(_10186_),
    .X(_01743_));
 sky130_fd_sc_hd__mux2_1 _23641_ (.A0(_09282_),
    .A1(\datamem.data_ram[59][12] ),
    .S(_10182_),
    .X(_10187_));
 sky130_fd_sc_hd__clkbuf_1 _23642_ (.A(_10187_),
    .X(_01744_));
 sky130_fd_sc_hd__mux2_1 _23643_ (.A0(_09285_),
    .A1(\datamem.data_ram[59][13] ),
    .S(_10182_),
    .X(_10188_));
 sky130_fd_sc_hd__clkbuf_1 _23644_ (.A(_10188_),
    .X(_01745_));
 sky130_fd_sc_hd__mux2_1 _23645_ (.A0(_09288_),
    .A1(\datamem.data_ram[59][14] ),
    .S(_10182_),
    .X(_10189_));
 sky130_fd_sc_hd__clkbuf_1 _23646_ (.A(_10189_),
    .X(_01746_));
 sky130_fd_sc_hd__mux2_1 _23647_ (.A0(_09291_),
    .A1(\datamem.data_ram[59][15] ),
    .S(_10182_),
    .X(_10190_));
 sky130_fd_sc_hd__clkbuf_1 _23648_ (.A(_10190_),
    .X(_01747_));
 sky130_fd_sc_hd__inv_2 _23649_ (.A(_10181_),
    .Y(_00548_));
 sky130_fd_sc_hd__inv_2 _23650_ (.A(_10181_),
    .Y(_00549_));
 sky130_fd_sc_hd__inv_2 _23651_ (.A(_10181_),
    .Y(_00550_));
 sky130_fd_sc_hd__inv_2 _23652_ (.A(_10181_),
    .Y(_00551_));
 sky130_fd_sc_hd__inv_2 _23653_ (.A(_10181_),
    .Y(_00552_));
 sky130_fd_sc_hd__inv_2 _23654_ (.A(_10181_),
    .Y(_00553_));
 sky130_fd_sc_hd__buf_1 _23655_ (.A(_10172_),
    .X(_10191_));
 sky130_fd_sc_hd__inv_2 _23656_ (.A(_10191_),
    .Y(_00554_));
 sky130_fd_sc_hd__inv_2 _23657_ (.A(_10191_),
    .Y(_00555_));
 sky130_fd_sc_hd__inv_2 _23658_ (.A(_10191_),
    .Y(_00556_));
 sky130_fd_sc_hd__inv_2 _23659_ (.A(_10191_),
    .Y(_00557_));
 sky130_fd_sc_hd__inv_2 _23660_ (.A(_10191_),
    .Y(_00558_));
 sky130_fd_sc_hd__inv_2 _23661_ (.A(_10191_),
    .Y(_00559_));
 sky130_fd_sc_hd__inv_2 _23662_ (.A(_10191_),
    .Y(_00560_));
 sky130_fd_sc_hd__inv_2 _23663_ (.A(_10191_),
    .Y(_00561_));
 sky130_fd_sc_hd__inv_2 _23664_ (.A(_10191_),
    .Y(_00562_));
 sky130_fd_sc_hd__inv_2 _23665_ (.A(_10191_),
    .Y(_00563_));
 sky130_fd_sc_hd__buf_1 _23666_ (.A(_10078_),
    .X(_10192_));
 sky130_fd_sc_hd__buf_1 _23667_ (.A(_10192_),
    .X(_10193_));
 sky130_fd_sc_hd__inv_2 _23668_ (.A(_10193_),
    .Y(_00564_));
 sky130_fd_sc_hd__inv_2 _23669_ (.A(_10193_),
    .Y(_00565_));
 sky130_fd_sc_hd__inv_2 _23670_ (.A(_10193_),
    .Y(_00566_));
 sky130_fd_sc_hd__inv_2 _23671_ (.A(_10193_),
    .Y(_00567_));
 sky130_fd_sc_hd__inv_2 _23672_ (.A(_10193_),
    .Y(_00568_));
 sky130_fd_sc_hd__inv_2 _23673_ (.A(_10193_),
    .Y(_00569_));
 sky130_fd_sc_hd__inv_2 _23674_ (.A(_10193_),
    .Y(_00570_));
 sky130_fd_sc_hd__inv_2 _23675_ (.A(_10193_),
    .Y(_00571_));
 sky130_fd_sc_hd__inv_2 _23676_ (.A(_10193_),
    .Y(_00572_));
 sky130_fd_sc_hd__inv_2 _23677_ (.A(_10193_),
    .Y(_00573_));
 sky130_fd_sc_hd__buf_1 _23678_ (.A(_10192_),
    .X(_10194_));
 sky130_fd_sc_hd__inv_2 _23679_ (.A(_10194_),
    .Y(_00574_));
 sky130_fd_sc_hd__inv_2 _23680_ (.A(_10194_),
    .Y(_00575_));
 sky130_fd_sc_hd__inv_2 _23681_ (.A(_10194_),
    .Y(_00576_));
 sky130_fd_sc_hd__inv_2 _23682_ (.A(_10194_),
    .Y(_00577_));
 sky130_fd_sc_hd__inv_2 _23683_ (.A(_10194_),
    .Y(_00578_));
 sky130_fd_sc_hd__inv_2 _23684_ (.A(_10194_),
    .Y(_00579_));
 sky130_fd_sc_hd__inv_2 _23685_ (.A(_10194_),
    .Y(_00580_));
 sky130_fd_sc_hd__inv_2 _23686_ (.A(_10194_),
    .Y(_00581_));
 sky130_fd_sc_hd__inv_2 _23687_ (.A(_10194_),
    .Y(_00582_));
 sky130_fd_sc_hd__inv_2 _23688_ (.A(_10194_),
    .Y(_00583_));
 sky130_fd_sc_hd__buf_1 _23689_ (.A(_10192_),
    .X(_10195_));
 sky130_fd_sc_hd__inv_2 _23690_ (.A(_10195_),
    .Y(_00584_));
 sky130_fd_sc_hd__inv_2 _23691_ (.A(_10195_),
    .Y(_00585_));
 sky130_fd_sc_hd__inv_2 _23692_ (.A(_10195_),
    .Y(_00586_));
 sky130_fd_sc_hd__inv_2 _23693_ (.A(_10195_),
    .Y(_00587_));
 sky130_fd_sc_hd__inv_2 _23694_ (.A(_10195_),
    .Y(_00588_));
 sky130_fd_sc_hd__inv_2 _23695_ (.A(_10195_),
    .Y(_00589_));
 sky130_fd_sc_hd__inv_2 _23696_ (.A(_10195_),
    .Y(_00590_));
 sky130_fd_sc_hd__inv_2 _23697_ (.A(_10195_),
    .Y(_00591_));
 sky130_fd_sc_hd__inv_2 _23698_ (.A(_10195_),
    .Y(_00592_));
 sky130_fd_sc_hd__inv_2 _23699_ (.A(_10195_),
    .Y(_00593_));
 sky130_fd_sc_hd__buf_1 _23700_ (.A(_10192_),
    .X(_10196_));
 sky130_fd_sc_hd__inv_2 _23701_ (.A(_10196_),
    .Y(_00594_));
 sky130_fd_sc_hd__inv_2 _23702_ (.A(_10196_),
    .Y(_00595_));
 sky130_fd_sc_hd__inv_2 _23703_ (.A(_10196_),
    .Y(_00596_));
 sky130_fd_sc_hd__inv_2 _23704_ (.A(_10196_),
    .Y(_00597_));
 sky130_fd_sc_hd__inv_2 _23705_ (.A(_10196_),
    .Y(_00598_));
 sky130_fd_sc_hd__inv_2 _23706_ (.A(_10196_),
    .Y(_00599_));
 sky130_fd_sc_hd__inv_2 _23707_ (.A(_10196_),
    .Y(_00600_));
 sky130_fd_sc_hd__inv_2 _23708_ (.A(_10196_),
    .Y(_00601_));
 sky130_fd_sc_hd__inv_2 _23709_ (.A(_10196_),
    .Y(_00602_));
 sky130_fd_sc_hd__inv_2 _23710_ (.A(_10196_),
    .Y(_00603_));
 sky130_fd_sc_hd__buf_1 _23711_ (.A(_10192_),
    .X(_10197_));
 sky130_fd_sc_hd__inv_2 _23712_ (.A(_10197_),
    .Y(_00604_));
 sky130_fd_sc_hd__inv_2 _23713_ (.A(_10197_),
    .Y(_00605_));
 sky130_fd_sc_hd__inv_2 _23714_ (.A(_10197_),
    .Y(_00606_));
 sky130_fd_sc_hd__inv_2 _23715_ (.A(_10197_),
    .Y(_00607_));
 sky130_fd_sc_hd__inv_2 _23716_ (.A(_10197_),
    .Y(_00608_));
 sky130_fd_sc_hd__inv_2 _23717_ (.A(_10197_),
    .Y(_00609_));
 sky130_fd_sc_hd__inv_2 _23718_ (.A(_10197_),
    .Y(_00610_));
 sky130_fd_sc_hd__inv_2 _23719_ (.A(_10197_),
    .Y(_00611_));
 sky130_fd_sc_hd__inv_2 _23720_ (.A(_10197_),
    .Y(_00612_));
 sky130_fd_sc_hd__inv_2 _23721_ (.A(_10197_),
    .Y(_00613_));
 sky130_fd_sc_hd__buf_1 _23722_ (.A(_10192_),
    .X(_10198_));
 sky130_fd_sc_hd__inv_2 _23723_ (.A(_10198_),
    .Y(_00614_));
 sky130_fd_sc_hd__inv_2 _23724_ (.A(_10198_),
    .Y(_00615_));
 sky130_fd_sc_hd__inv_2 _23725_ (.A(_10198_),
    .Y(_00616_));
 sky130_fd_sc_hd__inv_2 _23726_ (.A(_10198_),
    .Y(_00617_));
 sky130_fd_sc_hd__inv_2 _23727_ (.A(_10198_),
    .Y(_00618_));
 sky130_fd_sc_hd__inv_2 _23728_ (.A(_10198_),
    .Y(_00619_));
 sky130_fd_sc_hd__inv_2 _23729_ (.A(_10198_),
    .Y(_00620_));
 sky130_fd_sc_hd__inv_2 _23730_ (.A(_10198_),
    .Y(_00621_));
 sky130_fd_sc_hd__inv_2 _23731_ (.A(_10198_),
    .Y(_00622_));
 sky130_fd_sc_hd__inv_2 _23732_ (.A(_10198_),
    .Y(_00623_));
 sky130_fd_sc_hd__buf_1 _23733_ (.A(_10192_),
    .X(_10199_));
 sky130_fd_sc_hd__inv_2 _23734_ (.A(_10199_),
    .Y(_00624_));
 sky130_fd_sc_hd__inv_2 _23735_ (.A(_10199_),
    .Y(_00625_));
 sky130_fd_sc_hd__inv_2 _23736_ (.A(_10199_),
    .Y(_00626_));
 sky130_fd_sc_hd__inv_2 _23737_ (.A(_10199_),
    .Y(_00627_));
 sky130_fd_sc_hd__inv_2 _23738_ (.A(_10199_),
    .Y(_00628_));
 sky130_fd_sc_hd__inv_2 _23739_ (.A(_10199_),
    .Y(_00629_));
 sky130_fd_sc_hd__inv_2 _23740_ (.A(_10199_),
    .Y(_00630_));
 sky130_fd_sc_hd__inv_2 _23741_ (.A(_10199_),
    .Y(_00631_));
 sky130_fd_sc_hd__inv_2 _23742_ (.A(_10199_),
    .Y(_00632_));
 sky130_fd_sc_hd__inv_2 _23743_ (.A(_10199_),
    .Y(_00633_));
 sky130_fd_sc_hd__buf_1 _23744_ (.A(_10192_),
    .X(_10200_));
 sky130_fd_sc_hd__inv_2 _23745_ (.A(_10200_),
    .Y(_00634_));
 sky130_fd_sc_hd__inv_2 _23746_ (.A(_10200_),
    .Y(_00635_));
 sky130_fd_sc_hd__inv_2 _23747_ (.A(_10200_),
    .Y(_00636_));
 sky130_fd_sc_hd__inv_2 _23748_ (.A(_10200_),
    .Y(_00637_));
 sky130_fd_sc_hd__inv_2 _23749_ (.A(_10200_),
    .Y(_00638_));
 sky130_fd_sc_hd__inv_2 _23750_ (.A(_10200_),
    .Y(_00639_));
 sky130_fd_sc_hd__inv_2 _23751_ (.A(_10200_),
    .Y(_00640_));
 sky130_fd_sc_hd__inv_2 _23752_ (.A(_10200_),
    .Y(_00641_));
 sky130_fd_sc_hd__inv_2 _23753_ (.A(_10200_),
    .Y(_00642_));
 sky130_fd_sc_hd__inv_2 _23754_ (.A(_10200_),
    .Y(_00643_));
 sky130_fd_sc_hd__buf_1 _23755_ (.A(_10192_),
    .X(_10201_));
 sky130_fd_sc_hd__inv_2 _23756_ (.A(_10201_),
    .Y(_00644_));
 sky130_fd_sc_hd__inv_2 _23757_ (.A(_10201_),
    .Y(_00645_));
 sky130_fd_sc_hd__inv_2 _23758_ (.A(_10201_),
    .Y(_00646_));
 sky130_fd_sc_hd__inv_2 _23759_ (.A(_10201_),
    .Y(_00647_));
 sky130_fd_sc_hd__inv_2 _23760_ (.A(_10201_),
    .Y(_00648_));
 sky130_fd_sc_hd__inv_2 _23761_ (.A(_10201_),
    .Y(_00649_));
 sky130_fd_sc_hd__inv_2 _23762_ (.A(_10201_),
    .Y(_00650_));
 sky130_fd_sc_hd__inv_2 _23763_ (.A(_10201_),
    .Y(_00651_));
 sky130_fd_sc_hd__inv_2 _23764_ (.A(_10201_),
    .Y(_00652_));
 sky130_fd_sc_hd__inv_2 _23765_ (.A(_10201_),
    .Y(_00653_));
 sky130_fd_sc_hd__buf_1 _23766_ (.A(_10192_),
    .X(_10202_));
 sky130_fd_sc_hd__inv_2 _23767_ (.A(_10202_),
    .Y(_00654_));
 sky130_fd_sc_hd__inv_2 _23768_ (.A(_10202_),
    .Y(_00655_));
 sky130_fd_sc_hd__inv_2 _23769_ (.A(_10202_),
    .Y(_00656_));
 sky130_fd_sc_hd__inv_2 _23770_ (.A(_10202_),
    .Y(_00657_));
 sky130_fd_sc_hd__inv_2 _23771_ (.A(_10202_),
    .Y(_00658_));
 sky130_fd_sc_hd__inv_2 _23772_ (.A(_10202_),
    .Y(_00659_));
 sky130_fd_sc_hd__inv_2 _23773_ (.A(_10202_),
    .Y(_00660_));
 sky130_fd_sc_hd__inv_2 _23774_ (.A(_10202_),
    .Y(_00661_));
 sky130_fd_sc_hd__inv_2 _23775_ (.A(_10202_),
    .Y(_00662_));
 sky130_fd_sc_hd__inv_2 _23776_ (.A(_10202_),
    .Y(_00663_));
 sky130_fd_sc_hd__buf_1 _23777_ (.A(_10078_),
    .X(_10203_));
 sky130_fd_sc_hd__buf_1 _23778_ (.A(_10203_),
    .X(_10204_));
 sky130_fd_sc_hd__inv_2 _23779_ (.A(_10204_),
    .Y(_00664_));
 sky130_fd_sc_hd__inv_2 _23780_ (.A(_10204_),
    .Y(_00665_));
 sky130_fd_sc_hd__inv_2 _23781_ (.A(_10204_),
    .Y(_00666_));
 sky130_fd_sc_hd__inv_2 _23782_ (.A(_10204_),
    .Y(_00667_));
 sky130_fd_sc_hd__inv_2 _23783_ (.A(_10204_),
    .Y(_00668_));
 sky130_fd_sc_hd__inv_2 _23784_ (.A(_10204_),
    .Y(_00669_));
 sky130_fd_sc_hd__inv_2 _23785_ (.A(_10204_),
    .Y(_00670_));
 sky130_fd_sc_hd__inv_2 _23786_ (.A(_10204_),
    .Y(_00671_));
 sky130_fd_sc_hd__inv_2 _23787_ (.A(_10204_),
    .Y(_00672_));
 sky130_fd_sc_hd__inv_2 _23788_ (.A(_10204_),
    .Y(_00673_));
 sky130_fd_sc_hd__buf_1 _23789_ (.A(_10203_),
    .X(_10205_));
 sky130_fd_sc_hd__inv_2 _23790_ (.A(_10205_),
    .Y(_00674_));
 sky130_fd_sc_hd__inv_2 _23791_ (.A(_10205_),
    .Y(_00675_));
 sky130_fd_sc_hd__inv_2 _23792_ (.A(_10205_),
    .Y(_00676_));
 sky130_fd_sc_hd__inv_2 _23793_ (.A(_10205_),
    .Y(_00677_));
 sky130_fd_sc_hd__inv_2 _23794_ (.A(_10205_),
    .Y(_00678_));
 sky130_fd_sc_hd__inv_2 _23795_ (.A(_10205_),
    .Y(_00679_));
 sky130_fd_sc_hd__inv_2 _23796_ (.A(_10205_),
    .Y(_00680_));
 sky130_fd_sc_hd__inv_2 _23797_ (.A(_10205_),
    .Y(_00681_));
 sky130_fd_sc_hd__inv_2 _23798_ (.A(_10205_),
    .Y(_00682_));
 sky130_fd_sc_hd__inv_2 _23799_ (.A(_10205_),
    .Y(_00683_));
 sky130_fd_sc_hd__buf_1 _23800_ (.A(_10203_),
    .X(_10206_));
 sky130_fd_sc_hd__inv_2 _23801_ (.A(_10206_),
    .Y(_00684_));
 sky130_fd_sc_hd__inv_2 _23802_ (.A(_10206_),
    .Y(_00685_));
 sky130_fd_sc_hd__inv_2 _23803_ (.A(_10206_),
    .Y(_00686_));
 sky130_fd_sc_hd__inv_2 _23804_ (.A(_10206_),
    .Y(_00687_));
 sky130_fd_sc_hd__inv_2 _23805_ (.A(_10206_),
    .Y(_00688_));
 sky130_fd_sc_hd__inv_2 _23806_ (.A(_10206_),
    .Y(_00689_));
 sky130_fd_sc_hd__inv_2 _23807_ (.A(_10206_),
    .Y(_00690_));
 sky130_fd_sc_hd__inv_2 _23808_ (.A(_10206_),
    .Y(_00691_));
 sky130_fd_sc_hd__inv_2 _23809_ (.A(_10206_),
    .Y(_00692_));
 sky130_fd_sc_hd__inv_2 _23810_ (.A(_10206_),
    .Y(_00693_));
 sky130_fd_sc_hd__buf_1 _23811_ (.A(_10203_),
    .X(_10207_));
 sky130_fd_sc_hd__inv_2 _23812_ (.A(_10207_),
    .Y(_00694_));
 sky130_fd_sc_hd__inv_2 _23813_ (.A(_10207_),
    .Y(_00695_));
 sky130_fd_sc_hd__inv_2 _23814_ (.A(_10207_),
    .Y(_00696_));
 sky130_fd_sc_hd__inv_2 _23815_ (.A(_10207_),
    .Y(_00697_));
 sky130_fd_sc_hd__inv_2 _23816_ (.A(_10207_),
    .Y(_00698_));
 sky130_fd_sc_hd__inv_2 _23817_ (.A(_10207_),
    .Y(_00699_));
 sky130_fd_sc_hd__inv_2 _23818_ (.A(_10207_),
    .Y(_00700_));
 sky130_fd_sc_hd__inv_2 _23819_ (.A(_10207_),
    .Y(_00701_));
 sky130_fd_sc_hd__inv_2 _23820_ (.A(_10207_),
    .Y(_00702_));
 sky130_fd_sc_hd__inv_2 _23821_ (.A(_10207_),
    .Y(_00703_));
 sky130_fd_sc_hd__buf_1 _23822_ (.A(_10203_),
    .X(_10208_));
 sky130_fd_sc_hd__inv_2 _23823_ (.A(_10208_),
    .Y(_00704_));
 sky130_fd_sc_hd__inv_2 _23824_ (.A(_10208_),
    .Y(_00705_));
 sky130_fd_sc_hd__inv_2 _23825_ (.A(_10208_),
    .Y(_00706_));
 sky130_fd_sc_hd__inv_2 _23826_ (.A(_10208_),
    .Y(_00707_));
 sky130_fd_sc_hd__buf_8 _23827_ (.A(_07136_),
    .X(_10209_));
 sky130_fd_sc_hd__a21oi_4 _23828_ (.A1(_10209_),
    .A2(_09301_),
    .B1(_09361_),
    .Y(_10210_));
 sky130_fd_sc_hd__mux2_1 _23829_ (.A0(_09298_),
    .A1(\datamem.data_ram[58][24] ),
    .S(_10210_),
    .X(_10211_));
 sky130_fd_sc_hd__clkbuf_1 _23830_ (.A(_10211_),
    .X(_01908_));
 sky130_fd_sc_hd__mux2_1 _23831_ (.A0(_09306_),
    .A1(\datamem.data_ram[58][25] ),
    .S(_10210_),
    .X(_10212_));
 sky130_fd_sc_hd__clkbuf_1 _23832_ (.A(_10212_),
    .X(_01909_));
 sky130_fd_sc_hd__mux2_1 _23833_ (.A0(_09310_),
    .A1(\datamem.data_ram[58][26] ),
    .S(_10210_),
    .X(_10213_));
 sky130_fd_sc_hd__clkbuf_1 _23834_ (.A(_10213_),
    .X(_01910_));
 sky130_fd_sc_hd__mux2_1 _23835_ (.A0(_09314_),
    .A1(\datamem.data_ram[58][27] ),
    .S(_10210_),
    .X(_10214_));
 sky130_fd_sc_hd__clkbuf_1 _23836_ (.A(_10214_),
    .X(_01911_));
 sky130_fd_sc_hd__mux2_1 _23837_ (.A0(_09318_),
    .A1(\datamem.data_ram[58][28] ),
    .S(_10210_),
    .X(_10215_));
 sky130_fd_sc_hd__clkbuf_1 _23838_ (.A(_10215_),
    .X(_01912_));
 sky130_fd_sc_hd__mux2_1 _23839_ (.A0(_09322_),
    .A1(\datamem.data_ram[58][29] ),
    .S(_10210_),
    .X(_10216_));
 sky130_fd_sc_hd__clkbuf_1 _23840_ (.A(_10216_),
    .X(_01913_));
 sky130_fd_sc_hd__mux2_1 _23841_ (.A0(_09326_),
    .A1(\datamem.data_ram[58][30] ),
    .S(_10210_),
    .X(_10217_));
 sky130_fd_sc_hd__clkbuf_1 _23842_ (.A(_10217_),
    .X(_01914_));
 sky130_fd_sc_hd__mux2_1 _23843_ (.A0(_09330_),
    .A1(\datamem.data_ram[58][31] ),
    .S(_10210_),
    .X(_10218_));
 sky130_fd_sc_hd__clkbuf_1 _23844_ (.A(_10218_),
    .X(_01915_));
 sky130_fd_sc_hd__inv_2 _23845_ (.A(_10208_),
    .Y(_00708_));
 sky130_fd_sc_hd__inv_2 _23846_ (.A(_10208_),
    .Y(_00709_));
 sky130_fd_sc_hd__inv_2 _23847_ (.A(_10208_),
    .Y(_00710_));
 sky130_fd_sc_hd__inv_2 _23848_ (.A(_10208_),
    .Y(_00711_));
 sky130_fd_sc_hd__inv_2 _23849_ (.A(_10208_),
    .Y(_00712_));
 sky130_fd_sc_hd__inv_2 _23850_ (.A(_10208_),
    .Y(_00713_));
 sky130_fd_sc_hd__buf_1 _23851_ (.A(_10203_),
    .X(_10219_));
 sky130_fd_sc_hd__inv_2 _23852_ (.A(_10219_),
    .Y(_00714_));
 sky130_fd_sc_hd__inv_2 _23853_ (.A(_10219_),
    .Y(_00715_));
 sky130_fd_sc_hd__inv_2 _23854_ (.A(_10219_),
    .Y(_00716_));
 sky130_fd_sc_hd__inv_2 _23855_ (.A(_10219_),
    .Y(_00717_));
 sky130_fd_sc_hd__inv_2 _23856_ (.A(_10219_),
    .Y(_00718_));
 sky130_fd_sc_hd__inv_2 _23857_ (.A(_10219_),
    .Y(_00719_));
 sky130_fd_sc_hd__inv_2 _23858_ (.A(_10219_),
    .Y(_00720_));
 sky130_fd_sc_hd__inv_2 _23859_ (.A(_10219_),
    .Y(_00721_));
 sky130_fd_sc_hd__inv_2 _23860_ (.A(_10219_),
    .Y(_00722_));
 sky130_fd_sc_hd__inv_2 _23861_ (.A(_10219_),
    .Y(_00723_));
 sky130_fd_sc_hd__buf_1 _23862_ (.A(_10203_),
    .X(_10220_));
 sky130_fd_sc_hd__inv_2 _23863_ (.A(_10220_),
    .Y(_00724_));
 sky130_fd_sc_hd__inv_2 _23864_ (.A(_10220_),
    .Y(_00725_));
 sky130_fd_sc_hd__inv_2 _23865_ (.A(_10220_),
    .Y(_00726_));
 sky130_fd_sc_hd__inv_2 _23866_ (.A(_10220_),
    .Y(_00727_));
 sky130_fd_sc_hd__inv_2 _23867_ (.A(_10220_),
    .Y(_00728_));
 sky130_fd_sc_hd__inv_2 _23868_ (.A(_10220_),
    .Y(_00729_));
 sky130_fd_sc_hd__inv_2 _23869_ (.A(_10220_),
    .Y(_00730_));
 sky130_fd_sc_hd__inv_2 _23870_ (.A(_10220_),
    .Y(_00731_));
 sky130_fd_sc_hd__inv_2 _23871_ (.A(_10220_),
    .Y(_00732_));
 sky130_fd_sc_hd__inv_2 _23872_ (.A(_10220_),
    .Y(_00733_));
 sky130_fd_sc_hd__buf_1 _23873_ (.A(_10203_),
    .X(_10221_));
 sky130_fd_sc_hd__inv_2 _23874_ (.A(_10221_),
    .Y(_00734_));
 sky130_fd_sc_hd__inv_2 _23875_ (.A(_10221_),
    .Y(_00735_));
 sky130_fd_sc_hd__inv_2 _23876_ (.A(_10221_),
    .Y(_00736_));
 sky130_fd_sc_hd__inv_2 _23877_ (.A(_10221_),
    .Y(_00737_));
 sky130_fd_sc_hd__inv_2 _23878_ (.A(_10221_),
    .Y(_00738_));
 sky130_fd_sc_hd__inv_2 _23879_ (.A(_10221_),
    .Y(_00739_));
 sky130_fd_sc_hd__inv_2 _23880_ (.A(_10221_),
    .Y(_00740_));
 sky130_fd_sc_hd__inv_2 _23881_ (.A(_10221_),
    .Y(_00741_));
 sky130_fd_sc_hd__inv_2 _23882_ (.A(_10221_),
    .Y(_00742_));
 sky130_fd_sc_hd__inv_2 _23883_ (.A(_10221_),
    .Y(_00743_));
 sky130_fd_sc_hd__buf_1 _23884_ (.A(_10203_),
    .X(_10222_));
 sky130_fd_sc_hd__inv_2 _23885_ (.A(_10222_),
    .Y(_00744_));
 sky130_fd_sc_hd__inv_2 _23886_ (.A(_10222_),
    .Y(_00745_));
 sky130_fd_sc_hd__inv_2 _23887_ (.A(_10222_),
    .Y(_00746_));
 sky130_fd_sc_hd__inv_2 _23888_ (.A(_10222_),
    .Y(_00747_));
 sky130_fd_sc_hd__inv_2 _23889_ (.A(_10222_),
    .Y(_00748_));
 sky130_fd_sc_hd__inv_2 _23890_ (.A(_10222_),
    .Y(_00749_));
 sky130_fd_sc_hd__inv_2 _23891_ (.A(_10222_),
    .Y(_00750_));
 sky130_fd_sc_hd__inv_2 _23892_ (.A(_10222_),
    .Y(_00751_));
 sky130_fd_sc_hd__inv_2 _23893_ (.A(_10222_),
    .Y(_00752_));
 sky130_fd_sc_hd__inv_2 _23894_ (.A(_10222_),
    .Y(_00753_));
 sky130_fd_sc_hd__buf_1 _23895_ (.A(_10203_),
    .X(_10223_));
 sky130_fd_sc_hd__inv_2 _23896_ (.A(_10223_),
    .Y(_00754_));
 sky130_fd_sc_hd__inv_2 _23897_ (.A(_10223_),
    .Y(_00755_));
 sky130_fd_sc_hd__inv_2 _23898_ (.A(_10223_),
    .Y(_00756_));
 sky130_fd_sc_hd__inv_2 _23899_ (.A(_10223_),
    .Y(_00757_));
 sky130_fd_sc_hd__inv_2 _23900_ (.A(_10223_),
    .Y(_00758_));
 sky130_fd_sc_hd__inv_2 _23901_ (.A(_10223_),
    .Y(_00759_));
 sky130_fd_sc_hd__inv_2 _23902_ (.A(_10223_),
    .Y(_00760_));
 sky130_fd_sc_hd__inv_2 _23903_ (.A(_10223_),
    .Y(_00761_));
 sky130_fd_sc_hd__inv_2 _23904_ (.A(_10223_),
    .Y(_00762_));
 sky130_fd_sc_hd__inv_2 _23905_ (.A(_10223_),
    .Y(_00763_));
 sky130_fd_sc_hd__buf_1 _23906_ (.A(_10078_),
    .X(_10224_));
 sky130_fd_sc_hd__buf_1 _23907_ (.A(_10224_),
    .X(_10225_));
 sky130_fd_sc_hd__inv_2 _23908_ (.A(_10225_),
    .Y(_00764_));
 sky130_fd_sc_hd__inv_2 _23909_ (.A(_10225_),
    .Y(_00765_));
 sky130_fd_sc_hd__inv_2 _23910_ (.A(_10225_),
    .Y(_00766_));
 sky130_fd_sc_hd__inv_2 _23911_ (.A(_10225_),
    .Y(_00767_));
 sky130_fd_sc_hd__inv_2 _23912_ (.A(_10225_),
    .Y(_00768_));
 sky130_fd_sc_hd__inv_2 _23913_ (.A(_10225_),
    .Y(_00769_));
 sky130_fd_sc_hd__inv_2 _23914_ (.A(_10225_),
    .Y(_00770_));
 sky130_fd_sc_hd__inv_2 _23915_ (.A(_10225_),
    .Y(_00771_));
 sky130_fd_sc_hd__inv_2 _23916_ (.A(_10225_),
    .Y(_00772_));
 sky130_fd_sc_hd__inv_2 _23917_ (.A(_10225_),
    .Y(_00773_));
 sky130_fd_sc_hd__buf_1 _23918_ (.A(_10224_),
    .X(_10226_));
 sky130_fd_sc_hd__inv_2 _23919_ (.A(_10226_),
    .Y(_00774_));
 sky130_fd_sc_hd__inv_2 _23920_ (.A(_10226_),
    .Y(_00775_));
 sky130_fd_sc_hd__inv_2 _23921_ (.A(_10226_),
    .Y(_00776_));
 sky130_fd_sc_hd__inv_2 _23922_ (.A(_10226_),
    .Y(_00777_));
 sky130_fd_sc_hd__inv_2 _23923_ (.A(_10226_),
    .Y(_00778_));
 sky130_fd_sc_hd__inv_2 _23924_ (.A(_10226_),
    .Y(_00779_));
 sky130_fd_sc_hd__inv_2 _23925_ (.A(_10226_),
    .Y(_00780_));
 sky130_fd_sc_hd__inv_2 _23926_ (.A(_10226_),
    .Y(_00781_));
 sky130_fd_sc_hd__inv_2 _23927_ (.A(_10226_),
    .Y(_00782_));
 sky130_fd_sc_hd__inv_2 _23928_ (.A(_10226_),
    .Y(_00783_));
 sky130_fd_sc_hd__buf_1 _23929_ (.A(_10224_),
    .X(_10227_));
 sky130_fd_sc_hd__inv_2 _23930_ (.A(_10227_),
    .Y(_00784_));
 sky130_fd_sc_hd__inv_2 _23931_ (.A(_10227_),
    .Y(_00785_));
 sky130_fd_sc_hd__inv_2 _23932_ (.A(_10227_),
    .Y(_00786_));
 sky130_fd_sc_hd__inv_2 _23933_ (.A(_10227_),
    .Y(_00787_));
 sky130_fd_sc_hd__inv_2 _23934_ (.A(_10227_),
    .Y(_00788_));
 sky130_fd_sc_hd__inv_2 _23935_ (.A(_10227_),
    .Y(_00789_));
 sky130_fd_sc_hd__inv_2 _23936_ (.A(_10227_),
    .Y(_00790_));
 sky130_fd_sc_hd__inv_2 _23937_ (.A(_10227_),
    .Y(_00791_));
 sky130_fd_sc_hd__inv_2 _23938_ (.A(_10227_),
    .Y(_00792_));
 sky130_fd_sc_hd__inv_2 _23939_ (.A(_10227_),
    .Y(_00793_));
 sky130_fd_sc_hd__buf_1 _23940_ (.A(_10224_),
    .X(_10228_));
 sky130_fd_sc_hd__inv_2 _23941_ (.A(_10228_),
    .Y(_00794_));
 sky130_fd_sc_hd__inv_2 _23942_ (.A(_10228_),
    .Y(_00795_));
 sky130_fd_sc_hd__inv_2 _23943_ (.A(_10228_),
    .Y(_00796_));
 sky130_fd_sc_hd__inv_2 _23944_ (.A(_10228_),
    .Y(_00797_));
 sky130_fd_sc_hd__inv_2 _23945_ (.A(_10228_),
    .Y(_00798_));
 sky130_fd_sc_hd__inv_2 _23946_ (.A(_10228_),
    .Y(_00799_));
 sky130_fd_sc_hd__inv_2 _23947_ (.A(_10228_),
    .Y(_00800_));
 sky130_fd_sc_hd__inv_2 _23948_ (.A(_10228_),
    .Y(_00801_));
 sky130_fd_sc_hd__inv_2 _23949_ (.A(_10228_),
    .Y(_00802_));
 sky130_fd_sc_hd__inv_2 _23950_ (.A(_10228_),
    .Y(_00803_));
 sky130_fd_sc_hd__a21oi_4 _23951_ (.A1(_10209_),
    .A2(_09229_),
    .B1(_09361_),
    .Y(_10229_));
 sky130_fd_sc_hd__mux2_1 _23952_ (.A0(_09224_),
    .A1(\datamem.data_ram[58][16] ),
    .S(_10229_),
    .X(_10230_));
 sky130_fd_sc_hd__clkbuf_1 _23953_ (.A(_10230_),
    .X(_02012_));
 sky130_fd_sc_hd__mux2_1 _23954_ (.A0(_09236_),
    .A1(\datamem.data_ram[58][17] ),
    .S(_10229_),
    .X(_10231_));
 sky130_fd_sc_hd__clkbuf_1 _23955_ (.A(_10231_),
    .X(_02013_));
 sky130_fd_sc_hd__mux2_1 _23956_ (.A0(_09240_),
    .A1(\datamem.data_ram[58][18] ),
    .S(_10229_),
    .X(_10232_));
 sky130_fd_sc_hd__clkbuf_1 _23957_ (.A(_10232_),
    .X(_02014_));
 sky130_fd_sc_hd__mux2_1 _23958_ (.A0(_09244_),
    .A1(\datamem.data_ram[58][19] ),
    .S(_10229_),
    .X(_10233_));
 sky130_fd_sc_hd__clkbuf_1 _23959_ (.A(_10233_),
    .X(_02015_));
 sky130_fd_sc_hd__mux2_1 _23960_ (.A0(_09248_),
    .A1(\datamem.data_ram[58][20] ),
    .S(_10229_),
    .X(_10234_));
 sky130_fd_sc_hd__clkbuf_1 _23961_ (.A(_10234_),
    .X(_02016_));
 sky130_fd_sc_hd__mux2_1 _23962_ (.A0(_09252_),
    .A1(\datamem.data_ram[58][21] ),
    .S(_10229_),
    .X(_10235_));
 sky130_fd_sc_hd__clkbuf_1 _23963_ (.A(_10235_),
    .X(_02017_));
 sky130_fd_sc_hd__mux2_1 _23964_ (.A0(_09256_),
    .A1(\datamem.data_ram[58][22] ),
    .S(_10229_),
    .X(_10236_));
 sky130_fd_sc_hd__clkbuf_1 _23965_ (.A(_10236_),
    .X(_02018_));
 sky130_fd_sc_hd__mux2_1 _23966_ (.A0(_09260_),
    .A1(\datamem.data_ram[58][23] ),
    .S(_10229_),
    .X(_10237_));
 sky130_fd_sc_hd__clkbuf_1 _23967_ (.A(_10237_),
    .X(_02019_));
 sky130_fd_sc_hd__buf_1 _23968_ (.A(_10224_),
    .X(_10238_));
 sky130_fd_sc_hd__inv_2 _23969_ (.A(_10238_),
    .Y(_00804_));
 sky130_fd_sc_hd__inv_2 _23970_ (.A(_10238_),
    .Y(_00805_));
 sky130_fd_sc_hd__inv_2 _23971_ (.A(_10238_),
    .Y(_00806_));
 sky130_fd_sc_hd__inv_2 _23972_ (.A(_10238_),
    .Y(_00807_));
 sky130_fd_sc_hd__inv_2 _23973_ (.A(_10238_),
    .Y(_00808_));
 sky130_fd_sc_hd__inv_2 _23974_ (.A(_10238_),
    .Y(_00809_));
 sky130_fd_sc_hd__inv_2 _23975_ (.A(_10238_),
    .Y(_00810_));
 sky130_fd_sc_hd__inv_2 _23976_ (.A(_10238_),
    .Y(_00811_));
 sky130_fd_sc_hd__inv_2 _23977_ (.A(_10238_),
    .Y(_00812_));
 sky130_fd_sc_hd__inv_2 _23978_ (.A(_10238_),
    .Y(_00813_));
 sky130_fd_sc_hd__buf_1 _23979_ (.A(_10224_),
    .X(_10239_));
 sky130_fd_sc_hd__inv_2 _23980_ (.A(_10239_),
    .Y(_00814_));
 sky130_fd_sc_hd__inv_2 _23981_ (.A(_10239_),
    .Y(_00815_));
 sky130_fd_sc_hd__inv_2 _23982_ (.A(_10239_),
    .Y(_00816_));
 sky130_fd_sc_hd__inv_2 _23983_ (.A(_10239_),
    .Y(_00817_));
 sky130_fd_sc_hd__inv_2 _23984_ (.A(_10239_),
    .Y(_00818_));
 sky130_fd_sc_hd__inv_2 _23985_ (.A(_10239_),
    .Y(_00819_));
 sky130_fd_sc_hd__inv_2 _23986_ (.A(_10239_),
    .Y(_00820_));
 sky130_fd_sc_hd__inv_2 _23987_ (.A(_10239_),
    .Y(_00821_));
 sky130_fd_sc_hd__inv_2 _23988_ (.A(_10239_),
    .Y(_00822_));
 sky130_fd_sc_hd__inv_2 _23989_ (.A(_10239_),
    .Y(_00823_));
 sky130_fd_sc_hd__buf_1 _23990_ (.A(_10224_),
    .X(_10240_));
 sky130_fd_sc_hd__inv_2 _23991_ (.A(_10240_),
    .Y(_00824_));
 sky130_fd_sc_hd__inv_2 _23992_ (.A(_10240_),
    .Y(_00825_));
 sky130_fd_sc_hd__inv_2 _23993_ (.A(_10240_),
    .Y(_00826_));
 sky130_fd_sc_hd__inv_2 _23994_ (.A(_10240_),
    .Y(_00827_));
 sky130_fd_sc_hd__inv_2 _23995_ (.A(_10240_),
    .Y(_00828_));
 sky130_fd_sc_hd__inv_2 _23996_ (.A(_10240_),
    .Y(_00829_));
 sky130_fd_sc_hd__inv_2 _23997_ (.A(_10240_),
    .Y(_00830_));
 sky130_fd_sc_hd__inv_2 _23998_ (.A(_10240_),
    .Y(_00831_));
 sky130_fd_sc_hd__inv_2 _23999_ (.A(_10240_),
    .Y(_00832_));
 sky130_fd_sc_hd__inv_2 _24000_ (.A(_10240_),
    .Y(_00833_));
 sky130_fd_sc_hd__buf_1 _24001_ (.A(_10224_),
    .X(_10241_));
 sky130_fd_sc_hd__inv_2 _24002_ (.A(_10241_),
    .Y(_00834_));
 sky130_fd_sc_hd__inv_2 _24003_ (.A(_10241_),
    .Y(_00835_));
 sky130_fd_sc_hd__inv_2 _24004_ (.A(_10241_),
    .Y(_00836_));
 sky130_fd_sc_hd__inv_2 _24005_ (.A(_10241_),
    .Y(_00837_));
 sky130_fd_sc_hd__inv_2 _24006_ (.A(_10241_),
    .Y(_00838_));
 sky130_fd_sc_hd__inv_2 _24007_ (.A(_10241_),
    .Y(_00839_));
 sky130_fd_sc_hd__inv_2 _24008_ (.A(_10241_),
    .Y(_00840_));
 sky130_fd_sc_hd__inv_2 _24009_ (.A(_10241_),
    .Y(_00841_));
 sky130_fd_sc_hd__inv_2 _24010_ (.A(_10241_),
    .Y(_00842_));
 sky130_fd_sc_hd__inv_2 _24011_ (.A(_10241_),
    .Y(_00843_));
 sky130_fd_sc_hd__buf_1 _24012_ (.A(_10224_),
    .X(_10242_));
 sky130_fd_sc_hd__inv_2 _24013_ (.A(_10242_),
    .Y(_00844_));
 sky130_fd_sc_hd__inv_2 _24014_ (.A(_10242_),
    .Y(_00845_));
 sky130_fd_sc_hd__inv_2 _24015_ (.A(_10242_),
    .Y(_00846_));
 sky130_fd_sc_hd__inv_2 _24016_ (.A(_10242_),
    .Y(_00847_));
 sky130_fd_sc_hd__inv_2 _24017_ (.A(_10242_),
    .Y(_00848_));
 sky130_fd_sc_hd__inv_2 _24018_ (.A(_10242_),
    .Y(_00849_));
 sky130_fd_sc_hd__inv_2 _24019_ (.A(_10242_),
    .Y(_00850_));
 sky130_fd_sc_hd__inv_2 _24020_ (.A(_10242_),
    .Y(_00851_));
 sky130_fd_sc_hd__inv_2 _24021_ (.A(_10242_),
    .Y(_00852_));
 sky130_fd_sc_hd__inv_2 _24022_ (.A(_10242_),
    .Y(_00853_));
 sky130_fd_sc_hd__buf_1 _24023_ (.A(_10224_),
    .X(_10243_));
 sky130_fd_sc_hd__inv_2 _24024_ (.A(_10243_),
    .Y(_00854_));
 sky130_fd_sc_hd__inv_2 _24025_ (.A(_10243_),
    .Y(_00855_));
 sky130_fd_sc_hd__inv_2 _24026_ (.A(_10243_),
    .Y(_00856_));
 sky130_fd_sc_hd__inv_2 _24027_ (.A(_10243_),
    .Y(_00857_));
 sky130_fd_sc_hd__inv_2 _24028_ (.A(_10243_),
    .Y(_00858_));
 sky130_fd_sc_hd__inv_2 _24029_ (.A(_10243_),
    .Y(_00859_));
 sky130_fd_sc_hd__inv_2 _24030_ (.A(_10243_),
    .Y(_00860_));
 sky130_fd_sc_hd__inv_2 _24031_ (.A(_10243_),
    .Y(_00861_));
 sky130_fd_sc_hd__inv_2 _24032_ (.A(_10243_),
    .Y(_00862_));
 sky130_fd_sc_hd__inv_2 _24033_ (.A(_10243_),
    .Y(_00863_));
 sky130_fd_sc_hd__buf_1 _24034_ (.A(_10078_),
    .X(_10244_));
 sky130_fd_sc_hd__buf_1 _24035_ (.A(_10244_),
    .X(_10245_));
 sky130_fd_sc_hd__inv_2 _24036_ (.A(_10245_),
    .Y(_00864_));
 sky130_fd_sc_hd__inv_2 _24037_ (.A(_10245_),
    .Y(_00865_));
 sky130_fd_sc_hd__inv_2 _24038_ (.A(_10245_),
    .Y(_00866_));
 sky130_fd_sc_hd__inv_2 _24039_ (.A(_10245_),
    .Y(_00867_));
 sky130_fd_sc_hd__inv_2 _24040_ (.A(_10245_),
    .Y(_00868_));
 sky130_fd_sc_hd__inv_2 _24041_ (.A(_10245_),
    .Y(_00869_));
 sky130_fd_sc_hd__inv_2 _24042_ (.A(_10245_),
    .Y(_00870_));
 sky130_fd_sc_hd__inv_2 _24043_ (.A(_10245_),
    .Y(_00871_));
 sky130_fd_sc_hd__inv_2 _24044_ (.A(_10245_),
    .Y(_00872_));
 sky130_fd_sc_hd__inv_2 _24045_ (.A(_10245_),
    .Y(_00873_));
 sky130_fd_sc_hd__buf_1 _24046_ (.A(_10244_),
    .X(_10246_));
 sky130_fd_sc_hd__inv_2 _24047_ (.A(_10246_),
    .Y(_00874_));
 sky130_fd_sc_hd__inv_2 _24048_ (.A(_10246_),
    .Y(_00875_));
 sky130_fd_sc_hd__inv_2 _24049_ (.A(_10246_),
    .Y(_00876_));
 sky130_fd_sc_hd__inv_2 _24050_ (.A(_10246_),
    .Y(_00877_));
 sky130_fd_sc_hd__inv_2 _24051_ (.A(_10246_),
    .Y(_00878_));
 sky130_fd_sc_hd__inv_2 _24052_ (.A(_10246_),
    .Y(_00879_));
 sky130_fd_sc_hd__inv_2 _24053_ (.A(_10246_),
    .Y(_00880_));
 sky130_fd_sc_hd__inv_2 _24054_ (.A(_10246_),
    .Y(_00881_));
 sky130_fd_sc_hd__inv_2 _24055_ (.A(_10246_),
    .Y(_00882_));
 sky130_fd_sc_hd__inv_2 _24056_ (.A(_10246_),
    .Y(_00883_));
 sky130_fd_sc_hd__buf_1 _24057_ (.A(_10244_),
    .X(_10247_));
 sky130_fd_sc_hd__inv_2 _24058_ (.A(_10247_),
    .Y(_00884_));
 sky130_fd_sc_hd__inv_2 _24059_ (.A(_10247_),
    .Y(_00885_));
 sky130_fd_sc_hd__inv_2 _24060_ (.A(_10247_),
    .Y(_00886_));
 sky130_fd_sc_hd__inv_2 _24061_ (.A(_10247_),
    .Y(_00887_));
 sky130_fd_sc_hd__inv_2 _24062_ (.A(_10247_),
    .Y(_00888_));
 sky130_fd_sc_hd__inv_2 _24063_ (.A(_10247_),
    .Y(_00889_));
 sky130_fd_sc_hd__inv_2 _24064_ (.A(_10247_),
    .Y(_00890_));
 sky130_fd_sc_hd__inv_2 _24065_ (.A(_10247_),
    .Y(_00891_));
 sky130_fd_sc_hd__inv_2 _24066_ (.A(_10247_),
    .Y(_00892_));
 sky130_fd_sc_hd__inv_2 _24067_ (.A(_10247_),
    .Y(_00893_));
 sky130_fd_sc_hd__buf_1 _24068_ (.A(_10244_),
    .X(_10248_));
 sky130_fd_sc_hd__inv_2 _24069_ (.A(_10248_),
    .Y(_00894_));
 sky130_fd_sc_hd__inv_2 _24070_ (.A(_10248_),
    .Y(_00895_));
 sky130_fd_sc_hd__inv_2 _24071_ (.A(_10248_),
    .Y(_00896_));
 sky130_fd_sc_hd__inv_2 _24072_ (.A(_10248_),
    .Y(_00897_));
 sky130_fd_sc_hd__inv_2 _24073_ (.A(_10248_),
    .Y(_00898_));
 sky130_fd_sc_hd__inv_2 _24074_ (.A(_10248_),
    .Y(_00899_));
 sky130_fd_sc_hd__a21oi_4 _24075_ (.A1(_10209_),
    .A2(_09269_),
    .B1(_09361_),
    .Y(_10249_));
 sky130_fd_sc_hd__mux2_1 _24076_ (.A0(_09267_),
    .A1(\datamem.data_ram[58][8] ),
    .S(_10249_),
    .X(_10250_));
 sky130_fd_sc_hd__clkbuf_1 _24077_ (.A(_10250_),
    .X(_02116_));
 sky130_fd_sc_hd__mux2_1 _24078_ (.A0(_09273_),
    .A1(\datamem.data_ram[58][9] ),
    .S(_10249_),
    .X(_10251_));
 sky130_fd_sc_hd__clkbuf_1 _24079_ (.A(_10251_),
    .X(_02117_));
 sky130_fd_sc_hd__mux2_1 _24080_ (.A0(_09276_),
    .A1(\datamem.data_ram[58][10] ),
    .S(_10249_),
    .X(_10252_));
 sky130_fd_sc_hd__clkbuf_1 _24081_ (.A(_10252_),
    .X(_02118_));
 sky130_fd_sc_hd__mux2_1 _24082_ (.A0(_09279_),
    .A1(\datamem.data_ram[58][11] ),
    .S(_10249_),
    .X(_10253_));
 sky130_fd_sc_hd__clkbuf_1 _24083_ (.A(_10253_),
    .X(_02119_));
 sky130_fd_sc_hd__mux2_1 _24084_ (.A0(_09282_),
    .A1(\datamem.data_ram[58][12] ),
    .S(_10249_),
    .X(_10254_));
 sky130_fd_sc_hd__clkbuf_1 _24085_ (.A(_10254_),
    .X(_02120_));
 sky130_fd_sc_hd__mux2_1 _24086_ (.A0(_09285_),
    .A1(\datamem.data_ram[58][13] ),
    .S(_10249_),
    .X(_10255_));
 sky130_fd_sc_hd__clkbuf_1 _24087_ (.A(_10255_),
    .X(_02121_));
 sky130_fd_sc_hd__mux2_1 _24088_ (.A0(_09288_),
    .A1(\datamem.data_ram[58][14] ),
    .S(_10249_),
    .X(_10256_));
 sky130_fd_sc_hd__clkbuf_1 _24089_ (.A(_10256_),
    .X(_02122_));
 sky130_fd_sc_hd__mux2_1 _24090_ (.A0(_09291_),
    .A1(\datamem.data_ram[58][15] ),
    .S(_10249_),
    .X(_10257_));
 sky130_fd_sc_hd__clkbuf_1 _24091_ (.A(_10257_),
    .X(_02123_));
 sky130_fd_sc_hd__inv_2 _24092_ (.A(_10248_),
    .Y(_00900_));
 sky130_fd_sc_hd__inv_2 _24093_ (.A(_10248_),
    .Y(_00901_));
 sky130_fd_sc_hd__inv_2 _24094_ (.A(_10248_),
    .Y(_00902_));
 sky130_fd_sc_hd__inv_2 _24095_ (.A(_10248_),
    .Y(_00903_));
 sky130_fd_sc_hd__buf_1 _24096_ (.A(_10244_),
    .X(_10258_));
 sky130_fd_sc_hd__inv_2 _24097_ (.A(_10258_),
    .Y(_00904_));
 sky130_fd_sc_hd__inv_2 _24098_ (.A(_10258_),
    .Y(_00905_));
 sky130_fd_sc_hd__inv_2 _24099_ (.A(_10258_),
    .Y(_00906_));
 sky130_fd_sc_hd__inv_2 _24100_ (.A(_10258_),
    .Y(_00907_));
 sky130_fd_sc_hd__inv_2 _24101_ (.A(_10258_),
    .Y(_00908_));
 sky130_fd_sc_hd__inv_2 _24102_ (.A(_10258_),
    .Y(_00909_));
 sky130_fd_sc_hd__inv_2 _24103_ (.A(_10258_),
    .Y(_00910_));
 sky130_fd_sc_hd__inv_2 _24104_ (.A(_10258_),
    .Y(_00911_));
 sky130_fd_sc_hd__inv_2 _24105_ (.A(_10258_),
    .Y(_00912_));
 sky130_fd_sc_hd__inv_2 _24106_ (.A(_10258_),
    .Y(_00913_));
 sky130_fd_sc_hd__buf_1 _24107_ (.A(_10244_),
    .X(_10259_));
 sky130_fd_sc_hd__inv_2 _24108_ (.A(_10259_),
    .Y(_00914_));
 sky130_fd_sc_hd__inv_2 _24109_ (.A(_10259_),
    .Y(_00915_));
 sky130_fd_sc_hd__inv_2 _24110_ (.A(_10259_),
    .Y(_00916_));
 sky130_fd_sc_hd__inv_2 _24111_ (.A(_10259_),
    .Y(_00917_));
 sky130_fd_sc_hd__inv_2 _24112_ (.A(_10259_),
    .Y(_00918_));
 sky130_fd_sc_hd__inv_2 _24113_ (.A(_10259_),
    .Y(_00919_));
 sky130_fd_sc_hd__inv_2 _24114_ (.A(_10259_),
    .Y(_00920_));
 sky130_fd_sc_hd__inv_2 _24115_ (.A(_10259_),
    .Y(_00921_));
 sky130_fd_sc_hd__inv_2 _24116_ (.A(_10259_),
    .Y(_00922_));
 sky130_fd_sc_hd__inv_2 _24117_ (.A(_10259_),
    .Y(_00923_));
 sky130_fd_sc_hd__buf_1 _24118_ (.A(_10244_),
    .X(_10260_));
 sky130_fd_sc_hd__inv_2 _24119_ (.A(_10260_),
    .Y(_00924_));
 sky130_fd_sc_hd__inv_2 _24120_ (.A(_10260_),
    .Y(_00925_));
 sky130_fd_sc_hd__inv_2 _24121_ (.A(_10260_),
    .Y(_00926_));
 sky130_fd_sc_hd__inv_2 _24122_ (.A(_10260_),
    .Y(_00927_));
 sky130_fd_sc_hd__inv_2 _24123_ (.A(_10260_),
    .Y(_00928_));
 sky130_fd_sc_hd__inv_2 _24124_ (.A(_10260_),
    .Y(_00929_));
 sky130_fd_sc_hd__inv_2 _24125_ (.A(_10260_),
    .Y(_00930_));
 sky130_fd_sc_hd__inv_2 _24126_ (.A(_10260_),
    .Y(_00931_));
 sky130_fd_sc_hd__inv_2 _24127_ (.A(_10260_),
    .Y(_00932_));
 sky130_fd_sc_hd__inv_2 _24128_ (.A(_10260_),
    .Y(_00933_));
 sky130_fd_sc_hd__buf_1 _24129_ (.A(_10244_),
    .X(_10261_));
 sky130_fd_sc_hd__inv_2 _24130_ (.A(_10261_),
    .Y(_00934_));
 sky130_fd_sc_hd__inv_2 _24131_ (.A(_10261_),
    .Y(_00935_));
 sky130_fd_sc_hd__inv_2 _24132_ (.A(_10261_),
    .Y(_00936_));
 sky130_fd_sc_hd__inv_2 _24133_ (.A(_10261_),
    .Y(_00937_));
 sky130_fd_sc_hd__inv_2 _24134_ (.A(_10261_),
    .Y(_00938_));
 sky130_fd_sc_hd__inv_2 _24135_ (.A(_10261_),
    .Y(_00939_));
 sky130_fd_sc_hd__inv_2 _24136_ (.A(_10261_),
    .Y(_00940_));
 sky130_fd_sc_hd__inv_2 _24137_ (.A(_10261_),
    .Y(_00941_));
 sky130_fd_sc_hd__inv_2 _24138_ (.A(_10261_),
    .Y(_00942_));
 sky130_fd_sc_hd__inv_2 _24139_ (.A(_10261_),
    .Y(_00943_));
 sky130_fd_sc_hd__buf_1 _24140_ (.A(_10244_),
    .X(_10262_));
 sky130_fd_sc_hd__inv_2 _24141_ (.A(_10262_),
    .Y(_00944_));
 sky130_fd_sc_hd__inv_2 _24142_ (.A(_10262_),
    .Y(_00945_));
 sky130_fd_sc_hd__inv_2 _24143_ (.A(_10262_),
    .Y(_00946_));
 sky130_fd_sc_hd__inv_2 _24144_ (.A(_10262_),
    .Y(_00947_));
 sky130_fd_sc_hd__inv_2 _24145_ (.A(_10262_),
    .Y(_00948_));
 sky130_fd_sc_hd__inv_2 _24146_ (.A(_10262_),
    .Y(_00949_));
 sky130_fd_sc_hd__inv_2 _24147_ (.A(_10262_),
    .Y(_00950_));
 sky130_fd_sc_hd__inv_2 _24148_ (.A(_10262_),
    .Y(_00951_));
 sky130_fd_sc_hd__inv_2 _24149_ (.A(_10262_),
    .Y(_00952_));
 sky130_fd_sc_hd__inv_2 _24150_ (.A(_10262_),
    .Y(_00953_));
 sky130_fd_sc_hd__buf_1 _24151_ (.A(_10244_),
    .X(_10263_));
 sky130_fd_sc_hd__inv_2 _24152_ (.A(_10263_),
    .Y(_00954_));
 sky130_fd_sc_hd__inv_2 _24153_ (.A(_10263_),
    .Y(_00955_));
 sky130_fd_sc_hd__inv_2 _24154_ (.A(_10263_),
    .Y(_00956_));
 sky130_fd_sc_hd__inv_2 _24155_ (.A(_10263_),
    .Y(_00957_));
 sky130_fd_sc_hd__inv_2 _24156_ (.A(_10263_),
    .Y(_00958_));
 sky130_fd_sc_hd__inv_2 _24157_ (.A(_10263_),
    .Y(_00959_));
 sky130_fd_sc_hd__inv_2 _24158_ (.A(_10263_),
    .Y(_00960_));
 sky130_fd_sc_hd__inv_2 _24159_ (.A(_10263_),
    .Y(_00961_));
 sky130_fd_sc_hd__inv_2 _24160_ (.A(_10263_),
    .Y(_00962_));
 sky130_fd_sc_hd__inv_2 _24161_ (.A(_10263_),
    .Y(_00963_));
 sky130_fd_sc_hd__buf_1 _24162_ (.A(_10079_),
    .X(_10264_));
 sky130_fd_sc_hd__inv_2 _24163_ (.A(_10264_),
    .Y(_00964_));
 sky130_fd_sc_hd__inv_2 _24164_ (.A(_10264_),
    .Y(_00965_));
 sky130_fd_sc_hd__inv_2 _24165_ (.A(_10264_),
    .Y(_00966_));
 sky130_fd_sc_hd__inv_2 _24166_ (.A(_10264_),
    .Y(_00967_));
 sky130_fd_sc_hd__inv_2 _24167_ (.A(_10264_),
    .Y(_00968_));
 sky130_fd_sc_hd__inv_2 _24168_ (.A(_10264_),
    .Y(_00969_));
 sky130_fd_sc_hd__inv_2 _24169_ (.A(_10264_),
    .Y(_00970_));
 sky130_fd_sc_hd__inv_2 _24170_ (.A(_10264_),
    .Y(_00971_));
 sky130_fd_sc_hd__inv_2 _24171_ (.A(_10264_),
    .Y(_00972_));
 sky130_fd_sc_hd__inv_2 _24172_ (.A(_10264_),
    .Y(_00973_));
 sky130_fd_sc_hd__buf_1 _24173_ (.A(_10079_),
    .X(_10265_));
 sky130_fd_sc_hd__inv_2 _24174_ (.A(_10265_),
    .Y(_00974_));
 sky130_fd_sc_hd__inv_2 _24175_ (.A(_10265_),
    .Y(_00975_));
 sky130_fd_sc_hd__inv_2 _24176_ (.A(_10265_),
    .Y(_00976_));
 sky130_fd_sc_hd__inv_2 _24177_ (.A(_10265_),
    .Y(_00977_));
 sky130_fd_sc_hd__inv_2 _24178_ (.A(_10265_),
    .Y(_00978_));
 sky130_fd_sc_hd__inv_2 _24179_ (.A(_10265_),
    .Y(_00979_));
 sky130_fd_sc_hd__inv_2 _24180_ (.A(_10265_),
    .Y(_00980_));
 sky130_fd_sc_hd__inv_2 _24181_ (.A(_10265_),
    .Y(_00981_));
 sky130_fd_sc_hd__inv_2 _24182_ (.A(_10265_),
    .Y(_00982_));
 sky130_fd_sc_hd__inv_2 _24183_ (.A(_10265_),
    .Y(_00983_));
 sky130_fd_sc_hd__buf_1 _24184_ (.A(_10079_),
    .X(_10266_));
 sky130_fd_sc_hd__inv_2 _24185_ (.A(_10266_),
    .Y(_00984_));
 sky130_fd_sc_hd__inv_2 _24186_ (.A(_10266_),
    .Y(_00985_));
 sky130_fd_sc_hd__inv_2 _24187_ (.A(_10266_),
    .Y(_00986_));
 sky130_fd_sc_hd__inv_2 _24188_ (.A(_10266_),
    .Y(_00987_));
 sky130_fd_sc_hd__inv_2 _24189_ (.A(_10266_),
    .Y(_00988_));
 sky130_fd_sc_hd__inv_2 _24190_ (.A(_10266_),
    .Y(_00989_));
 sky130_fd_sc_hd__inv_2 _24191_ (.A(_10266_),
    .Y(_00990_));
 sky130_fd_sc_hd__inv_2 _24192_ (.A(_10266_),
    .Y(_00991_));
 sky130_fd_sc_hd__inv_2 _24193_ (.A(_10266_),
    .Y(_00992_));
 sky130_fd_sc_hd__inv_2 _24194_ (.A(_10266_),
    .Y(_00993_));
 sky130_fd_sc_hd__buf_1 _24195_ (.A(_10079_),
    .X(_10267_));
 sky130_fd_sc_hd__inv_2 _24196_ (.A(_10267_),
    .Y(_00994_));
 sky130_fd_sc_hd__inv_2 _24197_ (.A(_10267_),
    .Y(_00995_));
 sky130_fd_sc_hd__buf_8 _24198_ (.A(_06997_),
    .X(_10268_));
 sky130_fd_sc_hd__buf_8 _24199_ (.A(_09230_),
    .X(_10269_));
 sky130_fd_sc_hd__a21oi_4 _24200_ (.A1(_10268_),
    .A2(_09301_),
    .B1(_10269_),
    .Y(_10270_));
 sky130_fd_sc_hd__mux2_1 _24201_ (.A0(_09298_),
    .A1(\datamem.data_ram[57][24] ),
    .S(_10270_),
    .X(_10271_));
 sky130_fd_sc_hd__clkbuf_1 _24202_ (.A(_10271_),
    .X(_02220_));
 sky130_fd_sc_hd__mux2_1 _24203_ (.A0(_09306_),
    .A1(\datamem.data_ram[57][25] ),
    .S(_10270_),
    .X(_10272_));
 sky130_fd_sc_hd__clkbuf_1 _24204_ (.A(_10272_),
    .X(_02221_));
 sky130_fd_sc_hd__mux2_1 _24205_ (.A0(_09310_),
    .A1(\datamem.data_ram[57][26] ),
    .S(_10270_),
    .X(_10273_));
 sky130_fd_sc_hd__clkbuf_1 _24206_ (.A(_10273_),
    .X(_02222_));
 sky130_fd_sc_hd__mux2_1 _24207_ (.A0(_09314_),
    .A1(\datamem.data_ram[57][27] ),
    .S(_10270_),
    .X(_10274_));
 sky130_fd_sc_hd__clkbuf_1 _24208_ (.A(_10274_),
    .X(_02223_));
 sky130_fd_sc_hd__mux2_1 _24209_ (.A0(_09318_),
    .A1(\datamem.data_ram[57][28] ),
    .S(_10270_),
    .X(_10275_));
 sky130_fd_sc_hd__clkbuf_1 _24210_ (.A(_10275_),
    .X(_02224_));
 sky130_fd_sc_hd__mux2_1 _24211_ (.A0(_09322_),
    .A1(\datamem.data_ram[57][29] ),
    .S(_10270_),
    .X(_10276_));
 sky130_fd_sc_hd__clkbuf_1 _24212_ (.A(_10276_),
    .X(_02225_));
 sky130_fd_sc_hd__mux2_1 _24213_ (.A0(_09326_),
    .A1(\datamem.data_ram[57][30] ),
    .S(_10270_),
    .X(_10277_));
 sky130_fd_sc_hd__clkbuf_1 _24214_ (.A(_10277_),
    .X(_02226_));
 sky130_fd_sc_hd__mux2_1 _24215_ (.A0(_09330_),
    .A1(\datamem.data_ram[57][31] ),
    .S(_10270_),
    .X(_10278_));
 sky130_fd_sc_hd__clkbuf_1 _24216_ (.A(_10278_),
    .X(_02227_));
 sky130_fd_sc_hd__a21oi_4 _24217_ (.A1(_10268_),
    .A2(_09229_),
    .B1(_10269_),
    .Y(_10279_));
 sky130_fd_sc_hd__mux2_1 _24218_ (.A0(_09224_),
    .A1(\datamem.data_ram[57][16] ),
    .S(_10279_),
    .X(_10280_));
 sky130_fd_sc_hd__clkbuf_1 _24219_ (.A(_10280_),
    .X(_02228_));
 sky130_fd_sc_hd__mux2_1 _24220_ (.A0(_09236_),
    .A1(\datamem.data_ram[57][17] ),
    .S(_10279_),
    .X(_10281_));
 sky130_fd_sc_hd__clkbuf_1 _24221_ (.A(_10281_),
    .X(_02229_));
 sky130_fd_sc_hd__mux2_1 _24222_ (.A0(_09240_),
    .A1(\datamem.data_ram[57][18] ),
    .S(_10279_),
    .X(_10282_));
 sky130_fd_sc_hd__clkbuf_1 _24223_ (.A(_10282_),
    .X(_02230_));
 sky130_fd_sc_hd__mux2_1 _24224_ (.A0(_09244_),
    .A1(\datamem.data_ram[57][19] ),
    .S(_10279_),
    .X(_10283_));
 sky130_fd_sc_hd__clkbuf_1 _24225_ (.A(_10283_),
    .X(_02231_));
 sky130_fd_sc_hd__mux2_1 _24226_ (.A0(_09248_),
    .A1(\datamem.data_ram[57][20] ),
    .S(_10279_),
    .X(_10284_));
 sky130_fd_sc_hd__clkbuf_1 _24227_ (.A(_10284_),
    .X(_02232_));
 sky130_fd_sc_hd__mux2_1 _24228_ (.A0(_09252_),
    .A1(\datamem.data_ram[57][21] ),
    .S(_10279_),
    .X(_10285_));
 sky130_fd_sc_hd__clkbuf_1 _24229_ (.A(_10285_),
    .X(_02233_));
 sky130_fd_sc_hd__mux2_1 _24230_ (.A0(_09256_),
    .A1(\datamem.data_ram[57][22] ),
    .S(_10279_),
    .X(_10286_));
 sky130_fd_sc_hd__clkbuf_1 _24231_ (.A(_10286_),
    .X(_02234_));
 sky130_fd_sc_hd__mux2_1 _24232_ (.A0(_09260_),
    .A1(\datamem.data_ram[57][23] ),
    .S(_10279_),
    .X(_10287_));
 sky130_fd_sc_hd__clkbuf_1 _24233_ (.A(_10287_),
    .X(_02235_));
 sky130_fd_sc_hd__a21oi_4 _24234_ (.A1(_10268_),
    .A2(_09269_),
    .B1(_10269_),
    .Y(_10288_));
 sky130_fd_sc_hd__mux2_1 _24235_ (.A0(_09267_),
    .A1(\datamem.data_ram[57][8] ),
    .S(_10288_),
    .X(_10289_));
 sky130_fd_sc_hd__clkbuf_1 _24236_ (.A(_10289_),
    .X(_02236_));
 sky130_fd_sc_hd__mux2_1 _24237_ (.A0(_09273_),
    .A1(\datamem.data_ram[57][9] ),
    .S(_10288_),
    .X(_10290_));
 sky130_fd_sc_hd__clkbuf_1 _24238_ (.A(_10290_),
    .X(_02237_));
 sky130_fd_sc_hd__mux2_1 _24239_ (.A0(_09276_),
    .A1(\datamem.data_ram[57][10] ),
    .S(_10288_),
    .X(_10291_));
 sky130_fd_sc_hd__clkbuf_1 _24240_ (.A(_10291_),
    .X(_02238_));
 sky130_fd_sc_hd__mux2_1 _24241_ (.A0(_09279_),
    .A1(\datamem.data_ram[57][11] ),
    .S(_10288_),
    .X(_10292_));
 sky130_fd_sc_hd__clkbuf_1 _24242_ (.A(_10292_),
    .X(_02239_));
 sky130_fd_sc_hd__mux2_1 _24243_ (.A0(_09282_),
    .A1(\datamem.data_ram[57][12] ),
    .S(_10288_),
    .X(_10293_));
 sky130_fd_sc_hd__clkbuf_1 _24244_ (.A(_10293_),
    .X(_02240_));
 sky130_fd_sc_hd__mux2_1 _24245_ (.A0(_09285_),
    .A1(\datamem.data_ram[57][13] ),
    .S(_10288_),
    .X(_10294_));
 sky130_fd_sc_hd__clkbuf_1 _24246_ (.A(_10294_),
    .X(_02241_));
 sky130_fd_sc_hd__mux2_1 _24247_ (.A0(_09288_),
    .A1(\datamem.data_ram[57][14] ),
    .S(_10288_),
    .X(_10295_));
 sky130_fd_sc_hd__clkbuf_1 _24248_ (.A(_10295_),
    .X(_02242_));
 sky130_fd_sc_hd__mux2_1 _24249_ (.A0(_09291_),
    .A1(\datamem.data_ram[57][15] ),
    .S(_10288_),
    .X(_10296_));
 sky130_fd_sc_hd__clkbuf_1 _24250_ (.A(_10296_),
    .X(_02243_));
 sky130_fd_sc_hd__buf_8 _24251_ (.A(_07122_),
    .X(_10297_));
 sky130_fd_sc_hd__a21oi_4 _24252_ (.A1(_10297_),
    .A2(_09301_),
    .B1(_10269_),
    .Y(_10298_));
 sky130_fd_sc_hd__mux2_1 _24253_ (.A0(_09298_),
    .A1(\datamem.data_ram[56][24] ),
    .S(_10298_),
    .X(_10299_));
 sky130_fd_sc_hd__clkbuf_1 _24254_ (.A(_10299_),
    .X(_02244_));
 sky130_fd_sc_hd__mux2_1 _24255_ (.A0(_09306_),
    .A1(\datamem.data_ram[56][25] ),
    .S(_10298_),
    .X(_10300_));
 sky130_fd_sc_hd__clkbuf_1 _24256_ (.A(_10300_),
    .X(_02245_));
 sky130_fd_sc_hd__mux2_1 _24257_ (.A0(_09310_),
    .A1(\datamem.data_ram[56][26] ),
    .S(_10298_),
    .X(_10301_));
 sky130_fd_sc_hd__clkbuf_1 _24258_ (.A(_10301_),
    .X(_02246_));
 sky130_fd_sc_hd__mux2_1 _24259_ (.A0(_09314_),
    .A1(\datamem.data_ram[56][27] ),
    .S(_10298_),
    .X(_10302_));
 sky130_fd_sc_hd__clkbuf_1 _24260_ (.A(_10302_),
    .X(_02247_));
 sky130_fd_sc_hd__mux2_1 _24261_ (.A0(_09318_),
    .A1(\datamem.data_ram[56][28] ),
    .S(_10298_),
    .X(_10303_));
 sky130_fd_sc_hd__clkbuf_1 _24262_ (.A(_10303_),
    .X(_02248_));
 sky130_fd_sc_hd__mux2_1 _24263_ (.A0(_09322_),
    .A1(\datamem.data_ram[56][29] ),
    .S(_10298_),
    .X(_10304_));
 sky130_fd_sc_hd__clkbuf_1 _24264_ (.A(_10304_),
    .X(_02249_));
 sky130_fd_sc_hd__mux2_1 _24265_ (.A0(_09326_),
    .A1(\datamem.data_ram[56][30] ),
    .S(_10298_),
    .X(_10305_));
 sky130_fd_sc_hd__clkbuf_1 _24266_ (.A(_10305_),
    .X(_02250_));
 sky130_fd_sc_hd__mux2_1 _24267_ (.A0(_09330_),
    .A1(\datamem.data_ram[56][31] ),
    .S(_10298_),
    .X(_10306_));
 sky130_fd_sc_hd__clkbuf_1 _24268_ (.A(_10306_),
    .X(_02251_));
 sky130_fd_sc_hd__a21oi_4 _24269_ (.A1(_10297_),
    .A2(_09229_),
    .B1(_10269_),
    .Y(_10307_));
 sky130_fd_sc_hd__mux2_1 _24270_ (.A0(_09224_),
    .A1(\datamem.data_ram[56][16] ),
    .S(_10307_),
    .X(_10308_));
 sky130_fd_sc_hd__clkbuf_1 _24271_ (.A(_10308_),
    .X(_02252_));
 sky130_fd_sc_hd__mux2_1 _24272_ (.A0(_09236_),
    .A1(\datamem.data_ram[56][17] ),
    .S(_10307_),
    .X(_10309_));
 sky130_fd_sc_hd__clkbuf_1 _24273_ (.A(_10309_),
    .X(_02253_));
 sky130_fd_sc_hd__mux2_1 _24274_ (.A0(_09240_),
    .A1(\datamem.data_ram[56][18] ),
    .S(_10307_),
    .X(_10310_));
 sky130_fd_sc_hd__clkbuf_1 _24275_ (.A(_10310_),
    .X(_02254_));
 sky130_fd_sc_hd__mux2_1 _24276_ (.A0(_09244_),
    .A1(\datamem.data_ram[56][19] ),
    .S(_10307_),
    .X(_10311_));
 sky130_fd_sc_hd__clkbuf_1 _24277_ (.A(_10311_),
    .X(_02255_));
 sky130_fd_sc_hd__mux2_1 _24278_ (.A0(_09248_),
    .A1(\datamem.data_ram[56][20] ),
    .S(_10307_),
    .X(_10312_));
 sky130_fd_sc_hd__clkbuf_1 _24279_ (.A(_10312_),
    .X(_02256_));
 sky130_fd_sc_hd__mux2_1 _24280_ (.A0(_09252_),
    .A1(\datamem.data_ram[56][21] ),
    .S(_10307_),
    .X(_10313_));
 sky130_fd_sc_hd__clkbuf_1 _24281_ (.A(_10313_),
    .X(_02257_));
 sky130_fd_sc_hd__mux2_1 _24282_ (.A0(_09256_),
    .A1(\datamem.data_ram[56][22] ),
    .S(_10307_),
    .X(_10314_));
 sky130_fd_sc_hd__clkbuf_1 _24283_ (.A(_10314_),
    .X(_02258_));
 sky130_fd_sc_hd__mux2_1 _24284_ (.A0(_09260_),
    .A1(\datamem.data_ram[56][23] ),
    .S(_10307_),
    .X(_10315_));
 sky130_fd_sc_hd__clkbuf_1 _24285_ (.A(_10315_),
    .X(_02259_));
 sky130_fd_sc_hd__a21oi_4 _24286_ (.A1(_10297_),
    .A2(_09269_),
    .B1(_10269_),
    .Y(_10316_));
 sky130_fd_sc_hd__mux2_1 _24287_ (.A0(_09267_),
    .A1(\datamem.data_ram[56][8] ),
    .S(_10316_),
    .X(_10317_));
 sky130_fd_sc_hd__clkbuf_1 _24288_ (.A(_10317_),
    .X(_02260_));
 sky130_fd_sc_hd__mux2_1 _24289_ (.A0(_09273_),
    .A1(\datamem.data_ram[56][9] ),
    .S(_10316_),
    .X(_10318_));
 sky130_fd_sc_hd__clkbuf_1 _24290_ (.A(_10318_),
    .X(_02261_));
 sky130_fd_sc_hd__mux2_1 _24291_ (.A0(_09276_),
    .A1(\datamem.data_ram[56][10] ),
    .S(_10316_),
    .X(_10319_));
 sky130_fd_sc_hd__clkbuf_1 _24292_ (.A(_10319_),
    .X(_02262_));
 sky130_fd_sc_hd__mux2_1 _24293_ (.A0(_09279_),
    .A1(\datamem.data_ram[56][11] ),
    .S(_10316_),
    .X(_10320_));
 sky130_fd_sc_hd__clkbuf_1 _24294_ (.A(_10320_),
    .X(_02263_));
 sky130_fd_sc_hd__mux2_1 _24295_ (.A0(_09282_),
    .A1(\datamem.data_ram[56][12] ),
    .S(_10316_),
    .X(_10321_));
 sky130_fd_sc_hd__clkbuf_1 _24296_ (.A(_10321_),
    .X(_02264_));
 sky130_fd_sc_hd__mux2_1 _24297_ (.A0(_09285_),
    .A1(\datamem.data_ram[56][13] ),
    .S(_10316_),
    .X(_10322_));
 sky130_fd_sc_hd__clkbuf_1 _24298_ (.A(_10322_),
    .X(_02265_));
 sky130_fd_sc_hd__mux2_1 _24299_ (.A0(_09288_),
    .A1(\datamem.data_ram[56][14] ),
    .S(_10316_),
    .X(_10323_));
 sky130_fd_sc_hd__clkbuf_1 _24300_ (.A(_10323_),
    .X(_02266_));
 sky130_fd_sc_hd__mux2_1 _24301_ (.A0(_09291_),
    .A1(\datamem.data_ram[56][15] ),
    .S(_10316_),
    .X(_10324_));
 sky130_fd_sc_hd__clkbuf_1 _24302_ (.A(_10324_),
    .X(_02267_));
 sky130_fd_sc_hd__buf_6 _24303_ (.A(_07125_),
    .X(_10325_));
 sky130_fd_sc_hd__nand2_8 _24304_ (.A(_06681_),
    .B(_08355_),
    .Y(_10326_));
 sky130_fd_sc_hd__nor2_8 _24305_ (.A(_10326_),
    .B(net107),
    .Y(_10327_));
 sky130_fd_sc_hd__a21oi_4 _24306_ (.A1(_10325_),
    .A2(_10327_),
    .B1(_10269_),
    .Y(_10328_));
 sky130_fd_sc_hd__mux2_1 _24307_ (.A0(_09298_),
    .A1(\datamem.data_ram[55][24] ),
    .S(_10328_),
    .X(_10329_));
 sky130_fd_sc_hd__clkbuf_1 _24308_ (.A(_10329_),
    .X(_02268_));
 sky130_fd_sc_hd__mux2_1 _24309_ (.A0(_09306_),
    .A1(\datamem.data_ram[55][25] ),
    .S(_10328_),
    .X(_10330_));
 sky130_fd_sc_hd__clkbuf_1 _24310_ (.A(_10330_),
    .X(_02269_));
 sky130_fd_sc_hd__mux2_1 _24311_ (.A0(_09310_),
    .A1(\datamem.data_ram[55][26] ),
    .S(_10328_),
    .X(_10331_));
 sky130_fd_sc_hd__clkbuf_1 _24312_ (.A(_10331_),
    .X(_02270_));
 sky130_fd_sc_hd__mux2_1 _24313_ (.A0(_09314_),
    .A1(\datamem.data_ram[55][27] ),
    .S(_10328_),
    .X(_10332_));
 sky130_fd_sc_hd__clkbuf_1 _24314_ (.A(_10332_),
    .X(_02271_));
 sky130_fd_sc_hd__mux2_1 _24315_ (.A0(_09318_),
    .A1(\datamem.data_ram[55][28] ),
    .S(_10328_),
    .X(_10333_));
 sky130_fd_sc_hd__clkbuf_1 _24316_ (.A(_10333_),
    .X(_02272_));
 sky130_fd_sc_hd__mux2_1 _24317_ (.A0(_09322_),
    .A1(\datamem.data_ram[55][29] ),
    .S(_10328_),
    .X(_10334_));
 sky130_fd_sc_hd__clkbuf_1 _24318_ (.A(_10334_),
    .X(_02273_));
 sky130_fd_sc_hd__mux2_1 _24319_ (.A0(_09326_),
    .A1(\datamem.data_ram[55][30] ),
    .S(_10328_),
    .X(_10335_));
 sky130_fd_sc_hd__clkbuf_1 _24320_ (.A(_10335_),
    .X(_02274_));
 sky130_fd_sc_hd__mux2_1 _24321_ (.A0(_09330_),
    .A1(\datamem.data_ram[55][31] ),
    .S(_10328_),
    .X(_10336_));
 sky130_fd_sc_hd__clkbuf_1 _24322_ (.A(_10336_),
    .X(_02275_));
 sky130_fd_sc_hd__nor2_8 _24323_ (.A(_10326_),
    .B(net104),
    .Y(_10337_));
 sky130_fd_sc_hd__a21oi_4 _24324_ (.A1(_10325_),
    .A2(_10337_),
    .B1(_10269_),
    .Y(_10338_));
 sky130_fd_sc_hd__mux2_1 _24325_ (.A0(_09224_),
    .A1(\datamem.data_ram[55][16] ),
    .S(_10338_),
    .X(_10339_));
 sky130_fd_sc_hd__clkbuf_1 _24326_ (.A(_10339_),
    .X(_02276_));
 sky130_fd_sc_hd__mux2_1 _24327_ (.A0(_09236_),
    .A1(\datamem.data_ram[55][17] ),
    .S(_10338_),
    .X(_10340_));
 sky130_fd_sc_hd__clkbuf_1 _24328_ (.A(_10340_),
    .X(_02277_));
 sky130_fd_sc_hd__mux2_1 _24329_ (.A0(_09240_),
    .A1(\datamem.data_ram[55][18] ),
    .S(_10338_),
    .X(_10341_));
 sky130_fd_sc_hd__clkbuf_1 _24330_ (.A(_10341_),
    .X(_02278_));
 sky130_fd_sc_hd__mux2_1 _24331_ (.A0(_09244_),
    .A1(\datamem.data_ram[55][19] ),
    .S(_10338_),
    .X(_10342_));
 sky130_fd_sc_hd__clkbuf_1 _24332_ (.A(_10342_),
    .X(_02279_));
 sky130_fd_sc_hd__mux2_1 _24333_ (.A0(_09248_),
    .A1(\datamem.data_ram[55][20] ),
    .S(_10338_),
    .X(_10343_));
 sky130_fd_sc_hd__clkbuf_1 _24334_ (.A(_10343_),
    .X(_02280_));
 sky130_fd_sc_hd__mux2_1 _24335_ (.A0(_09252_),
    .A1(\datamem.data_ram[55][21] ),
    .S(_10338_),
    .X(_10344_));
 sky130_fd_sc_hd__clkbuf_1 _24336_ (.A(_10344_),
    .X(_02281_));
 sky130_fd_sc_hd__mux2_1 _24337_ (.A0(_09256_),
    .A1(\datamem.data_ram[55][22] ),
    .S(_10338_),
    .X(_10345_));
 sky130_fd_sc_hd__clkbuf_1 _24338_ (.A(_10345_),
    .X(_02282_));
 sky130_fd_sc_hd__mux2_1 _24339_ (.A0(_09260_),
    .A1(\datamem.data_ram[55][23] ),
    .S(_10338_),
    .X(_10346_));
 sky130_fd_sc_hd__clkbuf_1 _24340_ (.A(_10346_),
    .X(_02283_));
 sky130_fd_sc_hd__nor2_8 _24341_ (.A(_10326_),
    .B(net112),
    .Y(_10347_));
 sky130_fd_sc_hd__a21oi_4 _24342_ (.A1(_10325_),
    .A2(_10347_),
    .B1(_10269_),
    .Y(_10348_));
 sky130_fd_sc_hd__mux2_1 _24343_ (.A0(_09267_),
    .A1(\datamem.data_ram[55][8] ),
    .S(_10348_),
    .X(_10349_));
 sky130_fd_sc_hd__clkbuf_1 _24344_ (.A(_10349_),
    .X(_02284_));
 sky130_fd_sc_hd__mux2_1 _24345_ (.A0(_09273_),
    .A1(\datamem.data_ram[55][9] ),
    .S(_10348_),
    .X(_10350_));
 sky130_fd_sc_hd__clkbuf_1 _24346_ (.A(_10350_),
    .X(_02285_));
 sky130_fd_sc_hd__mux2_1 _24347_ (.A0(_09276_),
    .A1(\datamem.data_ram[55][10] ),
    .S(_10348_),
    .X(_10351_));
 sky130_fd_sc_hd__clkbuf_1 _24348_ (.A(_10351_),
    .X(_02286_));
 sky130_fd_sc_hd__mux2_1 _24349_ (.A0(_09279_),
    .A1(\datamem.data_ram[55][11] ),
    .S(_10348_),
    .X(_10352_));
 sky130_fd_sc_hd__clkbuf_1 _24350_ (.A(_10352_),
    .X(_02287_));
 sky130_fd_sc_hd__mux2_1 _24351_ (.A0(_09282_),
    .A1(\datamem.data_ram[55][12] ),
    .S(_10348_),
    .X(_10353_));
 sky130_fd_sc_hd__clkbuf_1 _24352_ (.A(_10353_),
    .X(_02288_));
 sky130_fd_sc_hd__mux2_1 _24353_ (.A0(_09285_),
    .A1(\datamem.data_ram[55][13] ),
    .S(_10348_),
    .X(_10354_));
 sky130_fd_sc_hd__clkbuf_1 _24354_ (.A(_10354_),
    .X(_02289_));
 sky130_fd_sc_hd__mux2_1 _24355_ (.A0(_09288_),
    .A1(\datamem.data_ram[55][14] ),
    .S(_10348_),
    .X(_10355_));
 sky130_fd_sc_hd__clkbuf_1 _24356_ (.A(_10355_),
    .X(_02290_));
 sky130_fd_sc_hd__mux2_1 _24357_ (.A0(_09291_),
    .A1(\datamem.data_ram[55][15] ),
    .S(_10348_),
    .X(_10356_));
 sky130_fd_sc_hd__clkbuf_1 _24358_ (.A(_10356_),
    .X(_02291_));
 sky130_fd_sc_hd__a21oi_2 _24359_ (.A1(_09226_),
    .A2(_10327_),
    .B1(_10269_),
    .Y(_10357_));
 sky130_fd_sc_hd__mux2_1 _24360_ (.A0(_09298_),
    .A1(\datamem.data_ram[54][24] ),
    .S(net61),
    .X(_10358_));
 sky130_fd_sc_hd__clkbuf_1 _24361_ (.A(_10358_),
    .X(_02292_));
 sky130_fd_sc_hd__mux2_1 _24362_ (.A0(_09306_),
    .A1(\datamem.data_ram[54][25] ),
    .S(net61),
    .X(_10359_));
 sky130_fd_sc_hd__clkbuf_1 _24363_ (.A(_10359_),
    .X(_02293_));
 sky130_fd_sc_hd__mux2_1 _24364_ (.A0(_09310_),
    .A1(\datamem.data_ram[54][26] ),
    .S(_10357_),
    .X(_10360_));
 sky130_fd_sc_hd__clkbuf_1 _24365_ (.A(_10360_),
    .X(_02294_));
 sky130_fd_sc_hd__mux2_1 _24366_ (.A0(_09314_),
    .A1(\datamem.data_ram[54][27] ),
    .S(net61),
    .X(_10361_));
 sky130_fd_sc_hd__clkbuf_1 _24367_ (.A(_10361_),
    .X(_02295_));
 sky130_fd_sc_hd__mux2_1 _24368_ (.A0(_09318_),
    .A1(\datamem.data_ram[54][28] ),
    .S(net61),
    .X(_10362_));
 sky130_fd_sc_hd__clkbuf_1 _24369_ (.A(_10362_),
    .X(_02296_));
 sky130_fd_sc_hd__mux2_1 _24370_ (.A0(_09322_),
    .A1(\datamem.data_ram[54][29] ),
    .S(net61),
    .X(_10363_));
 sky130_fd_sc_hd__clkbuf_1 _24371_ (.A(_10363_),
    .X(_02297_));
 sky130_fd_sc_hd__mux2_1 _24372_ (.A0(_09326_),
    .A1(\datamem.data_ram[54][30] ),
    .S(net61),
    .X(_10364_));
 sky130_fd_sc_hd__clkbuf_1 _24373_ (.A(_10364_),
    .X(_02298_));
 sky130_fd_sc_hd__mux2_1 _24374_ (.A0(_09330_),
    .A1(\datamem.data_ram[54][31] ),
    .S(_10357_),
    .X(_10365_));
 sky130_fd_sc_hd__clkbuf_1 _24375_ (.A(_10365_),
    .X(_02299_));
 sky130_fd_sc_hd__buf_8 _24376_ (.A(_09230_),
    .X(_10366_));
 sky130_fd_sc_hd__a21oi_4 _24377_ (.A1(_09226_),
    .A2(_10337_),
    .B1(_10366_),
    .Y(_10367_));
 sky130_fd_sc_hd__mux2_1 _24378_ (.A0(_09224_),
    .A1(\datamem.data_ram[54][16] ),
    .S(_10367_),
    .X(_10368_));
 sky130_fd_sc_hd__clkbuf_1 _24379_ (.A(_10368_),
    .X(_02300_));
 sky130_fd_sc_hd__mux2_1 _24380_ (.A0(_09236_),
    .A1(\datamem.data_ram[54][17] ),
    .S(_10367_),
    .X(_10369_));
 sky130_fd_sc_hd__clkbuf_1 _24381_ (.A(_10369_),
    .X(_02301_));
 sky130_fd_sc_hd__mux2_1 _24382_ (.A0(_09240_),
    .A1(\datamem.data_ram[54][18] ),
    .S(_10367_),
    .X(_10370_));
 sky130_fd_sc_hd__clkbuf_1 _24383_ (.A(_10370_),
    .X(_02302_));
 sky130_fd_sc_hd__mux2_1 _24384_ (.A0(_09244_),
    .A1(\datamem.data_ram[54][19] ),
    .S(_10367_),
    .X(_10371_));
 sky130_fd_sc_hd__clkbuf_1 _24385_ (.A(_10371_),
    .X(_02303_));
 sky130_fd_sc_hd__mux2_1 _24386_ (.A0(_09248_),
    .A1(\datamem.data_ram[54][20] ),
    .S(_10367_),
    .X(_10372_));
 sky130_fd_sc_hd__clkbuf_1 _24387_ (.A(_10372_),
    .X(_02304_));
 sky130_fd_sc_hd__mux2_1 _24388_ (.A0(_09252_),
    .A1(\datamem.data_ram[54][21] ),
    .S(_10367_),
    .X(_10373_));
 sky130_fd_sc_hd__clkbuf_1 _24389_ (.A(_10373_),
    .X(_02305_));
 sky130_fd_sc_hd__mux2_1 _24390_ (.A0(_09256_),
    .A1(\datamem.data_ram[54][22] ),
    .S(_10367_),
    .X(_10374_));
 sky130_fd_sc_hd__clkbuf_1 _24391_ (.A(_10374_),
    .X(_02306_));
 sky130_fd_sc_hd__mux2_1 _24392_ (.A0(_09260_),
    .A1(\datamem.data_ram[54][23] ),
    .S(_10367_),
    .X(_10375_));
 sky130_fd_sc_hd__clkbuf_1 _24393_ (.A(_10375_),
    .X(_02307_));
 sky130_fd_sc_hd__a21oi_4 _24394_ (.A1(_09226_),
    .A2(_10347_),
    .B1(_10366_),
    .Y(_10376_));
 sky130_fd_sc_hd__mux2_1 _24395_ (.A0(_09267_),
    .A1(\datamem.data_ram[54][8] ),
    .S(_10376_),
    .X(_10377_));
 sky130_fd_sc_hd__clkbuf_1 _24396_ (.A(_10377_),
    .X(_02308_));
 sky130_fd_sc_hd__mux2_1 _24397_ (.A0(_09273_),
    .A1(\datamem.data_ram[54][9] ),
    .S(_10376_),
    .X(_10378_));
 sky130_fd_sc_hd__clkbuf_1 _24398_ (.A(_10378_),
    .X(_02309_));
 sky130_fd_sc_hd__mux2_1 _24399_ (.A0(_09276_),
    .A1(\datamem.data_ram[54][10] ),
    .S(_10376_),
    .X(_10379_));
 sky130_fd_sc_hd__clkbuf_1 _24400_ (.A(_10379_),
    .X(_02310_));
 sky130_fd_sc_hd__mux2_1 _24401_ (.A0(_09279_),
    .A1(\datamem.data_ram[54][11] ),
    .S(_10376_),
    .X(_10380_));
 sky130_fd_sc_hd__clkbuf_1 _24402_ (.A(_10380_),
    .X(_02311_));
 sky130_fd_sc_hd__mux2_1 _24403_ (.A0(_09282_),
    .A1(\datamem.data_ram[54][12] ),
    .S(_10376_),
    .X(_10381_));
 sky130_fd_sc_hd__clkbuf_1 _24404_ (.A(_10381_),
    .X(_02312_));
 sky130_fd_sc_hd__mux2_1 _24405_ (.A0(_09285_),
    .A1(\datamem.data_ram[54][13] ),
    .S(_10376_),
    .X(_10382_));
 sky130_fd_sc_hd__clkbuf_1 _24406_ (.A(_10382_),
    .X(_02313_));
 sky130_fd_sc_hd__mux2_1 _24407_ (.A0(_09288_),
    .A1(\datamem.data_ram[54][14] ),
    .S(_10376_),
    .X(_10383_));
 sky130_fd_sc_hd__clkbuf_1 _24408_ (.A(_10383_),
    .X(_02314_));
 sky130_fd_sc_hd__mux2_1 _24409_ (.A0(_09291_),
    .A1(\datamem.data_ram[54][15] ),
    .S(_10376_),
    .X(_10384_));
 sky130_fd_sc_hd__clkbuf_1 _24410_ (.A(_10384_),
    .X(_02315_));
 sky130_fd_sc_hd__buf_2 _24411_ (.A(_09266_),
    .X(_10385_));
 sky130_fd_sc_hd__a21oi_4 _24412_ (.A1(_10113_),
    .A2(_10347_),
    .B1(_10366_),
    .Y(_10386_));
 sky130_fd_sc_hd__mux2_1 _24413_ (.A0(_10385_),
    .A1(\datamem.data_ram[53][8] ),
    .S(_10386_),
    .X(_10387_));
 sky130_fd_sc_hd__clkbuf_1 _24414_ (.A(_10387_),
    .X(_02316_));
 sky130_fd_sc_hd__buf_2 _24415_ (.A(_09272_),
    .X(_10388_));
 sky130_fd_sc_hd__mux2_1 _24416_ (.A0(_10388_),
    .A1(\datamem.data_ram[53][9] ),
    .S(_10386_),
    .X(_10389_));
 sky130_fd_sc_hd__clkbuf_1 _24417_ (.A(_10389_),
    .X(_02317_));
 sky130_fd_sc_hd__buf_2 _24418_ (.A(_09275_),
    .X(_10390_));
 sky130_fd_sc_hd__mux2_1 _24419_ (.A0(_10390_),
    .A1(\datamem.data_ram[53][10] ),
    .S(_10386_),
    .X(_10391_));
 sky130_fd_sc_hd__clkbuf_1 _24420_ (.A(_10391_),
    .X(_02318_));
 sky130_fd_sc_hd__clkbuf_4 _24421_ (.A(_09278_),
    .X(_10392_));
 sky130_fd_sc_hd__mux2_1 _24422_ (.A0(_10392_),
    .A1(\datamem.data_ram[53][11] ),
    .S(_10386_),
    .X(_10393_));
 sky130_fd_sc_hd__clkbuf_1 _24423_ (.A(_10393_),
    .X(_02319_));
 sky130_fd_sc_hd__buf_2 _24424_ (.A(_09281_),
    .X(_10394_));
 sky130_fd_sc_hd__mux2_1 _24425_ (.A0(_10394_),
    .A1(\datamem.data_ram[53][12] ),
    .S(_10386_),
    .X(_10395_));
 sky130_fd_sc_hd__clkbuf_1 _24426_ (.A(_10395_),
    .X(_02320_));
 sky130_fd_sc_hd__buf_2 _24427_ (.A(_09284_),
    .X(_10396_));
 sky130_fd_sc_hd__mux2_1 _24428_ (.A0(_10396_),
    .A1(\datamem.data_ram[53][13] ),
    .S(_10386_),
    .X(_10397_));
 sky130_fd_sc_hd__clkbuf_1 _24429_ (.A(_10397_),
    .X(_02321_));
 sky130_fd_sc_hd__buf_2 _24430_ (.A(_09287_),
    .X(_10398_));
 sky130_fd_sc_hd__mux2_1 _24431_ (.A0(_10398_),
    .A1(\datamem.data_ram[53][14] ),
    .S(_10386_),
    .X(_10399_));
 sky130_fd_sc_hd__clkbuf_1 _24432_ (.A(_10399_),
    .X(_02322_));
 sky130_fd_sc_hd__buf_2 _24433_ (.A(_09290_),
    .X(_10400_));
 sky130_fd_sc_hd__mux2_1 _24434_ (.A0(_10400_),
    .A1(\datamem.data_ram[53][15] ),
    .S(_10386_),
    .X(_10401_));
 sky130_fd_sc_hd__clkbuf_1 _24435_ (.A(_10401_),
    .X(_02323_));
 sky130_fd_sc_hd__buf_2 _24436_ (.A(_10326_),
    .X(_10402_));
 sky130_fd_sc_hd__or3_1 _24437_ (.A(_07019_),
    .B(_10402_),
    .C(_10044_),
    .X(_10403_));
 sky130_fd_sc_hd__clkbuf_2 _24438_ (.A(_10403_),
    .X(_10404_));
 sky130_fd_sc_hd__clkbuf_4 _24439_ (.A(_10047_),
    .X(_10405_));
 sky130_fd_sc_hd__and3_1 _24440_ (.A(_09299_),
    .B(_08059_),
    .C(_10052_),
    .X(_10406_));
 sky130_fd_sc_hd__and2_1 _24441_ (.A(_10405_),
    .B(_10406_),
    .X(_10407_));
 sky130_fd_sc_hd__a31o_1 _24442_ (.A1(_10056_),
    .A2(\datamem.data_ram[53][0] ),
    .A3(_10404_),
    .B1(_10407_),
    .X(_02324_));
 sky130_fd_sc_hd__buf_2 _24443_ (.A(_10057_),
    .X(_10408_));
 sky130_fd_sc_hd__and2_1 _24444_ (.A(_10408_),
    .B(_10406_),
    .X(_10409_));
 sky130_fd_sc_hd__a31o_1 _24445_ (.A1(_10056_),
    .A2(\datamem.data_ram[53][1] ),
    .A3(_10404_),
    .B1(_10409_),
    .X(_02325_));
 sky130_fd_sc_hd__clkbuf_4 _24446_ (.A(_10060_),
    .X(_10410_));
 sky130_fd_sc_hd__and2_1 _24447_ (.A(_10410_),
    .B(_10406_),
    .X(_10411_));
 sky130_fd_sc_hd__a31o_1 _24448_ (.A1(_10056_),
    .A2(\datamem.data_ram[53][2] ),
    .A3(_10404_),
    .B1(_10411_),
    .X(_02326_));
 sky130_fd_sc_hd__clkbuf_4 _24449_ (.A(_10055_),
    .X(_10412_));
 sky130_fd_sc_hd__buf_2 _24450_ (.A(_10063_),
    .X(_10413_));
 sky130_fd_sc_hd__and2_1 _24451_ (.A(_10413_),
    .B(_10406_),
    .X(_10414_));
 sky130_fd_sc_hd__a31o_1 _24452_ (.A1(_10412_),
    .A2(\datamem.data_ram[53][3] ),
    .A3(_10404_),
    .B1(_10414_),
    .X(_02327_));
 sky130_fd_sc_hd__and2_1 _24453_ (.A(_10067_),
    .B(_10406_),
    .X(_10415_));
 sky130_fd_sc_hd__a31o_1 _24454_ (.A1(_10412_),
    .A2(\datamem.data_ram[53][4] ),
    .A3(_10404_),
    .B1(_10415_),
    .X(_02328_));
 sky130_fd_sc_hd__buf_2 _24455_ (.A(_10069_),
    .X(_10416_));
 sky130_fd_sc_hd__and2_1 _24456_ (.A(_10416_),
    .B(_10406_),
    .X(_10417_));
 sky130_fd_sc_hd__a31o_1 _24457_ (.A1(_10412_),
    .A2(\datamem.data_ram[53][5] ),
    .A3(_10404_),
    .B1(_10417_),
    .X(_02329_));
 sky130_fd_sc_hd__clkbuf_4 _24458_ (.A(_10072_),
    .X(_10418_));
 sky130_fd_sc_hd__and2_1 _24459_ (.A(_10418_),
    .B(_10406_),
    .X(_10419_));
 sky130_fd_sc_hd__a31o_1 _24460_ (.A1(_10412_),
    .A2(\datamem.data_ram[53][6] ),
    .A3(_10404_),
    .B1(_10419_),
    .X(_02330_));
 sky130_fd_sc_hd__and2_1 _24461_ (.A(_10076_),
    .B(_10406_),
    .X(_10420_));
 sky130_fd_sc_hd__a31o_1 _24462_ (.A1(_10412_),
    .A2(\datamem.data_ram[53][7] ),
    .A3(_10404_),
    .B1(_10420_),
    .X(_02331_));
 sky130_fd_sc_hd__a21oi_4 _24463_ (.A1(_10113_),
    .A2(_10327_),
    .B1(_10366_),
    .Y(_10421_));
 sky130_fd_sc_hd__mux2_1 _24464_ (.A0(_09298_),
    .A1(\datamem.data_ram[53][24] ),
    .S(_10421_),
    .X(_10422_));
 sky130_fd_sc_hd__clkbuf_1 _24465_ (.A(_10422_),
    .X(_02332_));
 sky130_fd_sc_hd__mux2_1 _24466_ (.A0(_09306_),
    .A1(\datamem.data_ram[53][25] ),
    .S(_10421_),
    .X(_10423_));
 sky130_fd_sc_hd__clkbuf_1 _24467_ (.A(_10423_),
    .X(_02333_));
 sky130_fd_sc_hd__mux2_1 _24468_ (.A0(_09310_),
    .A1(\datamem.data_ram[53][26] ),
    .S(_10421_),
    .X(_10424_));
 sky130_fd_sc_hd__clkbuf_1 _24469_ (.A(_10424_),
    .X(_02334_));
 sky130_fd_sc_hd__mux2_1 _24470_ (.A0(_09314_),
    .A1(\datamem.data_ram[53][27] ),
    .S(_10421_),
    .X(_10425_));
 sky130_fd_sc_hd__clkbuf_1 _24471_ (.A(_10425_),
    .X(_02335_));
 sky130_fd_sc_hd__mux2_1 _24472_ (.A0(_09318_),
    .A1(\datamem.data_ram[53][28] ),
    .S(_10421_),
    .X(_10426_));
 sky130_fd_sc_hd__clkbuf_1 _24473_ (.A(_10426_),
    .X(_02336_));
 sky130_fd_sc_hd__mux2_1 _24474_ (.A0(_09322_),
    .A1(\datamem.data_ram[53][29] ),
    .S(_10421_),
    .X(_10427_));
 sky130_fd_sc_hd__clkbuf_1 _24475_ (.A(_10427_),
    .X(_02337_));
 sky130_fd_sc_hd__mux2_1 _24476_ (.A0(_09326_),
    .A1(\datamem.data_ram[53][30] ),
    .S(_10421_),
    .X(_10428_));
 sky130_fd_sc_hd__clkbuf_1 _24477_ (.A(_10428_),
    .X(_02338_));
 sky130_fd_sc_hd__mux2_1 _24478_ (.A0(_09330_),
    .A1(\datamem.data_ram[53][31] ),
    .S(_10421_),
    .X(_10429_));
 sky130_fd_sc_hd__clkbuf_1 _24479_ (.A(_10429_),
    .X(_02339_));
 sky130_fd_sc_hd__a21oi_4 _24480_ (.A1(_09351_),
    .A2(_10327_),
    .B1(_10366_),
    .Y(_10430_));
 sky130_fd_sc_hd__mux2_1 _24481_ (.A0(_09298_),
    .A1(\datamem.data_ram[52][24] ),
    .S(_10430_),
    .X(_10431_));
 sky130_fd_sc_hd__clkbuf_1 _24482_ (.A(_10431_),
    .X(_02340_));
 sky130_fd_sc_hd__mux2_1 _24483_ (.A0(_09306_),
    .A1(\datamem.data_ram[52][25] ),
    .S(_10430_),
    .X(_10432_));
 sky130_fd_sc_hd__clkbuf_1 _24484_ (.A(_10432_),
    .X(_02341_));
 sky130_fd_sc_hd__mux2_1 _24485_ (.A0(_09310_),
    .A1(\datamem.data_ram[52][26] ),
    .S(_10430_),
    .X(_10433_));
 sky130_fd_sc_hd__clkbuf_1 _24486_ (.A(_10433_),
    .X(_02342_));
 sky130_fd_sc_hd__mux2_1 _24487_ (.A0(_09314_),
    .A1(\datamem.data_ram[52][27] ),
    .S(_10430_),
    .X(_10434_));
 sky130_fd_sc_hd__clkbuf_1 _24488_ (.A(_10434_),
    .X(_02343_));
 sky130_fd_sc_hd__mux2_1 _24489_ (.A0(_09318_),
    .A1(\datamem.data_ram[52][28] ),
    .S(_10430_),
    .X(_10435_));
 sky130_fd_sc_hd__clkbuf_1 _24490_ (.A(_10435_),
    .X(_02344_));
 sky130_fd_sc_hd__mux2_1 _24491_ (.A0(_09322_),
    .A1(\datamem.data_ram[52][29] ),
    .S(_10430_),
    .X(_10436_));
 sky130_fd_sc_hd__clkbuf_1 _24492_ (.A(_10436_),
    .X(_02345_));
 sky130_fd_sc_hd__mux2_1 _24493_ (.A0(_09326_),
    .A1(\datamem.data_ram[52][30] ),
    .S(_10430_),
    .X(_10437_));
 sky130_fd_sc_hd__clkbuf_1 _24494_ (.A(_10437_),
    .X(_02346_));
 sky130_fd_sc_hd__mux2_1 _24495_ (.A0(_09330_),
    .A1(\datamem.data_ram[52][31] ),
    .S(_10430_),
    .X(_10438_));
 sky130_fd_sc_hd__clkbuf_1 _24496_ (.A(_10438_),
    .X(_02347_));
 sky130_fd_sc_hd__buf_2 _24497_ (.A(_09223_),
    .X(_10439_));
 sky130_fd_sc_hd__a21oi_4 _24498_ (.A1(_09351_),
    .A2(_10337_),
    .B1(_10366_),
    .Y(_10440_));
 sky130_fd_sc_hd__mux2_1 _24499_ (.A0(_10439_),
    .A1(\datamem.data_ram[52][16] ),
    .S(_10440_),
    .X(_10441_));
 sky130_fd_sc_hd__clkbuf_1 _24500_ (.A(_10441_),
    .X(_02348_));
 sky130_fd_sc_hd__buf_2 _24501_ (.A(_09235_),
    .X(_10442_));
 sky130_fd_sc_hd__mux2_1 _24502_ (.A0(_10442_),
    .A1(\datamem.data_ram[52][17] ),
    .S(_10440_),
    .X(_10443_));
 sky130_fd_sc_hd__clkbuf_1 _24503_ (.A(_10443_),
    .X(_02349_));
 sky130_fd_sc_hd__clkbuf_2 _24504_ (.A(_09239_),
    .X(_10444_));
 sky130_fd_sc_hd__mux2_1 _24505_ (.A0(_10444_),
    .A1(\datamem.data_ram[52][18] ),
    .S(_10440_),
    .X(_10445_));
 sky130_fd_sc_hd__clkbuf_1 _24506_ (.A(_10445_),
    .X(_02350_));
 sky130_fd_sc_hd__buf_2 _24507_ (.A(_09243_),
    .X(_10446_));
 sky130_fd_sc_hd__mux2_1 _24508_ (.A0(_10446_),
    .A1(\datamem.data_ram[52][19] ),
    .S(_10440_),
    .X(_10447_));
 sky130_fd_sc_hd__clkbuf_1 _24509_ (.A(_10447_),
    .X(_02351_));
 sky130_fd_sc_hd__clkbuf_2 _24510_ (.A(_09247_),
    .X(_10448_));
 sky130_fd_sc_hd__mux2_1 _24511_ (.A0(_10448_),
    .A1(\datamem.data_ram[52][20] ),
    .S(_10440_),
    .X(_10449_));
 sky130_fd_sc_hd__clkbuf_1 _24512_ (.A(_10449_),
    .X(_02352_));
 sky130_fd_sc_hd__clkbuf_2 _24513_ (.A(_09251_),
    .X(_10450_));
 sky130_fd_sc_hd__mux2_1 _24514_ (.A0(_10450_),
    .A1(\datamem.data_ram[52][21] ),
    .S(_10440_),
    .X(_10451_));
 sky130_fd_sc_hd__clkbuf_1 _24515_ (.A(_10451_),
    .X(_02353_));
 sky130_fd_sc_hd__clkbuf_2 _24516_ (.A(_09255_),
    .X(_10452_));
 sky130_fd_sc_hd__mux2_1 _24517_ (.A0(_10452_),
    .A1(\datamem.data_ram[52][22] ),
    .S(_10440_),
    .X(_10453_));
 sky130_fd_sc_hd__clkbuf_1 _24518_ (.A(_10453_),
    .X(_02354_));
 sky130_fd_sc_hd__buf_2 _24519_ (.A(_09259_),
    .X(_10454_));
 sky130_fd_sc_hd__mux2_1 _24520_ (.A0(_10454_),
    .A1(\datamem.data_ram[52][23] ),
    .S(_10440_),
    .X(_10455_));
 sky130_fd_sc_hd__clkbuf_1 _24521_ (.A(_10455_),
    .X(_02355_));
 sky130_fd_sc_hd__a21oi_4 _24522_ (.A1(_09351_),
    .A2(_10347_),
    .B1(_10366_),
    .Y(_10456_));
 sky130_fd_sc_hd__mux2_1 _24523_ (.A0(_10385_),
    .A1(\datamem.data_ram[52][8] ),
    .S(_10456_),
    .X(_10457_));
 sky130_fd_sc_hd__clkbuf_1 _24524_ (.A(_10457_),
    .X(_02356_));
 sky130_fd_sc_hd__mux2_1 _24525_ (.A0(_10388_),
    .A1(\datamem.data_ram[52][9] ),
    .S(_10456_),
    .X(_10458_));
 sky130_fd_sc_hd__clkbuf_1 _24526_ (.A(_10458_),
    .X(_02357_));
 sky130_fd_sc_hd__mux2_1 _24527_ (.A0(_10390_),
    .A1(\datamem.data_ram[52][10] ),
    .S(_10456_),
    .X(_10459_));
 sky130_fd_sc_hd__clkbuf_1 _24528_ (.A(_10459_),
    .X(_02358_));
 sky130_fd_sc_hd__mux2_1 _24529_ (.A0(_10392_),
    .A1(\datamem.data_ram[52][11] ),
    .S(_10456_),
    .X(_10460_));
 sky130_fd_sc_hd__clkbuf_1 _24530_ (.A(_10460_),
    .X(_02359_));
 sky130_fd_sc_hd__mux2_1 _24531_ (.A0(_10394_),
    .A1(\datamem.data_ram[52][12] ),
    .S(_10456_),
    .X(_10461_));
 sky130_fd_sc_hd__clkbuf_1 _24532_ (.A(_10461_),
    .X(_02360_));
 sky130_fd_sc_hd__mux2_1 _24533_ (.A0(_10396_),
    .A1(\datamem.data_ram[52][13] ),
    .S(_10456_),
    .X(_10462_));
 sky130_fd_sc_hd__clkbuf_1 _24534_ (.A(_10462_),
    .X(_02361_));
 sky130_fd_sc_hd__mux2_1 _24535_ (.A0(_10398_),
    .A1(\datamem.data_ram[52][14] ),
    .S(_10456_),
    .X(_10463_));
 sky130_fd_sc_hd__clkbuf_1 _24536_ (.A(_10463_),
    .X(_02362_));
 sky130_fd_sc_hd__mux2_1 _24537_ (.A0(_10400_),
    .A1(\datamem.data_ram[52][15] ),
    .S(_10456_),
    .X(_10464_));
 sky130_fd_sc_hd__clkbuf_1 _24538_ (.A(_10464_),
    .X(_02363_));
 sky130_fd_sc_hd__buf_2 _24539_ (.A(_09297_),
    .X(_10465_));
 sky130_fd_sc_hd__a21oi_2 _24540_ (.A1(_10142_),
    .A2(_10327_),
    .B1(_10366_),
    .Y(_10466_));
 sky130_fd_sc_hd__mux2_1 _24541_ (.A0(_10465_),
    .A1(\datamem.data_ram[51][24] ),
    .S(net60),
    .X(_10467_));
 sky130_fd_sc_hd__clkbuf_1 _24542_ (.A(_10467_),
    .X(_02364_));
 sky130_fd_sc_hd__clkbuf_2 _24543_ (.A(_09305_),
    .X(_10468_));
 sky130_fd_sc_hd__mux2_1 _24544_ (.A0(_10468_),
    .A1(\datamem.data_ram[51][25] ),
    .S(net60),
    .X(_10469_));
 sky130_fd_sc_hd__clkbuf_1 _24545_ (.A(_10469_),
    .X(_02365_));
 sky130_fd_sc_hd__buf_2 _24546_ (.A(_09309_),
    .X(_10470_));
 sky130_fd_sc_hd__mux2_1 _24547_ (.A0(_10470_),
    .A1(\datamem.data_ram[51][26] ),
    .S(_10466_),
    .X(_10471_));
 sky130_fd_sc_hd__clkbuf_1 _24548_ (.A(_10471_),
    .X(_02366_));
 sky130_fd_sc_hd__clkbuf_2 _24549_ (.A(_09313_),
    .X(_10472_));
 sky130_fd_sc_hd__mux2_1 _24550_ (.A0(_10472_),
    .A1(\datamem.data_ram[51][27] ),
    .S(net60),
    .X(_10473_));
 sky130_fd_sc_hd__clkbuf_1 _24551_ (.A(_10473_),
    .X(_02367_));
 sky130_fd_sc_hd__clkbuf_2 _24552_ (.A(_09317_),
    .X(_10474_));
 sky130_fd_sc_hd__mux2_1 _24553_ (.A0(_10474_),
    .A1(\datamem.data_ram[51][28] ),
    .S(net60),
    .X(_10475_));
 sky130_fd_sc_hd__clkbuf_1 _24554_ (.A(_10475_),
    .X(_02368_));
 sky130_fd_sc_hd__clkbuf_2 _24555_ (.A(_09321_),
    .X(_10476_));
 sky130_fd_sc_hd__mux2_1 _24556_ (.A0(_10476_),
    .A1(\datamem.data_ram[51][29] ),
    .S(net60),
    .X(_10477_));
 sky130_fd_sc_hd__clkbuf_1 _24557_ (.A(_10477_),
    .X(_02369_));
 sky130_fd_sc_hd__clkbuf_2 _24558_ (.A(_09325_),
    .X(_10478_));
 sky130_fd_sc_hd__mux2_1 _24559_ (.A0(_10478_),
    .A1(\datamem.data_ram[51][30] ),
    .S(net60),
    .X(_10479_));
 sky130_fd_sc_hd__clkbuf_1 _24560_ (.A(_10479_),
    .X(_02370_));
 sky130_fd_sc_hd__clkbuf_2 _24561_ (.A(_09329_),
    .X(_10480_));
 sky130_fd_sc_hd__mux2_1 _24562_ (.A0(_10480_),
    .A1(\datamem.data_ram[51][31] ),
    .S(_10466_),
    .X(_10481_));
 sky130_fd_sc_hd__clkbuf_1 _24563_ (.A(_10481_),
    .X(_02371_));
 sky130_fd_sc_hd__a21oi_4 _24564_ (.A1(_10142_),
    .A2(_10337_),
    .B1(_10366_),
    .Y(_10482_));
 sky130_fd_sc_hd__mux2_1 _24565_ (.A0(_10439_),
    .A1(\datamem.data_ram[51][16] ),
    .S(_10482_),
    .X(_10483_));
 sky130_fd_sc_hd__clkbuf_1 _24566_ (.A(_10483_),
    .X(_02372_));
 sky130_fd_sc_hd__mux2_1 _24567_ (.A0(_10442_),
    .A1(\datamem.data_ram[51][17] ),
    .S(_10482_),
    .X(_10484_));
 sky130_fd_sc_hd__clkbuf_1 _24568_ (.A(_10484_),
    .X(_02373_));
 sky130_fd_sc_hd__mux2_1 _24569_ (.A0(_10444_),
    .A1(\datamem.data_ram[51][18] ),
    .S(_10482_),
    .X(_10485_));
 sky130_fd_sc_hd__clkbuf_1 _24570_ (.A(_10485_),
    .X(_02374_));
 sky130_fd_sc_hd__mux2_1 _24571_ (.A0(_10446_),
    .A1(\datamem.data_ram[51][19] ),
    .S(_10482_),
    .X(_10486_));
 sky130_fd_sc_hd__clkbuf_1 _24572_ (.A(_10486_),
    .X(_02375_));
 sky130_fd_sc_hd__mux2_1 _24573_ (.A0(_10448_),
    .A1(\datamem.data_ram[51][20] ),
    .S(_10482_),
    .X(_10487_));
 sky130_fd_sc_hd__clkbuf_1 _24574_ (.A(_10487_),
    .X(_02376_));
 sky130_fd_sc_hd__mux2_1 _24575_ (.A0(_10450_),
    .A1(\datamem.data_ram[51][21] ),
    .S(_10482_),
    .X(_10488_));
 sky130_fd_sc_hd__clkbuf_1 _24576_ (.A(_10488_),
    .X(_02377_));
 sky130_fd_sc_hd__mux2_1 _24577_ (.A0(_10452_),
    .A1(\datamem.data_ram[51][22] ),
    .S(_10482_),
    .X(_10489_));
 sky130_fd_sc_hd__clkbuf_1 _24578_ (.A(_10489_),
    .X(_02378_));
 sky130_fd_sc_hd__mux2_1 _24579_ (.A0(_10454_),
    .A1(\datamem.data_ram[51][23] ),
    .S(_10482_),
    .X(_10490_));
 sky130_fd_sc_hd__clkbuf_1 _24580_ (.A(_10490_),
    .X(_02379_));
 sky130_fd_sc_hd__a21oi_4 _24581_ (.A1(_10142_),
    .A2(_10347_),
    .B1(_10366_),
    .Y(_10491_));
 sky130_fd_sc_hd__mux2_1 _24582_ (.A0(_10385_),
    .A1(\datamem.data_ram[51][8] ),
    .S(_10491_),
    .X(_10492_));
 sky130_fd_sc_hd__clkbuf_1 _24583_ (.A(_10492_),
    .X(_02380_));
 sky130_fd_sc_hd__mux2_1 _24584_ (.A0(_10388_),
    .A1(\datamem.data_ram[51][9] ),
    .S(_10491_),
    .X(_10493_));
 sky130_fd_sc_hd__clkbuf_1 _24585_ (.A(_10493_),
    .X(_02381_));
 sky130_fd_sc_hd__mux2_1 _24586_ (.A0(_10390_),
    .A1(\datamem.data_ram[51][10] ),
    .S(_10491_),
    .X(_10494_));
 sky130_fd_sc_hd__clkbuf_1 _24587_ (.A(_10494_),
    .X(_02382_));
 sky130_fd_sc_hd__mux2_1 _24588_ (.A0(_10392_),
    .A1(\datamem.data_ram[51][11] ),
    .S(_10491_),
    .X(_10495_));
 sky130_fd_sc_hd__clkbuf_1 _24589_ (.A(_10495_),
    .X(_02383_));
 sky130_fd_sc_hd__mux2_1 _24590_ (.A0(_10394_),
    .A1(\datamem.data_ram[51][12] ),
    .S(_10491_),
    .X(_10496_));
 sky130_fd_sc_hd__clkbuf_1 _24591_ (.A(_10496_),
    .X(_02384_));
 sky130_fd_sc_hd__mux2_1 _24592_ (.A0(_10396_),
    .A1(\datamem.data_ram[51][13] ),
    .S(_10491_),
    .X(_10497_));
 sky130_fd_sc_hd__clkbuf_1 _24593_ (.A(_10497_),
    .X(_02385_));
 sky130_fd_sc_hd__mux2_1 _24594_ (.A0(_10398_),
    .A1(\datamem.data_ram[51][14] ),
    .S(_10491_),
    .X(_10498_));
 sky130_fd_sc_hd__clkbuf_1 _24595_ (.A(_10498_),
    .X(_02386_));
 sky130_fd_sc_hd__mux2_1 _24596_ (.A0(_10400_),
    .A1(\datamem.data_ram[51][15] ),
    .S(_10491_),
    .X(_10499_));
 sky130_fd_sc_hd__clkbuf_1 _24597_ (.A(_10499_),
    .X(_02387_));
 sky130_fd_sc_hd__buf_4 _24598_ (.A(_06591_),
    .X(_10500_));
 sky130_fd_sc_hd__buf_8 _24599_ (.A(_10500_),
    .X(_10501_));
 sky130_fd_sc_hd__a21oi_4 _24600_ (.A1(_10209_),
    .A2(_10327_),
    .B1(_10501_),
    .Y(_10502_));
 sky130_fd_sc_hd__mux2_1 _24601_ (.A0(_10465_),
    .A1(\datamem.data_ram[50][24] ),
    .S(_10502_),
    .X(_10503_));
 sky130_fd_sc_hd__clkbuf_1 _24602_ (.A(_10503_),
    .X(_02388_));
 sky130_fd_sc_hd__mux2_1 _24603_ (.A0(_10468_),
    .A1(\datamem.data_ram[50][25] ),
    .S(_10502_),
    .X(_10504_));
 sky130_fd_sc_hd__clkbuf_1 _24604_ (.A(_10504_),
    .X(_02389_));
 sky130_fd_sc_hd__mux2_1 _24605_ (.A0(_10470_),
    .A1(\datamem.data_ram[50][26] ),
    .S(_10502_),
    .X(_10505_));
 sky130_fd_sc_hd__clkbuf_1 _24606_ (.A(_10505_),
    .X(_02390_));
 sky130_fd_sc_hd__mux2_1 _24607_ (.A0(_10472_),
    .A1(\datamem.data_ram[50][27] ),
    .S(_10502_),
    .X(_10506_));
 sky130_fd_sc_hd__clkbuf_1 _24608_ (.A(_10506_),
    .X(_02391_));
 sky130_fd_sc_hd__mux2_1 _24609_ (.A0(_10474_),
    .A1(\datamem.data_ram[50][28] ),
    .S(_10502_),
    .X(_10507_));
 sky130_fd_sc_hd__clkbuf_1 _24610_ (.A(_10507_),
    .X(_02392_));
 sky130_fd_sc_hd__mux2_1 _24611_ (.A0(_10476_),
    .A1(\datamem.data_ram[50][29] ),
    .S(_10502_),
    .X(_10508_));
 sky130_fd_sc_hd__clkbuf_1 _24612_ (.A(_10508_),
    .X(_02393_));
 sky130_fd_sc_hd__mux2_1 _24613_ (.A0(_10478_),
    .A1(\datamem.data_ram[50][30] ),
    .S(_10502_),
    .X(_10509_));
 sky130_fd_sc_hd__clkbuf_1 _24614_ (.A(_10509_),
    .X(_02394_));
 sky130_fd_sc_hd__mux2_1 _24615_ (.A0(_10480_),
    .A1(\datamem.data_ram[50][31] ),
    .S(_10502_),
    .X(_10510_));
 sky130_fd_sc_hd__clkbuf_1 _24616_ (.A(_10510_),
    .X(_02395_));
 sky130_fd_sc_hd__a21oi_4 _24617_ (.A1(_10209_),
    .A2(_10337_),
    .B1(_10501_),
    .Y(_10511_));
 sky130_fd_sc_hd__mux2_1 _24618_ (.A0(_10439_),
    .A1(\datamem.data_ram[50][16] ),
    .S(_10511_),
    .X(_10512_));
 sky130_fd_sc_hd__clkbuf_1 _24619_ (.A(_10512_),
    .X(_02396_));
 sky130_fd_sc_hd__mux2_1 _24620_ (.A0(_10442_),
    .A1(\datamem.data_ram[50][17] ),
    .S(_10511_),
    .X(_10513_));
 sky130_fd_sc_hd__clkbuf_1 _24621_ (.A(_10513_),
    .X(_02397_));
 sky130_fd_sc_hd__mux2_1 _24622_ (.A0(_10444_),
    .A1(\datamem.data_ram[50][18] ),
    .S(_10511_),
    .X(_10514_));
 sky130_fd_sc_hd__clkbuf_1 _24623_ (.A(_10514_),
    .X(_02398_));
 sky130_fd_sc_hd__mux2_1 _24624_ (.A0(_10446_),
    .A1(\datamem.data_ram[50][19] ),
    .S(_10511_),
    .X(_10515_));
 sky130_fd_sc_hd__clkbuf_1 _24625_ (.A(_10515_),
    .X(_02399_));
 sky130_fd_sc_hd__mux2_1 _24626_ (.A0(_10448_),
    .A1(\datamem.data_ram[50][20] ),
    .S(_10511_),
    .X(_10516_));
 sky130_fd_sc_hd__clkbuf_1 _24627_ (.A(_10516_),
    .X(_02400_));
 sky130_fd_sc_hd__mux2_1 _24628_ (.A0(_10450_),
    .A1(\datamem.data_ram[50][21] ),
    .S(_10511_),
    .X(_10517_));
 sky130_fd_sc_hd__clkbuf_1 _24629_ (.A(_10517_),
    .X(_02401_));
 sky130_fd_sc_hd__mux2_1 _24630_ (.A0(_10452_),
    .A1(\datamem.data_ram[50][22] ),
    .S(_10511_),
    .X(_10518_));
 sky130_fd_sc_hd__clkbuf_1 _24631_ (.A(_10518_),
    .X(_02402_));
 sky130_fd_sc_hd__mux2_1 _24632_ (.A0(_10454_),
    .A1(\datamem.data_ram[50][23] ),
    .S(_10511_),
    .X(_10519_));
 sky130_fd_sc_hd__clkbuf_1 _24633_ (.A(_10519_),
    .X(_02403_));
 sky130_fd_sc_hd__buf_8 _24634_ (.A(_07136_),
    .X(_10520_));
 sky130_fd_sc_hd__a21oi_4 _24635_ (.A1(_10520_),
    .A2(_10347_),
    .B1(_10501_),
    .Y(_10521_));
 sky130_fd_sc_hd__mux2_1 _24636_ (.A0(_10385_),
    .A1(\datamem.data_ram[50][8] ),
    .S(_10521_),
    .X(_10522_));
 sky130_fd_sc_hd__clkbuf_1 _24637_ (.A(_10522_),
    .X(_02404_));
 sky130_fd_sc_hd__mux2_1 _24638_ (.A0(_10388_),
    .A1(\datamem.data_ram[50][9] ),
    .S(_10521_),
    .X(_10523_));
 sky130_fd_sc_hd__clkbuf_1 _24639_ (.A(_10523_),
    .X(_02405_));
 sky130_fd_sc_hd__mux2_1 _24640_ (.A0(_10390_),
    .A1(\datamem.data_ram[50][10] ),
    .S(_10521_),
    .X(_10524_));
 sky130_fd_sc_hd__clkbuf_1 _24641_ (.A(_10524_),
    .X(_02406_));
 sky130_fd_sc_hd__mux2_1 _24642_ (.A0(_10392_),
    .A1(\datamem.data_ram[50][11] ),
    .S(_10521_),
    .X(_10525_));
 sky130_fd_sc_hd__clkbuf_1 _24643_ (.A(_10525_),
    .X(_02407_));
 sky130_fd_sc_hd__mux2_1 _24644_ (.A0(_10394_),
    .A1(\datamem.data_ram[50][12] ),
    .S(_10521_),
    .X(_10526_));
 sky130_fd_sc_hd__clkbuf_1 _24645_ (.A(_10526_),
    .X(_02408_));
 sky130_fd_sc_hd__mux2_1 _24646_ (.A0(_10396_),
    .A1(\datamem.data_ram[50][13] ),
    .S(_10521_),
    .X(_10527_));
 sky130_fd_sc_hd__clkbuf_1 _24647_ (.A(_10527_),
    .X(_02409_));
 sky130_fd_sc_hd__mux2_1 _24648_ (.A0(_10398_),
    .A1(\datamem.data_ram[50][14] ),
    .S(_10521_),
    .X(_10528_));
 sky130_fd_sc_hd__clkbuf_1 _24649_ (.A(_10528_),
    .X(_02410_));
 sky130_fd_sc_hd__mux2_1 _24650_ (.A0(_10400_),
    .A1(\datamem.data_ram[50][15] ),
    .S(_10521_),
    .X(_10529_));
 sky130_fd_sc_hd__clkbuf_1 _24651_ (.A(_10529_),
    .X(_02411_));
 sky130_fd_sc_hd__or3_1 _24652_ (.A(_07182_),
    .B(_10042_),
    .C(_10044_),
    .X(_10530_));
 sky130_fd_sc_hd__buf_2 _24653_ (.A(_10530_),
    .X(_10531_));
 sky130_fd_sc_hd__and3_2 _24654_ (.A(_09351_),
    .B(_10049_),
    .C(_10052_),
    .X(_10532_));
 sky130_fd_sc_hd__and2_1 _24655_ (.A(_10405_),
    .B(_10532_),
    .X(_10533_));
 sky130_fd_sc_hd__a31o_1 _24656_ (.A1(_10412_),
    .A2(\datamem.data_ram[4][0] ),
    .A3(_10531_),
    .B1(_10533_),
    .X(_02412_));
 sky130_fd_sc_hd__and2_1 _24657_ (.A(_10408_),
    .B(_10532_),
    .X(_10534_));
 sky130_fd_sc_hd__a31o_1 _24658_ (.A1(_10412_),
    .A2(\datamem.data_ram[4][1] ),
    .A3(_10531_),
    .B1(_10534_),
    .X(_02413_));
 sky130_fd_sc_hd__and2_1 _24659_ (.A(_10410_),
    .B(_10532_),
    .X(_10535_));
 sky130_fd_sc_hd__a31o_1 _24660_ (.A1(_10412_),
    .A2(\datamem.data_ram[4][2] ),
    .A3(_10531_),
    .B1(_10535_),
    .X(_02414_));
 sky130_fd_sc_hd__and2_1 _24661_ (.A(_10413_),
    .B(_10532_),
    .X(_10536_));
 sky130_fd_sc_hd__a31o_1 _24662_ (.A1(_10412_),
    .A2(\datamem.data_ram[4][3] ),
    .A3(_10531_),
    .B1(_10536_),
    .X(_02415_));
 sky130_fd_sc_hd__and2_1 _24663_ (.A(_10067_),
    .B(_10532_),
    .X(_10537_));
 sky130_fd_sc_hd__a31o_1 _24664_ (.A1(_10412_),
    .A2(\datamem.data_ram[4][4] ),
    .A3(_10531_),
    .B1(_10537_),
    .X(_02416_));
 sky130_fd_sc_hd__buf_2 _24665_ (.A(_10055_),
    .X(_10538_));
 sky130_fd_sc_hd__and2_1 _24666_ (.A(_10416_),
    .B(_10532_),
    .X(_10539_));
 sky130_fd_sc_hd__a31o_1 _24667_ (.A1(_10538_),
    .A2(\datamem.data_ram[4][5] ),
    .A3(_10531_),
    .B1(_10539_),
    .X(_02417_));
 sky130_fd_sc_hd__and2_1 _24668_ (.A(_10418_),
    .B(_10532_),
    .X(_10540_));
 sky130_fd_sc_hd__a31o_1 _24669_ (.A1(_10538_),
    .A2(\datamem.data_ram[4][6] ),
    .A3(_10531_),
    .B1(_10540_),
    .X(_02418_));
 sky130_fd_sc_hd__and2_1 _24670_ (.A(_10076_),
    .B(_10532_),
    .X(_10541_));
 sky130_fd_sc_hd__a31o_1 _24671_ (.A1(_10538_),
    .A2(\datamem.data_ram[4][7] ),
    .A3(_10531_),
    .B1(_10541_),
    .X(_02419_));
 sky130_fd_sc_hd__buf_8 _24672_ (.A(_07123_),
    .X(_10542_));
 sky130_fd_sc_hd__a21oi_4 _24673_ (.A1(_10542_),
    .A2(_10092_),
    .B1(_10501_),
    .Y(_10543_));
 sky130_fd_sc_hd__mux2_1 _24674_ (.A0(_10385_),
    .A1(\datamem.data_ram[4][8] ),
    .S(_10543_),
    .X(_10544_));
 sky130_fd_sc_hd__clkbuf_1 _24675_ (.A(_10544_),
    .X(_02420_));
 sky130_fd_sc_hd__mux2_1 _24676_ (.A0(_10388_),
    .A1(\datamem.data_ram[4][9] ),
    .S(_10543_),
    .X(_10545_));
 sky130_fd_sc_hd__clkbuf_1 _24677_ (.A(_10545_),
    .X(_02421_));
 sky130_fd_sc_hd__mux2_1 _24678_ (.A0(_10390_),
    .A1(\datamem.data_ram[4][10] ),
    .S(_10543_),
    .X(_10546_));
 sky130_fd_sc_hd__clkbuf_1 _24679_ (.A(_10546_),
    .X(_02422_));
 sky130_fd_sc_hd__mux2_1 _24680_ (.A0(_10392_),
    .A1(\datamem.data_ram[4][11] ),
    .S(_10543_),
    .X(_10547_));
 sky130_fd_sc_hd__clkbuf_1 _24681_ (.A(_10547_),
    .X(_02423_));
 sky130_fd_sc_hd__mux2_1 _24682_ (.A0(_10394_),
    .A1(\datamem.data_ram[4][12] ),
    .S(_10543_),
    .X(_10548_));
 sky130_fd_sc_hd__clkbuf_1 _24683_ (.A(_10548_),
    .X(_02424_));
 sky130_fd_sc_hd__mux2_1 _24684_ (.A0(_10396_),
    .A1(\datamem.data_ram[4][13] ),
    .S(_10543_),
    .X(_10549_));
 sky130_fd_sc_hd__clkbuf_1 _24685_ (.A(_10549_),
    .X(_02425_));
 sky130_fd_sc_hd__mux2_1 _24686_ (.A0(_10398_),
    .A1(\datamem.data_ram[4][14] ),
    .S(_10543_),
    .X(_10550_));
 sky130_fd_sc_hd__clkbuf_1 _24687_ (.A(_10550_),
    .X(_02426_));
 sky130_fd_sc_hd__mux2_1 _24688_ (.A0(_10400_),
    .A1(\datamem.data_ram[4][15] ),
    .S(_10543_),
    .X(_10551_));
 sky130_fd_sc_hd__clkbuf_1 _24689_ (.A(_10551_),
    .X(_02427_));
 sky130_fd_sc_hd__a21oi_4 _24690_ (.A1(_10542_),
    .A2(_10114_),
    .B1(_10501_),
    .Y(_10552_));
 sky130_fd_sc_hd__mux2_1 _24691_ (.A0(_10439_),
    .A1(\datamem.data_ram[4][16] ),
    .S(_10552_),
    .X(_10553_));
 sky130_fd_sc_hd__clkbuf_1 _24692_ (.A(_10553_),
    .X(_02428_));
 sky130_fd_sc_hd__mux2_1 _24693_ (.A0(_10442_),
    .A1(\datamem.data_ram[4][17] ),
    .S(_10552_),
    .X(_10554_));
 sky130_fd_sc_hd__clkbuf_1 _24694_ (.A(_10554_),
    .X(_02429_));
 sky130_fd_sc_hd__mux2_1 _24695_ (.A0(_10444_),
    .A1(\datamem.data_ram[4][18] ),
    .S(_10552_),
    .X(_10555_));
 sky130_fd_sc_hd__clkbuf_1 _24696_ (.A(_10555_),
    .X(_02430_));
 sky130_fd_sc_hd__mux2_1 _24697_ (.A0(_10446_),
    .A1(\datamem.data_ram[4][19] ),
    .S(_10552_),
    .X(_10556_));
 sky130_fd_sc_hd__clkbuf_1 _24698_ (.A(_10556_),
    .X(_02431_));
 sky130_fd_sc_hd__mux2_1 _24699_ (.A0(_10448_),
    .A1(\datamem.data_ram[4][20] ),
    .S(_10552_),
    .X(_10557_));
 sky130_fd_sc_hd__clkbuf_1 _24700_ (.A(_10557_),
    .X(_02432_));
 sky130_fd_sc_hd__mux2_1 _24701_ (.A0(_10450_),
    .A1(\datamem.data_ram[4][21] ),
    .S(_10552_),
    .X(_10558_));
 sky130_fd_sc_hd__clkbuf_1 _24702_ (.A(_10558_),
    .X(_02433_));
 sky130_fd_sc_hd__mux2_1 _24703_ (.A0(_10452_),
    .A1(\datamem.data_ram[4][22] ),
    .S(_10552_),
    .X(_10559_));
 sky130_fd_sc_hd__clkbuf_1 _24704_ (.A(_10559_),
    .X(_02434_));
 sky130_fd_sc_hd__mux2_1 _24705_ (.A0(_10454_),
    .A1(\datamem.data_ram[4][23] ),
    .S(_10552_),
    .X(_10560_));
 sky130_fd_sc_hd__clkbuf_1 _24706_ (.A(_10560_),
    .X(_02435_));
 sky130_fd_sc_hd__a21oi_2 _24707_ (.A1(_10268_),
    .A2(_10327_),
    .B1(_10501_),
    .Y(_10561_));
 sky130_fd_sc_hd__mux2_1 _24708_ (.A0(_10465_),
    .A1(\datamem.data_ram[49][24] ),
    .S(net59),
    .X(_10562_));
 sky130_fd_sc_hd__clkbuf_1 _24709_ (.A(_10562_),
    .X(_02436_));
 sky130_fd_sc_hd__mux2_1 _24710_ (.A0(_10468_),
    .A1(\datamem.data_ram[49][25] ),
    .S(net59),
    .X(_10563_));
 sky130_fd_sc_hd__clkbuf_1 _24711_ (.A(_10563_),
    .X(_02437_));
 sky130_fd_sc_hd__mux2_1 _24712_ (.A0(_10470_),
    .A1(\datamem.data_ram[49][26] ),
    .S(_10561_),
    .X(_10564_));
 sky130_fd_sc_hd__clkbuf_1 _24713_ (.A(_10564_),
    .X(_02438_));
 sky130_fd_sc_hd__mux2_1 _24714_ (.A0(_10472_),
    .A1(\datamem.data_ram[49][27] ),
    .S(net59),
    .X(_10565_));
 sky130_fd_sc_hd__clkbuf_1 _24715_ (.A(_10565_),
    .X(_02439_));
 sky130_fd_sc_hd__mux2_1 _24716_ (.A0(_10474_),
    .A1(\datamem.data_ram[49][28] ),
    .S(net59),
    .X(_10566_));
 sky130_fd_sc_hd__clkbuf_1 _24717_ (.A(_10566_),
    .X(_02440_));
 sky130_fd_sc_hd__mux2_1 _24718_ (.A0(_10476_),
    .A1(\datamem.data_ram[49][29] ),
    .S(net59),
    .X(_10567_));
 sky130_fd_sc_hd__clkbuf_1 _24719_ (.A(_10567_),
    .X(_02441_));
 sky130_fd_sc_hd__mux2_1 _24720_ (.A0(_10478_),
    .A1(\datamem.data_ram[49][30] ),
    .S(net59),
    .X(_10568_));
 sky130_fd_sc_hd__clkbuf_1 _24721_ (.A(_10568_),
    .X(_02442_));
 sky130_fd_sc_hd__mux2_1 _24722_ (.A0(_10480_),
    .A1(\datamem.data_ram[49][31] ),
    .S(_10561_),
    .X(_10569_));
 sky130_fd_sc_hd__clkbuf_1 _24723_ (.A(_10569_),
    .X(_02443_));
 sky130_fd_sc_hd__buf_8 _24724_ (.A(_06997_),
    .X(_10570_));
 sky130_fd_sc_hd__a21oi_4 _24725_ (.A1(_10570_),
    .A2(_10337_),
    .B1(_10501_),
    .Y(_10571_));
 sky130_fd_sc_hd__mux2_1 _24726_ (.A0(_10439_),
    .A1(\datamem.data_ram[49][16] ),
    .S(_10571_),
    .X(_10572_));
 sky130_fd_sc_hd__clkbuf_1 _24727_ (.A(_10572_),
    .X(_02444_));
 sky130_fd_sc_hd__mux2_1 _24728_ (.A0(_10442_),
    .A1(\datamem.data_ram[49][17] ),
    .S(_10571_),
    .X(_10573_));
 sky130_fd_sc_hd__clkbuf_1 _24729_ (.A(_10573_),
    .X(_02445_));
 sky130_fd_sc_hd__mux2_1 _24730_ (.A0(_10444_),
    .A1(\datamem.data_ram[49][18] ),
    .S(_10571_),
    .X(_10574_));
 sky130_fd_sc_hd__clkbuf_1 _24731_ (.A(_10574_),
    .X(_02446_));
 sky130_fd_sc_hd__mux2_1 _24732_ (.A0(_10446_),
    .A1(\datamem.data_ram[49][19] ),
    .S(_10571_),
    .X(_10575_));
 sky130_fd_sc_hd__clkbuf_1 _24733_ (.A(_10575_),
    .X(_02447_));
 sky130_fd_sc_hd__mux2_1 _24734_ (.A0(_10448_),
    .A1(\datamem.data_ram[49][20] ),
    .S(_10571_),
    .X(_10576_));
 sky130_fd_sc_hd__clkbuf_1 _24735_ (.A(_10576_),
    .X(_02448_));
 sky130_fd_sc_hd__mux2_1 _24736_ (.A0(_10450_),
    .A1(\datamem.data_ram[49][21] ),
    .S(_10571_),
    .X(_10577_));
 sky130_fd_sc_hd__clkbuf_1 _24737_ (.A(_10577_),
    .X(_02449_));
 sky130_fd_sc_hd__mux2_1 _24738_ (.A0(_10452_),
    .A1(\datamem.data_ram[49][22] ),
    .S(_10571_),
    .X(_10578_));
 sky130_fd_sc_hd__clkbuf_1 _24739_ (.A(_10578_),
    .X(_02450_));
 sky130_fd_sc_hd__mux2_1 _24740_ (.A0(_10454_),
    .A1(\datamem.data_ram[49][23] ),
    .S(_10571_),
    .X(_10579_));
 sky130_fd_sc_hd__clkbuf_1 _24741_ (.A(_10579_),
    .X(_02451_));
 sky130_fd_sc_hd__a21oi_4 _24742_ (.A1(_10570_),
    .A2(_10347_),
    .B1(_10501_),
    .Y(_10580_));
 sky130_fd_sc_hd__mux2_1 _24743_ (.A0(_10385_),
    .A1(\datamem.data_ram[49][8] ),
    .S(_10580_),
    .X(_10581_));
 sky130_fd_sc_hd__clkbuf_1 _24744_ (.A(_10581_),
    .X(_02452_));
 sky130_fd_sc_hd__mux2_1 _24745_ (.A0(_10388_),
    .A1(\datamem.data_ram[49][9] ),
    .S(_10580_),
    .X(_10582_));
 sky130_fd_sc_hd__clkbuf_1 _24746_ (.A(_10582_),
    .X(_02453_));
 sky130_fd_sc_hd__mux2_1 _24747_ (.A0(_10390_),
    .A1(\datamem.data_ram[49][10] ),
    .S(_10580_),
    .X(_10583_));
 sky130_fd_sc_hd__clkbuf_1 _24748_ (.A(_10583_),
    .X(_02454_));
 sky130_fd_sc_hd__mux2_1 _24749_ (.A0(_10392_),
    .A1(\datamem.data_ram[49][11] ),
    .S(_10580_),
    .X(_10584_));
 sky130_fd_sc_hd__clkbuf_1 _24750_ (.A(_10584_),
    .X(_02455_));
 sky130_fd_sc_hd__mux2_1 _24751_ (.A0(_10394_),
    .A1(\datamem.data_ram[49][12] ),
    .S(_10580_),
    .X(_10585_));
 sky130_fd_sc_hd__clkbuf_1 _24752_ (.A(_10585_),
    .X(_02456_));
 sky130_fd_sc_hd__mux2_1 _24753_ (.A0(_10396_),
    .A1(\datamem.data_ram[49][13] ),
    .S(_10580_),
    .X(_10586_));
 sky130_fd_sc_hd__clkbuf_1 _24754_ (.A(_10586_),
    .X(_02457_));
 sky130_fd_sc_hd__mux2_1 _24755_ (.A0(_10398_),
    .A1(\datamem.data_ram[49][14] ),
    .S(_10580_),
    .X(_10587_));
 sky130_fd_sc_hd__clkbuf_1 _24756_ (.A(_10587_),
    .X(_02458_));
 sky130_fd_sc_hd__mux2_1 _24757_ (.A0(_10400_),
    .A1(\datamem.data_ram[49][15] ),
    .S(_10580_),
    .X(_10588_));
 sky130_fd_sc_hd__clkbuf_1 _24758_ (.A(_10588_),
    .X(_02459_));
 sky130_fd_sc_hd__a21oi_4 _24759_ (.A1(_10297_),
    .A2(_10327_),
    .B1(_10501_),
    .Y(_10589_));
 sky130_fd_sc_hd__mux2_1 _24760_ (.A0(_10465_),
    .A1(\datamem.data_ram[48][24] ),
    .S(_10589_),
    .X(_10590_));
 sky130_fd_sc_hd__clkbuf_1 _24761_ (.A(_10590_),
    .X(_02460_));
 sky130_fd_sc_hd__mux2_1 _24762_ (.A0(_10468_),
    .A1(\datamem.data_ram[48][25] ),
    .S(_10589_),
    .X(_10591_));
 sky130_fd_sc_hd__clkbuf_1 _24763_ (.A(_10591_),
    .X(_02461_));
 sky130_fd_sc_hd__mux2_1 _24764_ (.A0(_10470_),
    .A1(\datamem.data_ram[48][26] ),
    .S(_10589_),
    .X(_10592_));
 sky130_fd_sc_hd__clkbuf_1 _24765_ (.A(_10592_),
    .X(_02462_));
 sky130_fd_sc_hd__mux2_1 _24766_ (.A0(_10472_),
    .A1(\datamem.data_ram[48][27] ),
    .S(_10589_),
    .X(_10593_));
 sky130_fd_sc_hd__clkbuf_1 _24767_ (.A(_10593_),
    .X(_02463_));
 sky130_fd_sc_hd__mux2_1 _24768_ (.A0(_10474_),
    .A1(\datamem.data_ram[48][28] ),
    .S(_10589_),
    .X(_10594_));
 sky130_fd_sc_hd__clkbuf_1 _24769_ (.A(_10594_),
    .X(_02464_));
 sky130_fd_sc_hd__mux2_1 _24770_ (.A0(_10476_),
    .A1(\datamem.data_ram[48][29] ),
    .S(_10589_),
    .X(_10595_));
 sky130_fd_sc_hd__clkbuf_1 _24771_ (.A(_10595_),
    .X(_02465_));
 sky130_fd_sc_hd__mux2_1 _24772_ (.A0(_10478_),
    .A1(\datamem.data_ram[48][30] ),
    .S(_10589_),
    .X(_10596_));
 sky130_fd_sc_hd__clkbuf_1 _24773_ (.A(_10596_),
    .X(_02466_));
 sky130_fd_sc_hd__mux2_1 _24774_ (.A0(_10480_),
    .A1(\datamem.data_ram[48][31] ),
    .S(_10589_),
    .X(_10597_));
 sky130_fd_sc_hd__clkbuf_1 _24775_ (.A(_10597_),
    .X(_02467_));
 sky130_fd_sc_hd__buf_8 _24776_ (.A(_07125_),
    .X(_10598_));
 sky130_fd_sc_hd__nand2_2 _24777_ (.A(_08124_),
    .B(_07858_),
    .Y(_10599_));
 sky130_fd_sc_hd__buf_8 _24778_ (.A(_10599_),
    .X(_10600_));
 sky130_fd_sc_hd__nor2_2 _24779_ (.A(net108),
    .B(_10600_),
    .Y(_10601_));
 sky130_fd_sc_hd__a21oi_1 _24780_ (.A1(_10598_),
    .A2(_10601_),
    .B1(_10501_),
    .Y(_10602_));
 sky130_fd_sc_hd__mux2_1 _24781_ (.A0(_10465_),
    .A1(\datamem.data_ram[47][24] ),
    .S(net94),
    .X(_10603_));
 sky130_fd_sc_hd__clkbuf_1 _24782_ (.A(_10603_),
    .X(_02468_));
 sky130_fd_sc_hd__mux2_1 _24783_ (.A0(_10468_),
    .A1(\datamem.data_ram[47][25] ),
    .S(net94),
    .X(_10604_));
 sky130_fd_sc_hd__clkbuf_1 _24784_ (.A(_10604_),
    .X(_02469_));
 sky130_fd_sc_hd__mux2_1 _24785_ (.A0(_10470_),
    .A1(\datamem.data_ram[47][26] ),
    .S(net94),
    .X(_10605_));
 sky130_fd_sc_hd__clkbuf_1 _24786_ (.A(_10605_),
    .X(_02470_));
 sky130_fd_sc_hd__mux2_1 _24787_ (.A0(_10472_),
    .A1(\datamem.data_ram[47][27] ),
    .S(net94),
    .X(_10606_));
 sky130_fd_sc_hd__clkbuf_1 _24788_ (.A(_10606_),
    .X(_02471_));
 sky130_fd_sc_hd__mux2_1 _24789_ (.A0(_10474_),
    .A1(\datamem.data_ram[47][28] ),
    .S(net94),
    .X(_10607_));
 sky130_fd_sc_hd__clkbuf_1 _24790_ (.A(_10607_),
    .X(_02472_));
 sky130_fd_sc_hd__mux2_1 _24791_ (.A0(_10476_),
    .A1(\datamem.data_ram[47][29] ),
    .S(net94),
    .X(_10608_));
 sky130_fd_sc_hd__clkbuf_1 _24792_ (.A(_10608_),
    .X(_02473_));
 sky130_fd_sc_hd__mux2_1 _24793_ (.A0(_10478_),
    .A1(\datamem.data_ram[47][30] ),
    .S(_10602_),
    .X(_10609_));
 sky130_fd_sc_hd__clkbuf_1 _24794_ (.A(_10609_),
    .X(_02474_));
 sky130_fd_sc_hd__mux2_1 _24795_ (.A0(_10480_),
    .A1(\datamem.data_ram[47][31] ),
    .S(net94),
    .X(_10610_));
 sky130_fd_sc_hd__clkbuf_1 _24796_ (.A(_10610_),
    .X(_02475_));
 sky130_fd_sc_hd__buf_6 _24797_ (.A(_10500_),
    .X(_10611_));
 sky130_fd_sc_hd__a21oi_4 _24798_ (.A1(_10297_),
    .A2(_10337_),
    .B1(_10611_),
    .Y(_10612_));
 sky130_fd_sc_hd__mux2_1 _24799_ (.A0(_10439_),
    .A1(\datamem.data_ram[48][16] ),
    .S(_10612_),
    .X(_10613_));
 sky130_fd_sc_hd__clkbuf_1 _24800_ (.A(_10613_),
    .X(_02476_));
 sky130_fd_sc_hd__mux2_1 _24801_ (.A0(_10442_),
    .A1(\datamem.data_ram[48][17] ),
    .S(_10612_),
    .X(_10614_));
 sky130_fd_sc_hd__clkbuf_1 _24802_ (.A(_10614_),
    .X(_02477_));
 sky130_fd_sc_hd__mux2_1 _24803_ (.A0(_10444_),
    .A1(\datamem.data_ram[48][18] ),
    .S(_10612_),
    .X(_10615_));
 sky130_fd_sc_hd__clkbuf_1 _24804_ (.A(_10615_),
    .X(_02478_));
 sky130_fd_sc_hd__mux2_1 _24805_ (.A0(_10446_),
    .A1(\datamem.data_ram[48][19] ),
    .S(_10612_),
    .X(_10616_));
 sky130_fd_sc_hd__clkbuf_1 _24806_ (.A(_10616_),
    .X(_02479_));
 sky130_fd_sc_hd__mux2_1 _24807_ (.A0(_10448_),
    .A1(\datamem.data_ram[48][20] ),
    .S(_10612_),
    .X(_10617_));
 sky130_fd_sc_hd__clkbuf_1 _24808_ (.A(_10617_),
    .X(_02480_));
 sky130_fd_sc_hd__mux2_1 _24809_ (.A0(_10450_),
    .A1(\datamem.data_ram[48][21] ),
    .S(_10612_),
    .X(_10618_));
 sky130_fd_sc_hd__clkbuf_1 _24810_ (.A(_10618_),
    .X(_02481_));
 sky130_fd_sc_hd__mux2_1 _24811_ (.A0(_10452_),
    .A1(\datamem.data_ram[48][22] ),
    .S(_10612_),
    .X(_10619_));
 sky130_fd_sc_hd__clkbuf_1 _24812_ (.A(_10619_),
    .X(_02482_));
 sky130_fd_sc_hd__mux2_1 _24813_ (.A0(_10454_),
    .A1(\datamem.data_ram[48][23] ),
    .S(_10612_),
    .X(_10620_));
 sky130_fd_sc_hd__clkbuf_1 _24814_ (.A(_10620_),
    .X(_02483_));
 sky130_fd_sc_hd__a21oi_4 _24815_ (.A1(_10297_),
    .A2(_10347_),
    .B1(_10611_),
    .Y(_10621_));
 sky130_fd_sc_hd__mux2_1 _24816_ (.A0(_10385_),
    .A1(\datamem.data_ram[48][8] ),
    .S(_10621_),
    .X(_10622_));
 sky130_fd_sc_hd__clkbuf_1 _24817_ (.A(_10622_),
    .X(_02484_));
 sky130_fd_sc_hd__mux2_1 _24818_ (.A0(_10388_),
    .A1(\datamem.data_ram[48][9] ),
    .S(_10621_),
    .X(_10623_));
 sky130_fd_sc_hd__clkbuf_1 _24819_ (.A(_10623_),
    .X(_02485_));
 sky130_fd_sc_hd__mux2_1 _24820_ (.A0(_10390_),
    .A1(\datamem.data_ram[48][10] ),
    .S(_10621_),
    .X(_10624_));
 sky130_fd_sc_hd__clkbuf_1 _24821_ (.A(_10624_),
    .X(_02486_));
 sky130_fd_sc_hd__mux2_1 _24822_ (.A0(_10392_),
    .A1(\datamem.data_ram[48][11] ),
    .S(_10621_),
    .X(_10625_));
 sky130_fd_sc_hd__clkbuf_1 _24823_ (.A(_10625_),
    .X(_02487_));
 sky130_fd_sc_hd__mux2_1 _24824_ (.A0(_10394_),
    .A1(\datamem.data_ram[48][12] ),
    .S(_10621_),
    .X(_10626_));
 sky130_fd_sc_hd__clkbuf_1 _24825_ (.A(_10626_),
    .X(_02488_));
 sky130_fd_sc_hd__mux2_1 _24826_ (.A0(_10396_),
    .A1(\datamem.data_ram[48][13] ),
    .S(_10621_),
    .X(_10627_));
 sky130_fd_sc_hd__clkbuf_1 _24827_ (.A(_10627_),
    .X(_02489_));
 sky130_fd_sc_hd__mux2_1 _24828_ (.A0(_10398_),
    .A1(\datamem.data_ram[48][14] ),
    .S(_10621_),
    .X(_10628_));
 sky130_fd_sc_hd__clkbuf_1 _24829_ (.A(_10628_),
    .X(_02490_));
 sky130_fd_sc_hd__mux2_1 _24830_ (.A0(_10400_),
    .A1(\datamem.data_ram[48][15] ),
    .S(_10621_),
    .X(_10629_));
 sky130_fd_sc_hd__clkbuf_1 _24831_ (.A(_10629_),
    .X(_02491_));
 sky130_fd_sc_hd__nor2_8 _24832_ (.A(net104),
    .B(_10600_),
    .Y(_10630_));
 sky130_fd_sc_hd__a21oi_4 _24833_ (.A1(_10598_),
    .A2(_10630_),
    .B1(_10611_),
    .Y(_10631_));
 sky130_fd_sc_hd__mux2_1 _24834_ (.A0(_10439_),
    .A1(\datamem.data_ram[47][16] ),
    .S(_10631_),
    .X(_10632_));
 sky130_fd_sc_hd__clkbuf_1 _24835_ (.A(_10632_),
    .X(_02492_));
 sky130_fd_sc_hd__mux2_1 _24836_ (.A0(_10442_),
    .A1(\datamem.data_ram[47][17] ),
    .S(_10631_),
    .X(_10633_));
 sky130_fd_sc_hd__clkbuf_1 _24837_ (.A(_10633_),
    .X(_02493_));
 sky130_fd_sc_hd__mux2_1 _24838_ (.A0(_10444_),
    .A1(\datamem.data_ram[47][18] ),
    .S(_10631_),
    .X(_10634_));
 sky130_fd_sc_hd__clkbuf_1 _24839_ (.A(_10634_),
    .X(_02494_));
 sky130_fd_sc_hd__mux2_1 _24840_ (.A0(_10446_),
    .A1(\datamem.data_ram[47][19] ),
    .S(_10631_),
    .X(_10635_));
 sky130_fd_sc_hd__clkbuf_1 _24841_ (.A(_10635_),
    .X(_02495_));
 sky130_fd_sc_hd__mux2_1 _24842_ (.A0(_10448_),
    .A1(\datamem.data_ram[47][20] ),
    .S(_10631_),
    .X(_10636_));
 sky130_fd_sc_hd__clkbuf_1 _24843_ (.A(_10636_),
    .X(_02496_));
 sky130_fd_sc_hd__mux2_1 _24844_ (.A0(_10450_),
    .A1(\datamem.data_ram[47][21] ),
    .S(_10631_),
    .X(_10637_));
 sky130_fd_sc_hd__clkbuf_1 _24845_ (.A(_10637_),
    .X(_02497_));
 sky130_fd_sc_hd__mux2_1 _24846_ (.A0(_10452_),
    .A1(\datamem.data_ram[47][22] ),
    .S(_10631_),
    .X(_10638_));
 sky130_fd_sc_hd__clkbuf_1 _24847_ (.A(_10638_),
    .X(_02498_));
 sky130_fd_sc_hd__mux2_1 _24848_ (.A0(_10454_),
    .A1(\datamem.data_ram[47][23] ),
    .S(_10631_),
    .X(_10639_));
 sky130_fd_sc_hd__clkbuf_1 _24849_ (.A(_10639_),
    .X(_02499_));
 sky130_fd_sc_hd__nor2_8 _24850_ (.A(net112),
    .B(_10599_),
    .Y(_10640_));
 sky130_fd_sc_hd__a21oi_2 _24851_ (.A1(_10598_),
    .A2(_10640_),
    .B1(_10611_),
    .Y(_10641_));
 sky130_fd_sc_hd__mux2_1 _24852_ (.A0(_10385_),
    .A1(\datamem.data_ram[47][8] ),
    .S(net93),
    .X(_10642_));
 sky130_fd_sc_hd__clkbuf_1 _24853_ (.A(_10642_),
    .X(_02500_));
 sky130_fd_sc_hd__mux2_1 _24854_ (.A0(_10388_),
    .A1(\datamem.data_ram[47][9] ),
    .S(_10641_),
    .X(_10643_));
 sky130_fd_sc_hd__clkbuf_1 _24855_ (.A(_10643_),
    .X(_02501_));
 sky130_fd_sc_hd__mux2_1 _24856_ (.A0(_10390_),
    .A1(\datamem.data_ram[47][10] ),
    .S(net93),
    .X(_10644_));
 sky130_fd_sc_hd__clkbuf_1 _24857_ (.A(_10644_),
    .X(_02502_));
 sky130_fd_sc_hd__mux2_1 _24858_ (.A0(_10392_),
    .A1(\datamem.data_ram[47][11] ),
    .S(net93),
    .X(_10645_));
 sky130_fd_sc_hd__clkbuf_1 _24859_ (.A(_10645_),
    .X(_02503_));
 sky130_fd_sc_hd__mux2_1 _24860_ (.A0(_10394_),
    .A1(\datamem.data_ram[47][12] ),
    .S(net93),
    .X(_10646_));
 sky130_fd_sc_hd__clkbuf_1 _24861_ (.A(_10646_),
    .X(_02504_));
 sky130_fd_sc_hd__mux2_1 _24862_ (.A0(_10396_),
    .A1(\datamem.data_ram[47][13] ),
    .S(net93),
    .X(_10647_));
 sky130_fd_sc_hd__clkbuf_1 _24863_ (.A(_10647_),
    .X(_02505_));
 sky130_fd_sc_hd__mux2_1 _24864_ (.A0(_10398_),
    .A1(\datamem.data_ram[47][14] ),
    .S(_10641_),
    .X(_10648_));
 sky130_fd_sc_hd__clkbuf_1 _24865_ (.A(_10648_),
    .X(_02506_));
 sky130_fd_sc_hd__mux2_1 _24866_ (.A0(_10400_),
    .A1(\datamem.data_ram[47][15] ),
    .S(_10641_),
    .X(_10649_));
 sky130_fd_sc_hd__clkbuf_1 _24867_ (.A(_10649_),
    .X(_02507_));
 sky130_fd_sc_hd__a21oi_1 _24868_ (.A1(_09226_),
    .A2(_10601_),
    .B1(_10611_),
    .Y(_10650_));
 sky130_fd_sc_hd__mux2_1 _24869_ (.A0(_10465_),
    .A1(\datamem.data_ram[46][24] ),
    .S(net92),
    .X(_10651_));
 sky130_fd_sc_hd__clkbuf_1 _24870_ (.A(_10651_),
    .X(_02508_));
 sky130_fd_sc_hd__mux2_1 _24871_ (.A0(_10468_),
    .A1(\datamem.data_ram[46][25] ),
    .S(net92),
    .X(_10652_));
 sky130_fd_sc_hd__clkbuf_1 _24872_ (.A(_10652_),
    .X(_02509_));
 sky130_fd_sc_hd__mux2_1 _24873_ (.A0(_10470_),
    .A1(\datamem.data_ram[46][26] ),
    .S(net92),
    .X(_10653_));
 sky130_fd_sc_hd__clkbuf_1 _24874_ (.A(_10653_),
    .X(_02510_));
 sky130_fd_sc_hd__mux2_1 _24875_ (.A0(_10472_),
    .A1(\datamem.data_ram[46][27] ),
    .S(net92),
    .X(_10654_));
 sky130_fd_sc_hd__clkbuf_1 _24876_ (.A(_10654_),
    .X(_02511_));
 sky130_fd_sc_hd__mux2_1 _24877_ (.A0(_10474_),
    .A1(\datamem.data_ram[46][28] ),
    .S(net92),
    .X(_10655_));
 sky130_fd_sc_hd__clkbuf_1 _24878_ (.A(_10655_),
    .X(_02512_));
 sky130_fd_sc_hd__mux2_1 _24879_ (.A0(_10476_),
    .A1(\datamem.data_ram[46][29] ),
    .S(net92),
    .X(_10656_));
 sky130_fd_sc_hd__clkbuf_1 _24880_ (.A(_10656_),
    .X(_02513_));
 sky130_fd_sc_hd__mux2_1 _24881_ (.A0(_10478_),
    .A1(\datamem.data_ram[46][30] ),
    .S(_10650_),
    .X(_10657_));
 sky130_fd_sc_hd__clkbuf_1 _24882_ (.A(_10657_),
    .X(_02514_));
 sky130_fd_sc_hd__mux2_1 _24883_ (.A0(_10480_),
    .A1(\datamem.data_ram[46][31] ),
    .S(net92),
    .X(_10658_));
 sky130_fd_sc_hd__clkbuf_1 _24884_ (.A(_10658_),
    .X(_02515_));
 sky130_fd_sc_hd__a21oi_4 _24885_ (.A1(_09226_),
    .A2(_10630_),
    .B1(_10611_),
    .Y(_10659_));
 sky130_fd_sc_hd__mux2_1 _24886_ (.A0(_10439_),
    .A1(\datamem.data_ram[46][16] ),
    .S(_10659_),
    .X(_10660_));
 sky130_fd_sc_hd__clkbuf_1 _24887_ (.A(_10660_),
    .X(_02516_));
 sky130_fd_sc_hd__mux2_1 _24888_ (.A0(_10442_),
    .A1(\datamem.data_ram[46][17] ),
    .S(_10659_),
    .X(_10661_));
 sky130_fd_sc_hd__clkbuf_1 _24889_ (.A(_10661_),
    .X(_02517_));
 sky130_fd_sc_hd__mux2_1 _24890_ (.A0(_10444_),
    .A1(\datamem.data_ram[46][18] ),
    .S(_10659_),
    .X(_10662_));
 sky130_fd_sc_hd__clkbuf_1 _24891_ (.A(_10662_),
    .X(_02518_));
 sky130_fd_sc_hd__mux2_1 _24892_ (.A0(_10446_),
    .A1(\datamem.data_ram[46][19] ),
    .S(_10659_),
    .X(_10663_));
 sky130_fd_sc_hd__clkbuf_1 _24893_ (.A(_10663_),
    .X(_02519_));
 sky130_fd_sc_hd__mux2_1 _24894_ (.A0(_10448_),
    .A1(\datamem.data_ram[46][20] ),
    .S(_10659_),
    .X(_10664_));
 sky130_fd_sc_hd__clkbuf_1 _24895_ (.A(_10664_),
    .X(_02520_));
 sky130_fd_sc_hd__mux2_1 _24896_ (.A0(_10450_),
    .A1(\datamem.data_ram[46][21] ),
    .S(_10659_),
    .X(_10665_));
 sky130_fd_sc_hd__clkbuf_1 _24897_ (.A(_10665_),
    .X(_02521_));
 sky130_fd_sc_hd__mux2_1 _24898_ (.A0(_10452_),
    .A1(\datamem.data_ram[46][22] ),
    .S(_10659_),
    .X(_10666_));
 sky130_fd_sc_hd__clkbuf_1 _24899_ (.A(_10666_),
    .X(_02522_));
 sky130_fd_sc_hd__mux2_1 _24900_ (.A0(_10454_),
    .A1(\datamem.data_ram[46][23] ),
    .S(_10659_),
    .X(_10667_));
 sky130_fd_sc_hd__clkbuf_1 _24901_ (.A(_10667_),
    .X(_02523_));
 sky130_fd_sc_hd__buf_8 _24902_ (.A(_09225_),
    .X(_10668_));
 sky130_fd_sc_hd__a21oi_4 _24903_ (.A1(_10668_),
    .A2(_10640_),
    .B1(_10611_),
    .Y(_10669_));
 sky130_fd_sc_hd__mux2_1 _24904_ (.A0(_10385_),
    .A1(\datamem.data_ram[46][8] ),
    .S(_10669_),
    .X(_10670_));
 sky130_fd_sc_hd__clkbuf_1 _24905_ (.A(_10670_),
    .X(_02524_));
 sky130_fd_sc_hd__mux2_1 _24906_ (.A0(_10388_),
    .A1(\datamem.data_ram[46][9] ),
    .S(_10669_),
    .X(_10671_));
 sky130_fd_sc_hd__clkbuf_1 _24907_ (.A(_10671_),
    .X(_02525_));
 sky130_fd_sc_hd__mux2_1 _24908_ (.A0(_10390_),
    .A1(\datamem.data_ram[46][10] ),
    .S(_10669_),
    .X(_10672_));
 sky130_fd_sc_hd__clkbuf_1 _24909_ (.A(_10672_),
    .X(_02526_));
 sky130_fd_sc_hd__mux2_1 _24910_ (.A0(_10392_),
    .A1(\datamem.data_ram[46][11] ),
    .S(_10669_),
    .X(_10673_));
 sky130_fd_sc_hd__clkbuf_1 _24911_ (.A(_10673_),
    .X(_02527_));
 sky130_fd_sc_hd__mux2_1 _24912_ (.A0(_10394_),
    .A1(\datamem.data_ram[46][12] ),
    .S(_10669_),
    .X(_10674_));
 sky130_fd_sc_hd__clkbuf_1 _24913_ (.A(_10674_),
    .X(_02528_));
 sky130_fd_sc_hd__mux2_1 _24914_ (.A0(_10396_),
    .A1(\datamem.data_ram[46][13] ),
    .S(_10669_),
    .X(_10675_));
 sky130_fd_sc_hd__clkbuf_1 _24915_ (.A(_10675_),
    .X(_02529_));
 sky130_fd_sc_hd__mux2_1 _24916_ (.A0(_10398_),
    .A1(\datamem.data_ram[46][14] ),
    .S(_10669_),
    .X(_10676_));
 sky130_fd_sc_hd__clkbuf_1 _24917_ (.A(_10676_),
    .X(_02530_));
 sky130_fd_sc_hd__mux2_1 _24918_ (.A0(_10400_),
    .A1(\datamem.data_ram[46][15] ),
    .S(_10669_),
    .X(_10677_));
 sky130_fd_sc_hd__clkbuf_1 _24919_ (.A(_10677_),
    .X(_02531_));
 sky130_fd_sc_hd__a21oi_1 _24920_ (.A1(_10113_),
    .A2(_10601_),
    .B1(_10611_),
    .Y(_10678_));
 sky130_fd_sc_hd__mux2_1 _24921_ (.A0(_10465_),
    .A1(\datamem.data_ram[45][24] ),
    .S(net91),
    .X(_10679_));
 sky130_fd_sc_hd__clkbuf_1 _24922_ (.A(_10679_),
    .X(_02532_));
 sky130_fd_sc_hd__mux2_1 _24923_ (.A0(_10468_),
    .A1(\datamem.data_ram[45][25] ),
    .S(net91),
    .X(_10680_));
 sky130_fd_sc_hd__clkbuf_1 _24924_ (.A(_10680_),
    .X(_02533_));
 sky130_fd_sc_hd__mux2_1 _24925_ (.A0(_10470_),
    .A1(\datamem.data_ram[45][26] ),
    .S(net91),
    .X(_10681_));
 sky130_fd_sc_hd__clkbuf_1 _24926_ (.A(_10681_),
    .X(_02534_));
 sky130_fd_sc_hd__mux2_1 _24927_ (.A0(_10472_),
    .A1(\datamem.data_ram[45][27] ),
    .S(net91),
    .X(_10682_));
 sky130_fd_sc_hd__clkbuf_1 _24928_ (.A(_10682_),
    .X(_02535_));
 sky130_fd_sc_hd__mux2_1 _24929_ (.A0(_10474_),
    .A1(\datamem.data_ram[45][28] ),
    .S(net91),
    .X(_10683_));
 sky130_fd_sc_hd__clkbuf_1 _24930_ (.A(_10683_),
    .X(_02536_));
 sky130_fd_sc_hd__mux2_1 _24931_ (.A0(_10476_),
    .A1(\datamem.data_ram[45][29] ),
    .S(net91),
    .X(_10684_));
 sky130_fd_sc_hd__clkbuf_1 _24932_ (.A(_10684_),
    .X(_02537_));
 sky130_fd_sc_hd__mux2_1 _24933_ (.A0(_10478_),
    .A1(\datamem.data_ram[45][30] ),
    .S(_10678_),
    .X(_10685_));
 sky130_fd_sc_hd__clkbuf_1 _24934_ (.A(_10685_),
    .X(_02538_));
 sky130_fd_sc_hd__mux2_1 _24935_ (.A0(_10480_),
    .A1(\datamem.data_ram[45][31] ),
    .S(net91),
    .X(_10686_));
 sky130_fd_sc_hd__clkbuf_1 _24936_ (.A(_10686_),
    .X(_02539_));
 sky130_fd_sc_hd__a21oi_4 _24937_ (.A1(_10113_),
    .A2(_10630_),
    .B1(_10611_),
    .Y(_10687_));
 sky130_fd_sc_hd__mux2_1 _24938_ (.A0(_10439_),
    .A1(\datamem.data_ram[45][16] ),
    .S(_10687_),
    .X(_10688_));
 sky130_fd_sc_hd__clkbuf_1 _24939_ (.A(_10688_),
    .X(_02540_));
 sky130_fd_sc_hd__mux2_1 _24940_ (.A0(_10442_),
    .A1(\datamem.data_ram[45][17] ),
    .S(_10687_),
    .X(_10689_));
 sky130_fd_sc_hd__clkbuf_1 _24941_ (.A(_10689_),
    .X(_02541_));
 sky130_fd_sc_hd__mux2_1 _24942_ (.A0(_10444_),
    .A1(\datamem.data_ram[45][18] ),
    .S(_10687_),
    .X(_10690_));
 sky130_fd_sc_hd__clkbuf_1 _24943_ (.A(_10690_),
    .X(_02542_));
 sky130_fd_sc_hd__mux2_1 _24944_ (.A0(_10446_),
    .A1(\datamem.data_ram[45][19] ),
    .S(_10687_),
    .X(_10691_));
 sky130_fd_sc_hd__clkbuf_1 _24945_ (.A(_10691_),
    .X(_02543_));
 sky130_fd_sc_hd__mux2_1 _24946_ (.A0(_10448_),
    .A1(\datamem.data_ram[45][20] ),
    .S(_10687_),
    .X(_10692_));
 sky130_fd_sc_hd__clkbuf_1 _24947_ (.A(_10692_),
    .X(_02544_));
 sky130_fd_sc_hd__mux2_1 _24948_ (.A0(_10450_),
    .A1(\datamem.data_ram[45][21] ),
    .S(_10687_),
    .X(_10693_));
 sky130_fd_sc_hd__clkbuf_1 _24949_ (.A(_10693_),
    .X(_02545_));
 sky130_fd_sc_hd__mux2_1 _24950_ (.A0(_10452_),
    .A1(\datamem.data_ram[45][22] ),
    .S(_10687_),
    .X(_10694_));
 sky130_fd_sc_hd__clkbuf_1 _24951_ (.A(_10694_),
    .X(_02546_));
 sky130_fd_sc_hd__mux2_1 _24952_ (.A0(_10454_),
    .A1(\datamem.data_ram[45][23] ),
    .S(_10687_),
    .X(_10695_));
 sky130_fd_sc_hd__clkbuf_1 _24953_ (.A(_10695_),
    .X(_02547_));
 sky130_fd_sc_hd__a21oi_4 _24954_ (.A1(_10113_),
    .A2(_10640_),
    .B1(_10611_),
    .Y(_10696_));
 sky130_fd_sc_hd__mux2_1 _24955_ (.A0(_10385_),
    .A1(\datamem.data_ram[45][8] ),
    .S(_10696_),
    .X(_10697_));
 sky130_fd_sc_hd__clkbuf_1 _24956_ (.A(_10697_),
    .X(_02548_));
 sky130_fd_sc_hd__mux2_1 _24957_ (.A0(_10388_),
    .A1(\datamem.data_ram[45][9] ),
    .S(_10696_),
    .X(_10698_));
 sky130_fd_sc_hd__clkbuf_1 _24958_ (.A(_10698_),
    .X(_02549_));
 sky130_fd_sc_hd__mux2_1 _24959_ (.A0(_10390_),
    .A1(\datamem.data_ram[45][10] ),
    .S(_10696_),
    .X(_10699_));
 sky130_fd_sc_hd__clkbuf_1 _24960_ (.A(_10699_),
    .X(_02550_));
 sky130_fd_sc_hd__mux2_1 _24961_ (.A0(_10392_),
    .A1(\datamem.data_ram[45][11] ),
    .S(_10696_),
    .X(_10700_));
 sky130_fd_sc_hd__clkbuf_1 _24962_ (.A(_10700_),
    .X(_02551_));
 sky130_fd_sc_hd__mux2_1 _24963_ (.A0(_10394_),
    .A1(\datamem.data_ram[45][12] ),
    .S(_10696_),
    .X(_10701_));
 sky130_fd_sc_hd__clkbuf_1 _24964_ (.A(_10701_),
    .X(_02552_));
 sky130_fd_sc_hd__mux2_1 _24965_ (.A0(_10396_),
    .A1(\datamem.data_ram[45][13] ),
    .S(_10696_),
    .X(_10702_));
 sky130_fd_sc_hd__clkbuf_1 _24966_ (.A(_10702_),
    .X(_02553_));
 sky130_fd_sc_hd__mux2_1 _24967_ (.A0(_10398_),
    .A1(\datamem.data_ram[45][14] ),
    .S(_10696_),
    .X(_10703_));
 sky130_fd_sc_hd__clkbuf_1 _24968_ (.A(_10703_),
    .X(_02554_));
 sky130_fd_sc_hd__mux2_1 _24969_ (.A0(_10400_),
    .A1(\datamem.data_ram[45][15] ),
    .S(_10696_),
    .X(_10704_));
 sky130_fd_sc_hd__clkbuf_1 _24970_ (.A(_10704_),
    .X(_02555_));
 sky130_fd_sc_hd__buf_6 _24971_ (.A(_10500_),
    .X(_10705_));
 sky130_fd_sc_hd__a21oi_1 _24972_ (.A1(_10542_),
    .A2(_10601_),
    .B1(_10705_),
    .Y(_10706_));
 sky130_fd_sc_hd__mux2_1 _24973_ (.A0(_10465_),
    .A1(\datamem.data_ram[44][24] ),
    .S(net101),
    .X(_10707_));
 sky130_fd_sc_hd__clkbuf_1 _24974_ (.A(_10707_),
    .X(_02556_));
 sky130_fd_sc_hd__mux2_1 _24975_ (.A0(_10468_),
    .A1(\datamem.data_ram[44][25] ),
    .S(net101),
    .X(_10708_));
 sky130_fd_sc_hd__clkbuf_1 _24976_ (.A(_10708_),
    .X(_02557_));
 sky130_fd_sc_hd__mux2_1 _24977_ (.A0(_10470_),
    .A1(\datamem.data_ram[44][26] ),
    .S(net101),
    .X(_10709_));
 sky130_fd_sc_hd__clkbuf_1 _24978_ (.A(_10709_),
    .X(_02558_));
 sky130_fd_sc_hd__mux2_1 _24979_ (.A0(_10472_),
    .A1(\datamem.data_ram[44][27] ),
    .S(net101),
    .X(_10710_));
 sky130_fd_sc_hd__clkbuf_1 _24980_ (.A(_10710_),
    .X(_02559_));
 sky130_fd_sc_hd__mux2_1 _24981_ (.A0(_10474_),
    .A1(\datamem.data_ram[44][28] ),
    .S(net101),
    .X(_10711_));
 sky130_fd_sc_hd__clkbuf_1 _24982_ (.A(_10711_),
    .X(_02560_));
 sky130_fd_sc_hd__mux2_1 _24983_ (.A0(_10476_),
    .A1(\datamem.data_ram[44][29] ),
    .S(net101),
    .X(_10712_));
 sky130_fd_sc_hd__clkbuf_1 _24984_ (.A(_10712_),
    .X(_02561_));
 sky130_fd_sc_hd__mux2_1 _24985_ (.A0(_10478_),
    .A1(\datamem.data_ram[44][30] ),
    .S(_10706_),
    .X(_10713_));
 sky130_fd_sc_hd__clkbuf_1 _24986_ (.A(_10713_),
    .X(_02562_));
 sky130_fd_sc_hd__mux2_1 _24987_ (.A0(_10480_),
    .A1(\datamem.data_ram[44][31] ),
    .S(net101),
    .X(_10714_));
 sky130_fd_sc_hd__clkbuf_1 _24988_ (.A(_10714_),
    .X(_02563_));
 sky130_fd_sc_hd__a21oi_4 _24989_ (.A1(_10542_),
    .A2(_10630_),
    .B1(_10705_),
    .Y(_10715_));
 sky130_fd_sc_hd__mux2_1 _24990_ (.A0(_10439_),
    .A1(\datamem.data_ram[44][16] ),
    .S(_10715_),
    .X(_10716_));
 sky130_fd_sc_hd__clkbuf_1 _24991_ (.A(_10716_),
    .X(_02564_));
 sky130_fd_sc_hd__mux2_1 _24992_ (.A0(_10442_),
    .A1(\datamem.data_ram[44][17] ),
    .S(_10715_),
    .X(_10717_));
 sky130_fd_sc_hd__clkbuf_1 _24993_ (.A(_10717_),
    .X(_02565_));
 sky130_fd_sc_hd__mux2_1 _24994_ (.A0(_10444_),
    .A1(\datamem.data_ram[44][18] ),
    .S(_10715_),
    .X(_10718_));
 sky130_fd_sc_hd__clkbuf_1 _24995_ (.A(_10718_),
    .X(_02566_));
 sky130_fd_sc_hd__mux2_1 _24996_ (.A0(_10446_),
    .A1(\datamem.data_ram[44][19] ),
    .S(_10715_),
    .X(_10719_));
 sky130_fd_sc_hd__clkbuf_1 _24997_ (.A(_10719_),
    .X(_02567_));
 sky130_fd_sc_hd__mux2_1 _24998_ (.A0(_10448_),
    .A1(\datamem.data_ram[44][20] ),
    .S(_10715_),
    .X(_10720_));
 sky130_fd_sc_hd__clkbuf_1 _24999_ (.A(_10720_),
    .X(_02568_));
 sky130_fd_sc_hd__mux2_1 _25000_ (.A0(_10450_),
    .A1(\datamem.data_ram[44][21] ),
    .S(_10715_),
    .X(_10721_));
 sky130_fd_sc_hd__clkbuf_1 _25001_ (.A(_10721_),
    .X(_02569_));
 sky130_fd_sc_hd__mux2_1 _25002_ (.A0(_10452_),
    .A1(\datamem.data_ram[44][22] ),
    .S(_10715_),
    .X(_10722_));
 sky130_fd_sc_hd__clkbuf_1 _25003_ (.A(_10722_),
    .X(_02570_));
 sky130_fd_sc_hd__mux2_1 _25004_ (.A0(_10454_),
    .A1(\datamem.data_ram[44][23] ),
    .S(_10715_),
    .X(_10723_));
 sky130_fd_sc_hd__clkbuf_1 _25005_ (.A(_10723_),
    .X(_02571_));
 sky130_fd_sc_hd__buf_2 _25006_ (.A(_09266_),
    .X(_10724_));
 sky130_fd_sc_hd__a21oi_4 _25007_ (.A1(_10542_),
    .A2(_10640_),
    .B1(_10705_),
    .Y(_10725_));
 sky130_fd_sc_hd__mux2_1 _25008_ (.A0(_10724_),
    .A1(\datamem.data_ram[44][8] ),
    .S(net100),
    .X(_10726_));
 sky130_fd_sc_hd__clkbuf_1 _25009_ (.A(_10726_),
    .X(_02572_));
 sky130_fd_sc_hd__buf_2 _25010_ (.A(_09272_),
    .X(_10727_));
 sky130_fd_sc_hd__mux2_1 _25011_ (.A0(_10727_),
    .A1(\datamem.data_ram[44][9] ),
    .S(_10725_),
    .X(_10728_));
 sky130_fd_sc_hd__clkbuf_1 _25012_ (.A(_10728_),
    .X(_02573_));
 sky130_fd_sc_hd__buf_2 _25013_ (.A(_09275_),
    .X(_10729_));
 sky130_fd_sc_hd__mux2_1 _25014_ (.A0(_10729_),
    .A1(\datamem.data_ram[44][10] ),
    .S(net100),
    .X(_10730_));
 sky130_fd_sc_hd__clkbuf_1 _25015_ (.A(_10730_),
    .X(_02574_));
 sky130_fd_sc_hd__clkbuf_2 _25016_ (.A(_09278_),
    .X(_10731_));
 sky130_fd_sc_hd__mux2_1 _25017_ (.A0(_10731_),
    .A1(\datamem.data_ram[44][11] ),
    .S(net100),
    .X(_10732_));
 sky130_fd_sc_hd__clkbuf_1 _25018_ (.A(_10732_),
    .X(_02575_));
 sky130_fd_sc_hd__buf_2 _25019_ (.A(_09281_),
    .X(_10733_));
 sky130_fd_sc_hd__mux2_1 _25020_ (.A0(_10733_),
    .A1(\datamem.data_ram[44][12] ),
    .S(net100),
    .X(_10734_));
 sky130_fd_sc_hd__clkbuf_1 _25021_ (.A(_10734_),
    .X(_02576_));
 sky130_fd_sc_hd__buf_2 _25022_ (.A(_09284_),
    .X(_10735_));
 sky130_fd_sc_hd__mux2_1 _25023_ (.A0(_10735_),
    .A1(\datamem.data_ram[44][13] ),
    .S(net100),
    .X(_10736_));
 sky130_fd_sc_hd__clkbuf_1 _25024_ (.A(_10736_),
    .X(_02577_));
 sky130_fd_sc_hd__buf_2 _25025_ (.A(_09287_),
    .X(_10737_));
 sky130_fd_sc_hd__mux2_1 _25026_ (.A0(_10737_),
    .A1(\datamem.data_ram[44][14] ),
    .S(_10725_),
    .X(_10738_));
 sky130_fd_sc_hd__clkbuf_1 _25027_ (.A(_10738_),
    .X(_02578_));
 sky130_fd_sc_hd__buf_2 _25028_ (.A(_09290_),
    .X(_10739_));
 sky130_fd_sc_hd__mux2_1 _25029_ (.A0(_10739_),
    .A1(\datamem.data_ram[44][15] ),
    .S(_10725_),
    .X(_10740_));
 sky130_fd_sc_hd__clkbuf_1 _25030_ (.A(_10740_),
    .X(_02579_));
 sky130_fd_sc_hd__buf_8 _25031_ (.A(_07137_),
    .X(_10741_));
 sky130_fd_sc_hd__a21oi_1 _25032_ (.A1(_10741_),
    .A2(_10601_),
    .B1(_10705_),
    .Y(_10742_));
 sky130_fd_sc_hd__mux2_1 _25033_ (.A0(_10465_),
    .A1(\datamem.data_ram[43][24] ),
    .S(net90),
    .X(_10743_));
 sky130_fd_sc_hd__clkbuf_1 _25034_ (.A(_10743_),
    .X(_02580_));
 sky130_fd_sc_hd__mux2_1 _25035_ (.A0(_10468_),
    .A1(\datamem.data_ram[43][25] ),
    .S(net90),
    .X(_10744_));
 sky130_fd_sc_hd__clkbuf_1 _25036_ (.A(_10744_),
    .X(_02581_));
 sky130_fd_sc_hd__mux2_1 _25037_ (.A0(_10470_),
    .A1(\datamem.data_ram[43][26] ),
    .S(net90),
    .X(_10745_));
 sky130_fd_sc_hd__clkbuf_1 _25038_ (.A(_10745_),
    .X(_02582_));
 sky130_fd_sc_hd__mux2_1 _25039_ (.A0(_10472_),
    .A1(\datamem.data_ram[43][27] ),
    .S(net90),
    .X(_10746_));
 sky130_fd_sc_hd__clkbuf_1 _25040_ (.A(_10746_),
    .X(_02583_));
 sky130_fd_sc_hd__mux2_1 _25041_ (.A0(_10474_),
    .A1(\datamem.data_ram[43][28] ),
    .S(net90),
    .X(_10747_));
 sky130_fd_sc_hd__clkbuf_1 _25042_ (.A(_10747_),
    .X(_02584_));
 sky130_fd_sc_hd__mux2_1 _25043_ (.A0(_10476_),
    .A1(\datamem.data_ram[43][29] ),
    .S(net90),
    .X(_10748_));
 sky130_fd_sc_hd__clkbuf_1 _25044_ (.A(_10748_),
    .X(_02585_));
 sky130_fd_sc_hd__mux2_1 _25045_ (.A0(_10478_),
    .A1(\datamem.data_ram[43][30] ),
    .S(_10742_),
    .X(_10749_));
 sky130_fd_sc_hd__clkbuf_1 _25046_ (.A(_10749_),
    .X(_02586_));
 sky130_fd_sc_hd__mux2_1 _25047_ (.A0(_10480_),
    .A1(\datamem.data_ram[43][31] ),
    .S(net90),
    .X(_10750_));
 sky130_fd_sc_hd__clkbuf_1 _25048_ (.A(_10750_),
    .X(_02587_));
 sky130_fd_sc_hd__buf_2 _25049_ (.A(_09223_),
    .X(_10751_));
 sky130_fd_sc_hd__a21oi_4 _25050_ (.A1(_10741_),
    .A2(_10630_),
    .B1(_10705_),
    .Y(_10752_));
 sky130_fd_sc_hd__mux2_1 _25051_ (.A0(_10751_),
    .A1(\datamem.data_ram[43][16] ),
    .S(_10752_),
    .X(_10753_));
 sky130_fd_sc_hd__clkbuf_1 _25052_ (.A(_10753_),
    .X(_02588_));
 sky130_fd_sc_hd__buf_2 _25053_ (.A(_09235_),
    .X(_10754_));
 sky130_fd_sc_hd__mux2_1 _25054_ (.A0(_10754_),
    .A1(\datamem.data_ram[43][17] ),
    .S(_10752_),
    .X(_10755_));
 sky130_fd_sc_hd__clkbuf_1 _25055_ (.A(_10755_),
    .X(_02589_));
 sky130_fd_sc_hd__buf_2 _25056_ (.A(_09239_),
    .X(_10756_));
 sky130_fd_sc_hd__mux2_1 _25057_ (.A0(_10756_),
    .A1(\datamem.data_ram[43][18] ),
    .S(_10752_),
    .X(_10757_));
 sky130_fd_sc_hd__clkbuf_1 _25058_ (.A(_10757_),
    .X(_02590_));
 sky130_fd_sc_hd__buf_2 _25059_ (.A(_09243_),
    .X(_10758_));
 sky130_fd_sc_hd__mux2_1 _25060_ (.A0(_10758_),
    .A1(\datamem.data_ram[43][19] ),
    .S(_10752_),
    .X(_10759_));
 sky130_fd_sc_hd__clkbuf_1 _25061_ (.A(_10759_),
    .X(_02591_));
 sky130_fd_sc_hd__buf_2 _25062_ (.A(_09247_),
    .X(_10760_));
 sky130_fd_sc_hd__mux2_1 _25063_ (.A0(_10760_),
    .A1(\datamem.data_ram[43][20] ),
    .S(_10752_),
    .X(_10761_));
 sky130_fd_sc_hd__clkbuf_1 _25064_ (.A(_10761_),
    .X(_02592_));
 sky130_fd_sc_hd__buf_2 _25065_ (.A(_09251_),
    .X(_10762_));
 sky130_fd_sc_hd__mux2_1 _25066_ (.A0(_10762_),
    .A1(\datamem.data_ram[43][21] ),
    .S(_10752_),
    .X(_10763_));
 sky130_fd_sc_hd__clkbuf_1 _25067_ (.A(_10763_),
    .X(_02593_));
 sky130_fd_sc_hd__buf_2 _25068_ (.A(_09255_),
    .X(_10764_));
 sky130_fd_sc_hd__mux2_1 _25069_ (.A0(_10764_),
    .A1(\datamem.data_ram[43][22] ),
    .S(_10752_),
    .X(_10765_));
 sky130_fd_sc_hd__clkbuf_1 _25070_ (.A(_10765_),
    .X(_02594_));
 sky130_fd_sc_hd__buf_2 _25071_ (.A(_09259_),
    .X(_10766_));
 sky130_fd_sc_hd__mux2_1 _25072_ (.A0(_10766_),
    .A1(\datamem.data_ram[43][23] ),
    .S(_10752_),
    .X(_10767_));
 sky130_fd_sc_hd__clkbuf_1 _25073_ (.A(_10767_),
    .X(_02595_));
 sky130_fd_sc_hd__a21oi_4 _25074_ (.A1(_10741_),
    .A2(_10640_),
    .B1(_10705_),
    .Y(_10768_));
 sky130_fd_sc_hd__mux2_1 _25075_ (.A0(_10724_),
    .A1(\datamem.data_ram[43][8] ),
    .S(net89),
    .X(_10769_));
 sky130_fd_sc_hd__clkbuf_1 _25076_ (.A(_10769_),
    .X(_02596_));
 sky130_fd_sc_hd__mux2_1 _25077_ (.A0(_10727_),
    .A1(\datamem.data_ram[43][9] ),
    .S(_10768_),
    .X(_10770_));
 sky130_fd_sc_hd__clkbuf_1 _25078_ (.A(_10770_),
    .X(_02597_));
 sky130_fd_sc_hd__mux2_1 _25079_ (.A0(_10729_),
    .A1(\datamem.data_ram[43][10] ),
    .S(net89),
    .X(_10771_));
 sky130_fd_sc_hd__clkbuf_1 _25080_ (.A(_10771_),
    .X(_02598_));
 sky130_fd_sc_hd__mux2_1 _25081_ (.A0(_10731_),
    .A1(\datamem.data_ram[43][11] ),
    .S(net89),
    .X(_10772_));
 sky130_fd_sc_hd__clkbuf_1 _25082_ (.A(_10772_),
    .X(_02599_));
 sky130_fd_sc_hd__mux2_1 _25083_ (.A0(_10733_),
    .A1(\datamem.data_ram[43][12] ),
    .S(net89),
    .X(_10773_));
 sky130_fd_sc_hd__clkbuf_1 _25084_ (.A(_10773_),
    .X(_02600_));
 sky130_fd_sc_hd__mux2_1 _25085_ (.A0(_10735_),
    .A1(\datamem.data_ram[43][13] ),
    .S(net89),
    .X(_10774_));
 sky130_fd_sc_hd__clkbuf_1 _25086_ (.A(_10774_),
    .X(_02601_));
 sky130_fd_sc_hd__mux2_1 _25087_ (.A0(_10737_),
    .A1(\datamem.data_ram[43][14] ),
    .S(_10768_),
    .X(_10775_));
 sky130_fd_sc_hd__clkbuf_1 _25088_ (.A(_10775_),
    .X(_02602_));
 sky130_fd_sc_hd__mux2_1 _25089_ (.A0(_10739_),
    .A1(\datamem.data_ram[43][15] ),
    .S(_10768_),
    .X(_10776_));
 sky130_fd_sc_hd__clkbuf_1 _25090_ (.A(_10776_),
    .X(_02603_));
 sky130_fd_sc_hd__buf_8 _25091_ (.A(_07136_),
    .X(_10777_));
 sky130_fd_sc_hd__nand2_4 _25092_ (.A(_10777_),
    .B(_10051_),
    .Y(_10778_));
 sky130_fd_sc_hd__nor2_2 _25093_ (.A(_10600_),
    .B(_10778_),
    .Y(_10779_));
 sky130_fd_sc_hd__buf_4 _25094_ (.A(_09231_),
    .X(_10780_));
 sky130_fd_sc_hd__nor2_2 _25095_ (.A(_10780_),
    .B(_10779_),
    .Y(_10781_));
 sky130_fd_sc_hd__a22o_1 _25096_ (.A1(_10048_),
    .A2(_10779_),
    .B1(_10781_),
    .B2(\datamem.data_ram[42][0] ),
    .X(_02604_));
 sky130_fd_sc_hd__a22o_1 _25097_ (.A1(_10058_),
    .A2(_10779_),
    .B1(_10781_),
    .B2(\datamem.data_ram[42][1] ),
    .X(_02605_));
 sky130_fd_sc_hd__a22o_1 _25098_ (.A1(_10061_),
    .A2(_10779_),
    .B1(_10781_),
    .B2(\datamem.data_ram[42][2] ),
    .X(_02606_));
 sky130_fd_sc_hd__a22o_1 _25099_ (.A1(_10064_),
    .A2(_10779_),
    .B1(_10781_),
    .B2(\datamem.data_ram[42][3] ),
    .X(_02607_));
 sky130_fd_sc_hd__clkbuf_4 _25100_ (.A(_10067_),
    .X(_10782_));
 sky130_fd_sc_hd__a22o_1 _25101_ (.A1(_10782_),
    .A2(_10779_),
    .B1(_10781_),
    .B2(\datamem.data_ram[42][4] ),
    .X(_02608_));
 sky130_fd_sc_hd__a22o_1 _25102_ (.A1(_10070_),
    .A2(_10779_),
    .B1(_10781_),
    .B2(\datamem.data_ram[42][5] ),
    .X(_02609_));
 sky130_fd_sc_hd__a22o_1 _25103_ (.A1(_10073_),
    .A2(_10779_),
    .B1(_10781_),
    .B2(\datamem.data_ram[42][6] ),
    .X(_02610_));
 sky130_fd_sc_hd__clkbuf_4 _25104_ (.A(_10075_),
    .X(_10783_));
 sky130_fd_sc_hd__a22o_1 _25105_ (.A1(_10783_),
    .A2(_10779_),
    .B1(_10781_),
    .B2(\datamem.data_ram[42][7] ),
    .X(_02611_));
 sky130_fd_sc_hd__a21oi_4 _25106_ (.A1(_10520_),
    .A2(_10640_),
    .B1(_10705_),
    .Y(_10784_));
 sky130_fd_sc_hd__mux2_1 _25107_ (.A0(_10724_),
    .A1(\datamem.data_ram[42][8] ),
    .S(net88),
    .X(_10785_));
 sky130_fd_sc_hd__clkbuf_1 _25108_ (.A(_10785_),
    .X(_02612_));
 sky130_fd_sc_hd__mux2_1 _25109_ (.A0(_10727_),
    .A1(\datamem.data_ram[42][9] ),
    .S(_10784_),
    .X(_10786_));
 sky130_fd_sc_hd__clkbuf_1 _25110_ (.A(_10786_),
    .X(_02613_));
 sky130_fd_sc_hd__mux2_1 _25111_ (.A0(_10729_),
    .A1(\datamem.data_ram[42][10] ),
    .S(net88),
    .X(_10787_));
 sky130_fd_sc_hd__clkbuf_1 _25112_ (.A(_10787_),
    .X(_02614_));
 sky130_fd_sc_hd__mux2_1 _25113_ (.A0(_10731_),
    .A1(\datamem.data_ram[42][11] ),
    .S(net88),
    .X(_10788_));
 sky130_fd_sc_hd__clkbuf_1 _25114_ (.A(_10788_),
    .X(_02615_));
 sky130_fd_sc_hd__mux2_1 _25115_ (.A0(_10733_),
    .A1(\datamem.data_ram[42][12] ),
    .S(net88),
    .X(_10789_));
 sky130_fd_sc_hd__clkbuf_1 _25116_ (.A(_10789_),
    .X(_02616_));
 sky130_fd_sc_hd__mux2_1 _25117_ (.A0(_10735_),
    .A1(\datamem.data_ram[42][13] ),
    .S(net88),
    .X(_10790_));
 sky130_fd_sc_hd__clkbuf_1 _25118_ (.A(_10790_),
    .X(_02617_));
 sky130_fd_sc_hd__mux2_1 _25119_ (.A0(_10737_),
    .A1(\datamem.data_ram[42][14] ),
    .S(_10784_),
    .X(_10791_));
 sky130_fd_sc_hd__clkbuf_1 _25120_ (.A(_10791_),
    .X(_02618_));
 sky130_fd_sc_hd__mux2_1 _25121_ (.A0(_10739_),
    .A1(\datamem.data_ram[42][15] ),
    .S(_10784_),
    .X(_10792_));
 sky130_fd_sc_hd__clkbuf_1 _25122_ (.A(_10792_),
    .X(_02619_));
 sky130_fd_sc_hd__a21oi_2 _25123_ (.A1(_10520_),
    .A2(_10601_),
    .B1(_10705_),
    .Y(_10793_));
 sky130_fd_sc_hd__mux2_1 _25124_ (.A0(_10465_),
    .A1(\datamem.data_ram[42][24] ),
    .S(net87),
    .X(_10794_));
 sky130_fd_sc_hd__clkbuf_1 _25125_ (.A(_10794_),
    .X(_02620_));
 sky130_fd_sc_hd__mux2_1 _25126_ (.A0(_10468_),
    .A1(\datamem.data_ram[42][25] ),
    .S(net87),
    .X(_10795_));
 sky130_fd_sc_hd__clkbuf_1 _25127_ (.A(_10795_),
    .X(_02621_));
 sky130_fd_sc_hd__mux2_1 _25128_ (.A0(_10470_),
    .A1(\datamem.data_ram[42][26] ),
    .S(net87),
    .X(_10796_));
 sky130_fd_sc_hd__clkbuf_1 _25129_ (.A(_10796_),
    .X(_02622_));
 sky130_fd_sc_hd__mux2_1 _25130_ (.A0(_10472_),
    .A1(\datamem.data_ram[42][27] ),
    .S(net87),
    .X(_10797_));
 sky130_fd_sc_hd__clkbuf_1 _25131_ (.A(_10797_),
    .X(_02623_));
 sky130_fd_sc_hd__mux2_1 _25132_ (.A0(_10474_),
    .A1(\datamem.data_ram[42][28] ),
    .S(net87),
    .X(_10798_));
 sky130_fd_sc_hd__clkbuf_1 _25133_ (.A(_10798_),
    .X(_02624_));
 sky130_fd_sc_hd__mux2_1 _25134_ (.A0(_10476_),
    .A1(\datamem.data_ram[42][29] ),
    .S(net87),
    .X(_10799_));
 sky130_fd_sc_hd__clkbuf_1 _25135_ (.A(_10799_),
    .X(_02625_));
 sky130_fd_sc_hd__mux2_1 _25136_ (.A0(_10478_),
    .A1(\datamem.data_ram[42][30] ),
    .S(_10793_),
    .X(_10800_));
 sky130_fd_sc_hd__clkbuf_1 _25137_ (.A(_10800_),
    .X(_02626_));
 sky130_fd_sc_hd__mux2_1 _25138_ (.A0(_10480_),
    .A1(\datamem.data_ram[42][31] ),
    .S(_10793_),
    .X(_10801_));
 sky130_fd_sc_hd__clkbuf_1 _25139_ (.A(_10801_),
    .X(_02627_));
 sky130_fd_sc_hd__a21oi_4 _25140_ (.A1(_10570_),
    .A2(_10630_),
    .B1(_10705_),
    .Y(_10802_));
 sky130_fd_sc_hd__mux2_1 _25141_ (.A0(_10751_),
    .A1(\datamem.data_ram[41][16] ),
    .S(_10802_),
    .X(_10803_));
 sky130_fd_sc_hd__clkbuf_1 _25142_ (.A(_10803_),
    .X(_02628_));
 sky130_fd_sc_hd__mux2_1 _25143_ (.A0(_10754_),
    .A1(\datamem.data_ram[41][17] ),
    .S(_10802_),
    .X(_10804_));
 sky130_fd_sc_hd__clkbuf_1 _25144_ (.A(_10804_),
    .X(_02629_));
 sky130_fd_sc_hd__mux2_1 _25145_ (.A0(_10756_),
    .A1(\datamem.data_ram[41][18] ),
    .S(_10802_),
    .X(_10805_));
 sky130_fd_sc_hd__clkbuf_1 _25146_ (.A(_10805_),
    .X(_02630_));
 sky130_fd_sc_hd__mux2_1 _25147_ (.A0(_10758_),
    .A1(\datamem.data_ram[41][19] ),
    .S(_10802_),
    .X(_10806_));
 sky130_fd_sc_hd__clkbuf_1 _25148_ (.A(_10806_),
    .X(_02631_));
 sky130_fd_sc_hd__mux2_1 _25149_ (.A0(_10760_),
    .A1(\datamem.data_ram[41][20] ),
    .S(_10802_),
    .X(_10807_));
 sky130_fd_sc_hd__clkbuf_1 _25150_ (.A(_10807_),
    .X(_02632_));
 sky130_fd_sc_hd__mux2_1 _25151_ (.A0(_10762_),
    .A1(\datamem.data_ram[41][21] ),
    .S(_10802_),
    .X(_10808_));
 sky130_fd_sc_hd__clkbuf_1 _25152_ (.A(_10808_),
    .X(_02633_));
 sky130_fd_sc_hd__mux2_1 _25153_ (.A0(_10764_),
    .A1(\datamem.data_ram[41][22] ),
    .S(_10802_),
    .X(_10809_));
 sky130_fd_sc_hd__clkbuf_1 _25154_ (.A(_10809_),
    .X(_02634_));
 sky130_fd_sc_hd__mux2_1 _25155_ (.A0(_10766_),
    .A1(\datamem.data_ram[41][23] ),
    .S(_10802_),
    .X(_10810_));
 sky130_fd_sc_hd__clkbuf_1 _25156_ (.A(_10810_),
    .X(_02635_));
 sky130_fd_sc_hd__clkbuf_2 _25157_ (.A(_09297_),
    .X(_10811_));
 sky130_fd_sc_hd__a21oi_1 _25158_ (.A1(_10570_),
    .A2(_10601_),
    .B1(_10705_),
    .Y(_10812_));
 sky130_fd_sc_hd__mux2_1 _25159_ (.A0(_10811_),
    .A1(\datamem.data_ram[41][24] ),
    .S(net58),
    .X(_10813_));
 sky130_fd_sc_hd__clkbuf_1 _25160_ (.A(_10813_),
    .X(_02636_));
 sky130_fd_sc_hd__buf_2 _25161_ (.A(_09305_),
    .X(_10814_));
 sky130_fd_sc_hd__mux2_1 _25162_ (.A0(_10814_),
    .A1(\datamem.data_ram[41][25] ),
    .S(net58),
    .X(_10815_));
 sky130_fd_sc_hd__clkbuf_1 _25163_ (.A(_10815_),
    .X(_02637_));
 sky130_fd_sc_hd__buf_2 _25164_ (.A(_09309_),
    .X(_10816_));
 sky130_fd_sc_hd__mux2_1 _25165_ (.A0(_10816_),
    .A1(\datamem.data_ram[41][26] ),
    .S(net58),
    .X(_10817_));
 sky130_fd_sc_hd__clkbuf_1 _25166_ (.A(_10817_),
    .X(_02638_));
 sky130_fd_sc_hd__buf_2 _25167_ (.A(_09313_),
    .X(_10818_));
 sky130_fd_sc_hd__mux2_1 _25168_ (.A0(_10818_),
    .A1(\datamem.data_ram[41][27] ),
    .S(net58),
    .X(_10819_));
 sky130_fd_sc_hd__clkbuf_1 _25169_ (.A(_10819_),
    .X(_02639_));
 sky130_fd_sc_hd__buf_2 _25170_ (.A(_09317_),
    .X(_10820_));
 sky130_fd_sc_hd__mux2_1 _25171_ (.A0(_10820_),
    .A1(\datamem.data_ram[41][28] ),
    .S(net58),
    .X(_10821_));
 sky130_fd_sc_hd__clkbuf_1 _25172_ (.A(_10821_),
    .X(_02640_));
 sky130_fd_sc_hd__clkbuf_2 _25173_ (.A(_09321_),
    .X(_10822_));
 sky130_fd_sc_hd__mux2_1 _25174_ (.A0(_10822_),
    .A1(\datamem.data_ram[41][29] ),
    .S(net58),
    .X(_10823_));
 sky130_fd_sc_hd__clkbuf_1 _25175_ (.A(_10823_),
    .X(_02641_));
 sky130_fd_sc_hd__buf_2 _25176_ (.A(_09325_),
    .X(_10824_));
 sky130_fd_sc_hd__mux2_1 _25177_ (.A0(_10824_),
    .A1(\datamem.data_ram[41][30] ),
    .S(_10812_),
    .X(_10825_));
 sky130_fd_sc_hd__clkbuf_1 _25178_ (.A(_10825_),
    .X(_02642_));
 sky130_fd_sc_hd__clkbuf_2 _25179_ (.A(_09329_),
    .X(_10826_));
 sky130_fd_sc_hd__mux2_1 _25180_ (.A0(_10826_),
    .A1(\datamem.data_ram[41][31] ),
    .S(net58),
    .X(_10827_));
 sky130_fd_sc_hd__clkbuf_1 _25181_ (.A(_10827_),
    .X(_02643_));
 sky130_fd_sc_hd__buf_8 _25182_ (.A(_10500_),
    .X(_10828_));
 sky130_fd_sc_hd__a21oi_4 _25183_ (.A1(_10570_),
    .A2(_10640_),
    .B1(_10828_),
    .Y(_10829_));
 sky130_fd_sc_hd__mux2_1 _25184_ (.A0(_10724_),
    .A1(\datamem.data_ram[41][8] ),
    .S(net57),
    .X(_10830_));
 sky130_fd_sc_hd__clkbuf_1 _25185_ (.A(_10830_),
    .X(_02644_));
 sky130_fd_sc_hd__mux2_1 _25186_ (.A0(_10727_),
    .A1(\datamem.data_ram[41][9] ),
    .S(_10829_),
    .X(_10831_));
 sky130_fd_sc_hd__clkbuf_1 _25187_ (.A(_10831_),
    .X(_02645_));
 sky130_fd_sc_hd__mux2_1 _25188_ (.A0(_10729_),
    .A1(\datamem.data_ram[41][10] ),
    .S(net57),
    .X(_10832_));
 sky130_fd_sc_hd__clkbuf_1 _25189_ (.A(_10832_),
    .X(_02646_));
 sky130_fd_sc_hd__mux2_1 _25190_ (.A0(_10731_),
    .A1(\datamem.data_ram[41][11] ),
    .S(net57),
    .X(_10833_));
 sky130_fd_sc_hd__clkbuf_1 _25191_ (.A(_10833_),
    .X(_02647_));
 sky130_fd_sc_hd__mux2_1 _25192_ (.A0(_10733_),
    .A1(\datamem.data_ram[41][12] ),
    .S(net57),
    .X(_10834_));
 sky130_fd_sc_hd__clkbuf_1 _25193_ (.A(_10834_),
    .X(_02648_));
 sky130_fd_sc_hd__mux2_1 _25194_ (.A0(_10735_),
    .A1(\datamem.data_ram[41][13] ),
    .S(net57),
    .X(_10835_));
 sky130_fd_sc_hd__clkbuf_1 _25195_ (.A(_10835_),
    .X(_02649_));
 sky130_fd_sc_hd__mux2_1 _25196_ (.A0(_10737_),
    .A1(\datamem.data_ram[41][14] ),
    .S(_10829_),
    .X(_10836_));
 sky130_fd_sc_hd__clkbuf_1 _25197_ (.A(_10836_),
    .X(_02650_));
 sky130_fd_sc_hd__mux2_1 _25198_ (.A0(_10739_),
    .A1(\datamem.data_ram[41][15] ),
    .S(_10829_),
    .X(_10837_));
 sky130_fd_sc_hd__clkbuf_1 _25199_ (.A(_10837_),
    .X(_02651_));
 sky130_fd_sc_hd__buf_8 _25200_ (.A(_07122_),
    .X(_10838_));
 sky130_fd_sc_hd__a21oi_1 _25201_ (.A1(_10838_),
    .A2(_10601_),
    .B1(_10828_),
    .Y(_10839_));
 sky130_fd_sc_hd__mux2_1 _25202_ (.A0(_10811_),
    .A1(\datamem.data_ram[40][24] ),
    .S(net56),
    .X(_10840_));
 sky130_fd_sc_hd__clkbuf_1 _25203_ (.A(_10840_),
    .X(_02652_));
 sky130_fd_sc_hd__mux2_1 _25204_ (.A0(_10814_),
    .A1(\datamem.data_ram[40][25] ),
    .S(net56),
    .X(_10841_));
 sky130_fd_sc_hd__clkbuf_1 _25205_ (.A(_10841_),
    .X(_02653_));
 sky130_fd_sc_hd__mux2_1 _25206_ (.A0(_10816_),
    .A1(\datamem.data_ram[40][26] ),
    .S(net56),
    .X(_10842_));
 sky130_fd_sc_hd__clkbuf_1 _25207_ (.A(_10842_),
    .X(_02654_));
 sky130_fd_sc_hd__mux2_1 _25208_ (.A0(_10818_),
    .A1(\datamem.data_ram[40][27] ),
    .S(net56),
    .X(_10843_));
 sky130_fd_sc_hd__clkbuf_1 _25209_ (.A(_10843_),
    .X(_02655_));
 sky130_fd_sc_hd__mux2_1 _25210_ (.A0(_10820_),
    .A1(\datamem.data_ram[40][28] ),
    .S(net56),
    .X(_10844_));
 sky130_fd_sc_hd__clkbuf_1 _25211_ (.A(_10844_),
    .X(_02656_));
 sky130_fd_sc_hd__mux2_1 _25212_ (.A0(_10822_),
    .A1(\datamem.data_ram[40][29] ),
    .S(net56),
    .X(_10845_));
 sky130_fd_sc_hd__clkbuf_1 _25213_ (.A(_10845_),
    .X(_02657_));
 sky130_fd_sc_hd__mux2_1 _25214_ (.A0(_10824_),
    .A1(\datamem.data_ram[40][30] ),
    .S(_10839_),
    .X(_10846_));
 sky130_fd_sc_hd__clkbuf_1 _25215_ (.A(_10846_),
    .X(_02658_));
 sky130_fd_sc_hd__mux2_1 _25216_ (.A0(_10826_),
    .A1(\datamem.data_ram[40][31] ),
    .S(net56),
    .X(_10847_));
 sky130_fd_sc_hd__clkbuf_1 _25217_ (.A(_10847_),
    .X(_02659_));
 sky130_fd_sc_hd__a21oi_4 _25218_ (.A1(_10838_),
    .A2(_10630_),
    .B1(_10828_),
    .Y(_10848_));
 sky130_fd_sc_hd__mux2_1 _25219_ (.A0(_10751_),
    .A1(\datamem.data_ram[40][16] ),
    .S(_10848_),
    .X(_10849_));
 sky130_fd_sc_hd__clkbuf_1 _25220_ (.A(_10849_),
    .X(_02660_));
 sky130_fd_sc_hd__mux2_1 _25221_ (.A0(_10754_),
    .A1(\datamem.data_ram[40][17] ),
    .S(_10848_),
    .X(_10850_));
 sky130_fd_sc_hd__clkbuf_1 _25222_ (.A(_10850_),
    .X(_02661_));
 sky130_fd_sc_hd__mux2_1 _25223_ (.A0(_10756_),
    .A1(\datamem.data_ram[40][18] ),
    .S(_10848_),
    .X(_10851_));
 sky130_fd_sc_hd__clkbuf_1 _25224_ (.A(_10851_),
    .X(_02662_));
 sky130_fd_sc_hd__mux2_1 _25225_ (.A0(_10758_),
    .A1(\datamem.data_ram[40][19] ),
    .S(_10848_),
    .X(_10852_));
 sky130_fd_sc_hd__clkbuf_1 _25226_ (.A(_10852_),
    .X(_02663_));
 sky130_fd_sc_hd__mux2_1 _25227_ (.A0(_10760_),
    .A1(\datamem.data_ram[40][20] ),
    .S(_10848_),
    .X(_10853_));
 sky130_fd_sc_hd__clkbuf_1 _25228_ (.A(_10853_),
    .X(_02664_));
 sky130_fd_sc_hd__mux2_1 _25229_ (.A0(_10762_),
    .A1(\datamem.data_ram[40][21] ),
    .S(_10848_),
    .X(_10854_));
 sky130_fd_sc_hd__clkbuf_1 _25230_ (.A(_10854_),
    .X(_02665_));
 sky130_fd_sc_hd__mux2_1 _25231_ (.A0(_10764_),
    .A1(\datamem.data_ram[40][22] ),
    .S(_10848_),
    .X(_10855_));
 sky130_fd_sc_hd__clkbuf_1 _25232_ (.A(_10855_),
    .X(_02666_));
 sky130_fd_sc_hd__mux2_1 _25233_ (.A0(_10766_),
    .A1(\datamem.data_ram[40][23] ),
    .S(_10848_),
    .X(_10856_));
 sky130_fd_sc_hd__clkbuf_1 _25234_ (.A(_10856_),
    .X(_02667_));
 sky130_fd_sc_hd__a21oi_4 _25235_ (.A1(_10838_),
    .A2(_10640_),
    .B1(_10828_),
    .Y(_10857_));
 sky130_fd_sc_hd__mux2_1 _25236_ (.A0(_10724_),
    .A1(\datamem.data_ram[40][8] ),
    .S(net55),
    .X(_10858_));
 sky130_fd_sc_hd__clkbuf_1 _25237_ (.A(_10858_),
    .X(_02668_));
 sky130_fd_sc_hd__mux2_1 _25238_ (.A0(_10727_),
    .A1(\datamem.data_ram[40][9] ),
    .S(_10857_),
    .X(_10859_));
 sky130_fd_sc_hd__clkbuf_1 _25239_ (.A(_10859_),
    .X(_02669_));
 sky130_fd_sc_hd__mux2_1 _25240_ (.A0(_10729_),
    .A1(\datamem.data_ram[40][10] ),
    .S(net55),
    .X(_10860_));
 sky130_fd_sc_hd__clkbuf_1 _25241_ (.A(_10860_),
    .X(_02670_));
 sky130_fd_sc_hd__mux2_1 _25242_ (.A0(_10731_),
    .A1(\datamem.data_ram[40][11] ),
    .S(net55),
    .X(_10861_));
 sky130_fd_sc_hd__clkbuf_1 _25243_ (.A(_10861_),
    .X(_02671_));
 sky130_fd_sc_hd__mux2_1 _25244_ (.A0(_10733_),
    .A1(\datamem.data_ram[40][12] ),
    .S(net55),
    .X(_10862_));
 sky130_fd_sc_hd__clkbuf_1 _25245_ (.A(_10862_),
    .X(_02672_));
 sky130_fd_sc_hd__mux2_1 _25246_ (.A0(_10735_),
    .A1(\datamem.data_ram[40][13] ),
    .S(net55),
    .X(_10863_));
 sky130_fd_sc_hd__clkbuf_1 _25247_ (.A(_10863_),
    .X(_02673_));
 sky130_fd_sc_hd__mux2_1 _25248_ (.A0(_10737_),
    .A1(\datamem.data_ram[40][14] ),
    .S(_10857_),
    .X(_10864_));
 sky130_fd_sc_hd__clkbuf_1 _25249_ (.A(_10864_),
    .X(_02674_));
 sky130_fd_sc_hd__mux2_1 _25250_ (.A0(_10739_),
    .A1(\datamem.data_ram[40][15] ),
    .S(_10857_),
    .X(_10865_));
 sky130_fd_sc_hd__clkbuf_1 _25251_ (.A(_10865_),
    .X(_02675_));
 sky130_fd_sc_hd__or3_1 _25252_ (.A(_07077_),
    .B(_10042_),
    .C(_10044_),
    .X(_10866_));
 sky130_fd_sc_hd__buf_2 _25253_ (.A(_10866_),
    .X(_10867_));
 sky130_fd_sc_hd__and3_2 _25254_ (.A(_10142_),
    .B(_10049_),
    .C(_10052_),
    .X(_10868_));
 sky130_fd_sc_hd__and2_1 _25255_ (.A(_10405_),
    .B(_10868_),
    .X(_10869_));
 sky130_fd_sc_hd__a31o_1 _25256_ (.A1(_10538_),
    .A2(\datamem.data_ram[3][0] ),
    .A3(_10867_),
    .B1(_10869_),
    .X(_02676_));
 sky130_fd_sc_hd__and2_1 _25257_ (.A(_10408_),
    .B(_10868_),
    .X(_10870_));
 sky130_fd_sc_hd__a31o_1 _25258_ (.A1(_10538_),
    .A2(\datamem.data_ram[3][1] ),
    .A3(_10867_),
    .B1(_10870_),
    .X(_02677_));
 sky130_fd_sc_hd__and2_1 _25259_ (.A(_10410_),
    .B(_10868_),
    .X(_10871_));
 sky130_fd_sc_hd__a31o_1 _25260_ (.A1(_10538_),
    .A2(\datamem.data_ram[3][2] ),
    .A3(_10867_),
    .B1(_10871_),
    .X(_02678_));
 sky130_fd_sc_hd__and2_1 _25261_ (.A(_10413_),
    .B(_10868_),
    .X(_10872_));
 sky130_fd_sc_hd__a31o_1 _25262_ (.A1(_10538_),
    .A2(\datamem.data_ram[3][3] ),
    .A3(_10867_),
    .B1(_10872_),
    .X(_02679_));
 sky130_fd_sc_hd__and2_1 _25263_ (.A(_10067_),
    .B(_10868_),
    .X(_10873_));
 sky130_fd_sc_hd__a31o_1 _25264_ (.A1(_10538_),
    .A2(\datamem.data_ram[3][4] ),
    .A3(_10867_),
    .B1(_10873_),
    .X(_02680_));
 sky130_fd_sc_hd__and2_1 _25265_ (.A(_10416_),
    .B(_10868_),
    .X(_10874_));
 sky130_fd_sc_hd__a31o_1 _25266_ (.A1(_10538_),
    .A2(\datamem.data_ram[3][5] ),
    .A3(_10867_),
    .B1(_10874_),
    .X(_02681_));
 sky130_fd_sc_hd__and2_1 _25267_ (.A(_10418_),
    .B(_10868_),
    .X(_10875_));
 sky130_fd_sc_hd__a31o_1 _25268_ (.A1(_10538_),
    .A2(\datamem.data_ram[3][6] ),
    .A3(_10867_),
    .B1(_10875_),
    .X(_02682_));
 sky130_fd_sc_hd__clkbuf_4 _25269_ (.A(_10055_),
    .X(_10876_));
 sky130_fd_sc_hd__and2_1 _25270_ (.A(_10076_),
    .B(_10868_),
    .X(_10877_));
 sky130_fd_sc_hd__a31o_1 _25271_ (.A1(_10876_),
    .A2(\datamem.data_ram[3][7] ),
    .A3(_10867_),
    .B1(_10877_),
    .X(_02683_));
 sky130_fd_sc_hd__a21oi_4 _25272_ (.A1(_10741_),
    .A2(_10092_),
    .B1(_10828_),
    .Y(_10878_));
 sky130_fd_sc_hd__mux2_1 _25273_ (.A0(_10724_),
    .A1(\datamem.data_ram[3][8] ),
    .S(_10878_),
    .X(_10879_));
 sky130_fd_sc_hd__clkbuf_1 _25274_ (.A(_10879_),
    .X(_02684_));
 sky130_fd_sc_hd__mux2_1 _25275_ (.A0(_10727_),
    .A1(\datamem.data_ram[3][9] ),
    .S(_10878_),
    .X(_10880_));
 sky130_fd_sc_hd__clkbuf_1 _25276_ (.A(_10880_),
    .X(_02685_));
 sky130_fd_sc_hd__mux2_1 _25277_ (.A0(_10729_),
    .A1(\datamem.data_ram[3][10] ),
    .S(_10878_),
    .X(_10881_));
 sky130_fd_sc_hd__clkbuf_1 _25278_ (.A(_10881_),
    .X(_02686_));
 sky130_fd_sc_hd__mux2_1 _25279_ (.A0(_10731_),
    .A1(\datamem.data_ram[3][11] ),
    .S(_10878_),
    .X(_10882_));
 sky130_fd_sc_hd__clkbuf_1 _25280_ (.A(_10882_),
    .X(_02687_));
 sky130_fd_sc_hd__mux2_1 _25281_ (.A0(_10733_),
    .A1(\datamem.data_ram[3][12] ),
    .S(_10878_),
    .X(_10883_));
 sky130_fd_sc_hd__clkbuf_1 _25282_ (.A(_10883_),
    .X(_02688_));
 sky130_fd_sc_hd__mux2_1 _25283_ (.A0(_10735_),
    .A1(\datamem.data_ram[3][13] ),
    .S(_10878_),
    .X(_10884_));
 sky130_fd_sc_hd__clkbuf_1 _25284_ (.A(_10884_),
    .X(_02689_));
 sky130_fd_sc_hd__mux2_1 _25285_ (.A0(_10737_),
    .A1(\datamem.data_ram[3][14] ),
    .S(_10878_),
    .X(_10885_));
 sky130_fd_sc_hd__clkbuf_1 _25286_ (.A(_10885_),
    .X(_02690_));
 sky130_fd_sc_hd__mux2_1 _25287_ (.A0(_10739_),
    .A1(\datamem.data_ram[3][15] ),
    .S(_10878_),
    .X(_10886_));
 sky130_fd_sc_hd__clkbuf_1 _25288_ (.A(_10886_),
    .X(_02691_));
 sky130_fd_sc_hd__a21oi_4 _25289_ (.A1(_10741_),
    .A2(_10114_),
    .B1(_10828_),
    .Y(_10887_));
 sky130_fd_sc_hd__mux2_1 _25290_ (.A0(_10751_),
    .A1(\datamem.data_ram[3][16] ),
    .S(_10887_),
    .X(_10888_));
 sky130_fd_sc_hd__clkbuf_1 _25291_ (.A(_10888_),
    .X(_02692_));
 sky130_fd_sc_hd__mux2_1 _25292_ (.A0(_10754_),
    .A1(\datamem.data_ram[3][17] ),
    .S(_10887_),
    .X(_10889_));
 sky130_fd_sc_hd__clkbuf_1 _25293_ (.A(_10889_),
    .X(_02693_));
 sky130_fd_sc_hd__mux2_1 _25294_ (.A0(_10756_),
    .A1(\datamem.data_ram[3][18] ),
    .S(_10887_),
    .X(_10890_));
 sky130_fd_sc_hd__clkbuf_1 _25295_ (.A(_10890_),
    .X(_02694_));
 sky130_fd_sc_hd__mux2_1 _25296_ (.A0(_10758_),
    .A1(\datamem.data_ram[3][19] ),
    .S(_10887_),
    .X(_10891_));
 sky130_fd_sc_hd__clkbuf_1 _25297_ (.A(_10891_),
    .X(_02695_));
 sky130_fd_sc_hd__mux2_1 _25298_ (.A0(_10760_),
    .A1(\datamem.data_ram[3][20] ),
    .S(_10887_),
    .X(_10892_));
 sky130_fd_sc_hd__clkbuf_1 _25299_ (.A(_10892_),
    .X(_02696_));
 sky130_fd_sc_hd__mux2_1 _25300_ (.A0(_10762_),
    .A1(\datamem.data_ram[3][21] ),
    .S(_10887_),
    .X(_10893_));
 sky130_fd_sc_hd__clkbuf_1 _25301_ (.A(_10893_),
    .X(_02697_));
 sky130_fd_sc_hd__mux2_1 _25302_ (.A0(_10764_),
    .A1(\datamem.data_ram[3][22] ),
    .S(_10887_),
    .X(_10894_));
 sky130_fd_sc_hd__clkbuf_1 _25303_ (.A(_10894_),
    .X(_02698_));
 sky130_fd_sc_hd__mux2_1 _25304_ (.A0(_10766_),
    .A1(\datamem.data_ram[3][23] ),
    .S(_10887_),
    .X(_10895_));
 sky130_fd_sc_hd__clkbuf_1 _25305_ (.A(_10895_),
    .X(_02699_));
 sky130_fd_sc_hd__or2_2 _25306_ (.A(_08124_),
    .B(_07903_),
    .X(_10896_));
 sky130_fd_sc_hd__clkbuf_8 _25307_ (.A(_10896_),
    .X(_10897_));
 sky130_fd_sc_hd__nor2_4 _25308_ (.A(_09300_),
    .B(_10897_),
    .Y(_10898_));
 sky130_fd_sc_hd__a21oi_4 _25309_ (.A1(_10598_),
    .A2(_10898_),
    .B1(_10828_),
    .Y(_10899_));
 sky130_fd_sc_hd__mux2_1 _25310_ (.A0(_10811_),
    .A1(\datamem.data_ram[39][24] ),
    .S(_10899_),
    .X(_10900_));
 sky130_fd_sc_hd__clkbuf_1 _25311_ (.A(_10900_),
    .X(_02700_));
 sky130_fd_sc_hd__mux2_1 _25312_ (.A0(_10814_),
    .A1(\datamem.data_ram[39][25] ),
    .S(_10899_),
    .X(_10901_));
 sky130_fd_sc_hd__clkbuf_1 _25313_ (.A(_10901_),
    .X(_02701_));
 sky130_fd_sc_hd__mux2_1 _25314_ (.A0(_10816_),
    .A1(\datamem.data_ram[39][26] ),
    .S(_10899_),
    .X(_10902_));
 sky130_fd_sc_hd__clkbuf_1 _25315_ (.A(_10902_),
    .X(_02702_));
 sky130_fd_sc_hd__mux2_1 _25316_ (.A0(_10818_),
    .A1(\datamem.data_ram[39][27] ),
    .S(_10899_),
    .X(_10903_));
 sky130_fd_sc_hd__clkbuf_1 _25317_ (.A(_10903_),
    .X(_02703_));
 sky130_fd_sc_hd__mux2_1 _25318_ (.A0(_10820_),
    .A1(\datamem.data_ram[39][28] ),
    .S(_10899_),
    .X(_10904_));
 sky130_fd_sc_hd__clkbuf_1 _25319_ (.A(_10904_),
    .X(_02704_));
 sky130_fd_sc_hd__mux2_1 _25320_ (.A0(_10822_),
    .A1(\datamem.data_ram[39][29] ),
    .S(_10899_),
    .X(_10905_));
 sky130_fd_sc_hd__clkbuf_1 _25321_ (.A(_10905_),
    .X(_02705_));
 sky130_fd_sc_hd__mux2_1 _25322_ (.A0(_10824_),
    .A1(\datamem.data_ram[39][30] ),
    .S(_10899_),
    .X(_10906_));
 sky130_fd_sc_hd__clkbuf_1 _25323_ (.A(_10906_),
    .X(_02706_));
 sky130_fd_sc_hd__mux2_1 _25324_ (.A0(_10826_),
    .A1(\datamem.data_ram[39][31] ),
    .S(_10899_),
    .X(_10907_));
 sky130_fd_sc_hd__clkbuf_1 _25325_ (.A(_10907_),
    .X(_02707_));
 sky130_fd_sc_hd__nor2_8 _25326_ (.A(_09228_),
    .B(_10897_),
    .Y(_10908_));
 sky130_fd_sc_hd__a21oi_4 _25327_ (.A1(_10598_),
    .A2(_10908_),
    .B1(_10828_),
    .Y(_10909_));
 sky130_fd_sc_hd__mux2_1 _25328_ (.A0(_10751_),
    .A1(\datamem.data_ram[39][16] ),
    .S(_10909_),
    .X(_10910_));
 sky130_fd_sc_hd__clkbuf_1 _25329_ (.A(_10910_),
    .X(_02708_));
 sky130_fd_sc_hd__mux2_1 _25330_ (.A0(_10754_),
    .A1(\datamem.data_ram[39][17] ),
    .S(_10909_),
    .X(_10911_));
 sky130_fd_sc_hd__clkbuf_1 _25331_ (.A(_10911_),
    .X(_02709_));
 sky130_fd_sc_hd__mux2_1 _25332_ (.A0(_10756_),
    .A1(\datamem.data_ram[39][18] ),
    .S(_10909_),
    .X(_10912_));
 sky130_fd_sc_hd__clkbuf_1 _25333_ (.A(_10912_),
    .X(_02710_));
 sky130_fd_sc_hd__mux2_1 _25334_ (.A0(_10758_),
    .A1(\datamem.data_ram[39][19] ),
    .S(_10909_),
    .X(_10913_));
 sky130_fd_sc_hd__clkbuf_1 _25335_ (.A(_10913_),
    .X(_02711_));
 sky130_fd_sc_hd__mux2_1 _25336_ (.A0(_10760_),
    .A1(\datamem.data_ram[39][20] ),
    .S(_10909_),
    .X(_10914_));
 sky130_fd_sc_hd__clkbuf_1 _25337_ (.A(_10914_),
    .X(_02712_));
 sky130_fd_sc_hd__mux2_1 _25338_ (.A0(_10762_),
    .A1(\datamem.data_ram[39][21] ),
    .S(_10909_),
    .X(_10915_));
 sky130_fd_sc_hd__clkbuf_1 _25339_ (.A(_10915_),
    .X(_02713_));
 sky130_fd_sc_hd__mux2_1 _25340_ (.A0(_10764_),
    .A1(\datamem.data_ram[39][22] ),
    .S(_10909_),
    .X(_10916_));
 sky130_fd_sc_hd__clkbuf_1 _25341_ (.A(_10916_),
    .X(_02714_));
 sky130_fd_sc_hd__mux2_1 _25342_ (.A0(_10766_),
    .A1(\datamem.data_ram[39][23] ),
    .S(_10909_),
    .X(_10917_));
 sky130_fd_sc_hd__clkbuf_1 _25343_ (.A(_10917_),
    .X(_02715_));
 sky130_fd_sc_hd__buf_2 _25344_ (.A(_10043_),
    .X(_10918_));
 sky130_fd_sc_hd__or3_1 _25345_ (.A(_07791_),
    .B(_10918_),
    .C(_10897_),
    .X(_10919_));
 sky130_fd_sc_hd__buf_2 _25346_ (.A(_10919_),
    .X(_10920_));
 sky130_fd_sc_hd__buf_2 _25347_ (.A(_10051_),
    .X(_10921_));
 sky130_fd_sc_hd__nor2_2 _25348_ (.A(_08124_),
    .B(_07903_),
    .Y(_10922_));
 sky130_fd_sc_hd__and3_2 _25349_ (.A(_10325_),
    .B(_10921_),
    .C(_10922_),
    .X(_10923_));
 sky130_fd_sc_hd__and2_1 _25350_ (.A(_10405_),
    .B(_10923_),
    .X(_10924_));
 sky130_fd_sc_hd__a31o_1 _25351_ (.A1(_10876_),
    .A2(\datamem.data_ram[39][0] ),
    .A3(_10920_),
    .B1(_10924_),
    .X(_02716_));
 sky130_fd_sc_hd__and2_1 _25352_ (.A(_10408_),
    .B(_10923_),
    .X(_10925_));
 sky130_fd_sc_hd__a31o_1 _25353_ (.A1(_10876_),
    .A2(\datamem.data_ram[39][1] ),
    .A3(_10920_),
    .B1(_10925_),
    .X(_02717_));
 sky130_fd_sc_hd__and2_1 _25354_ (.A(_10410_),
    .B(_10923_),
    .X(_10926_));
 sky130_fd_sc_hd__a31o_1 _25355_ (.A1(_10876_),
    .A2(\datamem.data_ram[39][2] ),
    .A3(_10920_),
    .B1(_10926_),
    .X(_02718_));
 sky130_fd_sc_hd__and2_1 _25356_ (.A(_10413_),
    .B(_10923_),
    .X(_10927_));
 sky130_fd_sc_hd__a31o_1 _25357_ (.A1(_10876_),
    .A2(\datamem.data_ram[39][3] ),
    .A3(_10920_),
    .B1(_10927_),
    .X(_02719_));
 sky130_fd_sc_hd__and2_1 _25358_ (.A(_10067_),
    .B(_10923_),
    .X(_10928_));
 sky130_fd_sc_hd__a31o_1 _25359_ (.A1(_10876_),
    .A2(\datamem.data_ram[39][4] ),
    .A3(_10920_),
    .B1(_10928_),
    .X(_02720_));
 sky130_fd_sc_hd__and2_1 _25360_ (.A(_10416_),
    .B(_10923_),
    .X(_10929_));
 sky130_fd_sc_hd__a31o_1 _25361_ (.A1(_10876_),
    .A2(\datamem.data_ram[39][5] ),
    .A3(_10920_),
    .B1(_10929_),
    .X(_02721_));
 sky130_fd_sc_hd__and2_1 _25362_ (.A(_10418_),
    .B(_10923_),
    .X(_10930_));
 sky130_fd_sc_hd__a31o_1 _25363_ (.A1(_10876_),
    .A2(\datamem.data_ram[39][6] ),
    .A3(_10920_),
    .B1(_10930_),
    .X(_02722_));
 sky130_fd_sc_hd__and2_1 _25364_ (.A(_10076_),
    .B(_10923_),
    .X(_10931_));
 sky130_fd_sc_hd__a31o_1 _25365_ (.A1(_10876_),
    .A2(\datamem.data_ram[39][7] ),
    .A3(_10920_),
    .B1(_10931_),
    .X(_02723_));
 sky130_fd_sc_hd__clkbuf_8 _25366_ (.A(_08151_),
    .X(_10932_));
 sky130_fd_sc_hd__or3_1 _25367_ (.A(_07019_),
    .B(_10932_),
    .C(_10044_),
    .X(_10933_));
 sky130_fd_sc_hd__buf_2 _25368_ (.A(_10933_),
    .X(_10934_));
 sky130_fd_sc_hd__nor2_2 _25369_ (.A(_07131_),
    .B(_07154_),
    .Y(_10935_));
 sky130_fd_sc_hd__and3_2 _25370_ (.A(_09299_),
    .B(_10935_),
    .C(_10052_),
    .X(_10936_));
 sky130_fd_sc_hd__and2_1 _25371_ (.A(_10405_),
    .B(_10936_),
    .X(_10937_));
 sky130_fd_sc_hd__a31o_1 _25372_ (.A1(_10876_),
    .A2(\datamem.data_ram[13][0] ),
    .A3(_10934_),
    .B1(_10937_),
    .X(_02724_));
 sky130_fd_sc_hd__buf_2 _25373_ (.A(_10055_),
    .X(_10938_));
 sky130_fd_sc_hd__and2_1 _25374_ (.A(_10408_),
    .B(_10936_),
    .X(_10939_));
 sky130_fd_sc_hd__a31o_1 _25375_ (.A1(_10938_),
    .A2(\datamem.data_ram[13][1] ),
    .A3(_10934_),
    .B1(_10939_),
    .X(_02725_));
 sky130_fd_sc_hd__and2_1 _25376_ (.A(_10410_),
    .B(_10936_),
    .X(_10940_));
 sky130_fd_sc_hd__a31o_1 _25377_ (.A1(_10938_),
    .A2(\datamem.data_ram[13][2] ),
    .A3(_10934_),
    .B1(_10940_),
    .X(_02726_));
 sky130_fd_sc_hd__and2_1 _25378_ (.A(_10413_),
    .B(_10936_),
    .X(_10941_));
 sky130_fd_sc_hd__a31o_1 _25379_ (.A1(_10938_),
    .A2(\datamem.data_ram[13][3] ),
    .A3(_10934_),
    .B1(_10941_),
    .X(_02727_));
 sky130_fd_sc_hd__and2_1 _25380_ (.A(_10067_),
    .B(_10936_),
    .X(_10942_));
 sky130_fd_sc_hd__a31o_1 _25381_ (.A1(_10938_),
    .A2(\datamem.data_ram[13][4] ),
    .A3(_10934_),
    .B1(_10942_),
    .X(_02728_));
 sky130_fd_sc_hd__and2_1 _25382_ (.A(_10416_),
    .B(_10936_),
    .X(_10943_));
 sky130_fd_sc_hd__a31o_1 _25383_ (.A1(_10938_),
    .A2(\datamem.data_ram[13][5] ),
    .A3(_10934_),
    .B1(_10943_),
    .X(_02729_));
 sky130_fd_sc_hd__and2_1 _25384_ (.A(_10418_),
    .B(_10936_),
    .X(_10944_));
 sky130_fd_sc_hd__a31o_1 _25385_ (.A1(_10938_),
    .A2(\datamem.data_ram[13][6] ),
    .A3(_10934_),
    .B1(_10944_),
    .X(_02730_));
 sky130_fd_sc_hd__and2_1 _25386_ (.A(_10076_),
    .B(_10936_),
    .X(_10945_));
 sky130_fd_sc_hd__a31o_1 _25387_ (.A1(_10938_),
    .A2(\datamem.data_ram[13][7] ),
    .A3(_10934_),
    .B1(_10945_),
    .X(_02731_));
 sky130_fd_sc_hd__buf_2 _25388_ (.A(_08133_),
    .X(_10946_));
 sky130_fd_sc_hd__nand2_8 _25389_ (.A(_09225_),
    .B(_10051_),
    .Y(_10947_));
 sky130_fd_sc_hd__or2_1 _25390_ (.A(_10946_),
    .B(_10947_),
    .X(_10948_));
 sky130_fd_sc_hd__clkbuf_2 _25391_ (.A(_10948_),
    .X(_10949_));
 sky130_fd_sc_hd__nor2_1 _25392_ (.A(_10946_),
    .B(_10947_),
    .Y(_10950_));
 sky130_fd_sc_hd__and2_1 _25393_ (.A(_10405_),
    .B(_10950_),
    .X(_10951_));
 sky130_fd_sc_hd__a31o_1 _25394_ (.A1(_10938_),
    .A2(\datamem.data_ram[22][0] ),
    .A3(_10949_),
    .B1(_10951_),
    .X(_02732_));
 sky130_fd_sc_hd__and2_1 _25395_ (.A(_10408_),
    .B(_10950_),
    .X(_10952_));
 sky130_fd_sc_hd__a31o_1 _25396_ (.A1(_10938_),
    .A2(\datamem.data_ram[22][1] ),
    .A3(_10949_),
    .B1(_10952_),
    .X(_02733_));
 sky130_fd_sc_hd__and2_1 _25397_ (.A(_10410_),
    .B(_10950_),
    .X(_10953_));
 sky130_fd_sc_hd__a31o_1 _25398_ (.A1(_10938_),
    .A2(\datamem.data_ram[22][2] ),
    .A3(_10949_),
    .B1(_10953_),
    .X(_02734_));
 sky130_fd_sc_hd__buf_2 _25399_ (.A(_10055_),
    .X(_10954_));
 sky130_fd_sc_hd__and2_1 _25400_ (.A(_10413_),
    .B(_10950_),
    .X(_10955_));
 sky130_fd_sc_hd__a31o_1 _25401_ (.A1(_10954_),
    .A2(\datamem.data_ram[22][3] ),
    .A3(_10949_),
    .B1(_10955_),
    .X(_02735_));
 sky130_fd_sc_hd__and2_1 _25402_ (.A(_10067_),
    .B(_10950_),
    .X(_10956_));
 sky130_fd_sc_hd__a31o_1 _25403_ (.A1(_10954_),
    .A2(\datamem.data_ram[22][4] ),
    .A3(_10949_),
    .B1(_10956_),
    .X(_02736_));
 sky130_fd_sc_hd__and2_1 _25404_ (.A(_10416_),
    .B(_10950_),
    .X(_10957_));
 sky130_fd_sc_hd__a31o_1 _25405_ (.A1(_10954_),
    .A2(\datamem.data_ram[22][5] ),
    .A3(_10949_),
    .B1(_10957_),
    .X(_02737_));
 sky130_fd_sc_hd__and2_1 _25406_ (.A(_10418_),
    .B(_10950_),
    .X(_10958_));
 sky130_fd_sc_hd__a31o_1 _25407_ (.A1(_10954_),
    .A2(\datamem.data_ram[22][6] ),
    .A3(_10949_),
    .B1(_10958_),
    .X(_02738_));
 sky130_fd_sc_hd__and2_1 _25408_ (.A(_10076_),
    .B(_10950_),
    .X(_10959_));
 sky130_fd_sc_hd__a31o_1 _25409_ (.A1(_10954_),
    .A2(\datamem.data_ram[22][7] ),
    .A3(_10949_),
    .B1(_10959_),
    .X(_02739_));
 sky130_fd_sc_hd__nor2_8 _25410_ (.A(_10932_),
    .B(net104),
    .Y(_10960_));
 sky130_fd_sc_hd__a21oi_4 _25411_ (.A1(_10741_),
    .A2(_10960_),
    .B1(_10828_),
    .Y(_10961_));
 sky130_fd_sc_hd__mux2_1 _25412_ (.A0(_10751_),
    .A1(\datamem.data_ram[11][16] ),
    .S(_10961_),
    .X(_10962_));
 sky130_fd_sc_hd__clkbuf_1 _25413_ (.A(_10962_),
    .X(_02740_));
 sky130_fd_sc_hd__mux2_1 _25414_ (.A0(_10754_),
    .A1(\datamem.data_ram[11][17] ),
    .S(_10961_),
    .X(_10963_));
 sky130_fd_sc_hd__clkbuf_1 _25415_ (.A(_10963_),
    .X(_02741_));
 sky130_fd_sc_hd__mux2_1 _25416_ (.A0(_10756_),
    .A1(\datamem.data_ram[11][18] ),
    .S(_10961_),
    .X(_10964_));
 sky130_fd_sc_hd__clkbuf_1 _25417_ (.A(_10964_),
    .X(_02742_));
 sky130_fd_sc_hd__mux2_1 _25418_ (.A0(_10758_),
    .A1(\datamem.data_ram[11][19] ),
    .S(_10961_),
    .X(_10965_));
 sky130_fd_sc_hd__clkbuf_1 _25419_ (.A(_10965_),
    .X(_02743_));
 sky130_fd_sc_hd__mux2_1 _25420_ (.A0(_10760_),
    .A1(\datamem.data_ram[11][20] ),
    .S(_10961_),
    .X(_10966_));
 sky130_fd_sc_hd__clkbuf_1 _25421_ (.A(_10966_),
    .X(_02744_));
 sky130_fd_sc_hd__mux2_1 _25422_ (.A0(_10762_),
    .A1(\datamem.data_ram[11][21] ),
    .S(_10961_),
    .X(_10967_));
 sky130_fd_sc_hd__clkbuf_1 _25423_ (.A(_10967_),
    .X(_02745_));
 sky130_fd_sc_hd__mux2_1 _25424_ (.A0(_10764_),
    .A1(\datamem.data_ram[11][22] ),
    .S(_10961_),
    .X(_10968_));
 sky130_fd_sc_hd__clkbuf_1 _25425_ (.A(_10968_),
    .X(_02746_));
 sky130_fd_sc_hd__mux2_1 _25426_ (.A0(_10766_),
    .A1(\datamem.data_ram[11][23] ),
    .S(_10961_),
    .X(_10969_));
 sky130_fd_sc_hd__clkbuf_1 _25427_ (.A(_10969_),
    .X(_02747_));
 sky130_fd_sc_hd__a21oi_4 _25428_ (.A1(_10520_),
    .A2(_10630_),
    .B1(_10828_),
    .Y(_10970_));
 sky130_fd_sc_hd__mux2_1 _25429_ (.A0(_10751_),
    .A1(\datamem.data_ram[42][16] ),
    .S(_10970_),
    .X(_10971_));
 sky130_fd_sc_hd__clkbuf_1 _25430_ (.A(_10971_),
    .X(_02748_));
 sky130_fd_sc_hd__mux2_1 _25431_ (.A0(_10754_),
    .A1(\datamem.data_ram[42][17] ),
    .S(_10970_),
    .X(_10972_));
 sky130_fd_sc_hd__clkbuf_1 _25432_ (.A(_10972_),
    .X(_02749_));
 sky130_fd_sc_hd__mux2_1 _25433_ (.A0(_10756_),
    .A1(\datamem.data_ram[42][18] ),
    .S(_10970_),
    .X(_10973_));
 sky130_fd_sc_hd__clkbuf_1 _25434_ (.A(_10973_),
    .X(_02750_));
 sky130_fd_sc_hd__mux2_1 _25435_ (.A0(_10758_),
    .A1(\datamem.data_ram[42][19] ),
    .S(_10970_),
    .X(_10974_));
 sky130_fd_sc_hd__clkbuf_1 _25436_ (.A(_10974_),
    .X(_02751_));
 sky130_fd_sc_hd__mux2_1 _25437_ (.A0(_10760_),
    .A1(\datamem.data_ram[42][20] ),
    .S(_10970_),
    .X(_10975_));
 sky130_fd_sc_hd__clkbuf_1 _25438_ (.A(_10975_),
    .X(_02752_));
 sky130_fd_sc_hd__mux2_1 _25439_ (.A0(_10762_),
    .A1(\datamem.data_ram[42][21] ),
    .S(_10970_),
    .X(_10976_));
 sky130_fd_sc_hd__clkbuf_1 _25440_ (.A(_10976_),
    .X(_02753_));
 sky130_fd_sc_hd__mux2_1 _25441_ (.A0(_10764_),
    .A1(\datamem.data_ram[42][22] ),
    .S(_10970_),
    .X(_10977_));
 sky130_fd_sc_hd__clkbuf_1 _25442_ (.A(_10977_),
    .X(_02754_));
 sky130_fd_sc_hd__mux2_1 _25443_ (.A0(_10766_),
    .A1(\datamem.data_ram[42][23] ),
    .S(_10970_),
    .X(_10978_));
 sky130_fd_sc_hd__clkbuf_1 _25444_ (.A(_10978_),
    .X(_02755_));
 sky130_fd_sc_hd__clkbuf_16 _25445_ (.A(_07122_),
    .X(_10979_));
 sky130_fd_sc_hd__nand2_4 _25446_ (.A(_10979_),
    .B(_10051_),
    .Y(_10980_));
 sky130_fd_sc_hd__nor2_4 _25447_ (.A(_10600_),
    .B(_10980_),
    .Y(_10981_));
 sky130_fd_sc_hd__nor2_2 _25448_ (.A(_10780_),
    .B(_10981_),
    .Y(_10982_));
 sky130_fd_sc_hd__a22o_1 _25449_ (.A1(_10048_),
    .A2(_10981_),
    .B1(_10982_),
    .B2(\datamem.data_ram[40][0] ),
    .X(_02756_));
 sky130_fd_sc_hd__a22o_1 _25450_ (.A1(_10058_),
    .A2(_10981_),
    .B1(_10982_),
    .B2(\datamem.data_ram[40][1] ),
    .X(_02757_));
 sky130_fd_sc_hd__a22o_1 _25451_ (.A1(_10061_),
    .A2(_10981_),
    .B1(_10982_),
    .B2(\datamem.data_ram[40][2] ),
    .X(_02758_));
 sky130_fd_sc_hd__a22o_1 _25452_ (.A1(_10064_),
    .A2(_10981_),
    .B1(_10982_),
    .B2(\datamem.data_ram[40][3] ),
    .X(_02759_));
 sky130_fd_sc_hd__a22o_1 _25453_ (.A1(_10782_),
    .A2(_10981_),
    .B1(_10982_),
    .B2(\datamem.data_ram[40][4] ),
    .X(_02760_));
 sky130_fd_sc_hd__a22o_1 _25454_ (.A1(_10070_),
    .A2(_10981_),
    .B1(_10982_),
    .B2(\datamem.data_ram[40][5] ),
    .X(_02761_));
 sky130_fd_sc_hd__a22o_1 _25455_ (.A1(_10073_),
    .A2(_10981_),
    .B1(_10982_),
    .B2(\datamem.data_ram[40][6] ),
    .X(_02762_));
 sky130_fd_sc_hd__a22o_1 _25456_ (.A1(_10783_),
    .A2(_10981_),
    .B1(_10982_),
    .B2(\datamem.data_ram[40][7] ),
    .X(_02763_));
 sky130_fd_sc_hd__or3_1 _25457_ (.A(_07182_),
    .B(_10932_),
    .C(_10044_),
    .X(_10983_));
 sky130_fd_sc_hd__clkbuf_2 _25458_ (.A(_10983_),
    .X(_10984_));
 sky130_fd_sc_hd__and3_2 _25459_ (.A(_09351_),
    .B(_10935_),
    .C(_10052_),
    .X(_10985_));
 sky130_fd_sc_hd__and2_1 _25460_ (.A(_10405_),
    .B(_10985_),
    .X(_10986_));
 sky130_fd_sc_hd__a31o_1 _25461_ (.A1(_10954_),
    .A2(\datamem.data_ram[12][0] ),
    .A3(_10984_),
    .B1(_10986_),
    .X(_02764_));
 sky130_fd_sc_hd__and2_1 _25462_ (.A(_10408_),
    .B(_10985_),
    .X(_10987_));
 sky130_fd_sc_hd__a31o_1 _25463_ (.A1(_10954_),
    .A2(\datamem.data_ram[12][1] ),
    .A3(_10984_),
    .B1(_10987_),
    .X(_02765_));
 sky130_fd_sc_hd__and2_1 _25464_ (.A(_10410_),
    .B(_10985_),
    .X(_10988_));
 sky130_fd_sc_hd__a31o_1 _25465_ (.A1(_10954_),
    .A2(\datamem.data_ram[12][2] ),
    .A3(_10984_),
    .B1(_10988_),
    .X(_02766_));
 sky130_fd_sc_hd__and2_1 _25466_ (.A(_10413_),
    .B(_10985_),
    .X(_10989_));
 sky130_fd_sc_hd__a31o_1 _25467_ (.A1(_10954_),
    .A2(\datamem.data_ram[12][3] ),
    .A3(_10984_),
    .B1(_10989_),
    .X(_02767_));
 sky130_fd_sc_hd__and2_1 _25468_ (.A(_10067_),
    .B(_10985_),
    .X(_10990_));
 sky130_fd_sc_hd__a31o_1 _25469_ (.A1(_10954_),
    .A2(\datamem.data_ram[12][4] ),
    .A3(_10984_),
    .B1(_10990_),
    .X(_02768_));
 sky130_fd_sc_hd__clkbuf_4 _25470_ (.A(_10055_),
    .X(_10991_));
 sky130_fd_sc_hd__and2_1 _25471_ (.A(_10416_),
    .B(_10985_),
    .X(_10992_));
 sky130_fd_sc_hd__a31o_1 _25472_ (.A1(_10991_),
    .A2(\datamem.data_ram[12][5] ),
    .A3(_10984_),
    .B1(_10992_),
    .X(_02769_));
 sky130_fd_sc_hd__and2_1 _25473_ (.A(_10418_),
    .B(_10985_),
    .X(_10993_));
 sky130_fd_sc_hd__a31o_1 _25474_ (.A1(_10991_),
    .A2(\datamem.data_ram[12][6] ),
    .A3(_10984_),
    .B1(_10993_),
    .X(_02770_));
 sky130_fd_sc_hd__and2_1 _25475_ (.A(_10076_),
    .B(_10985_),
    .X(_10994_));
 sky130_fd_sc_hd__a31o_1 _25476_ (.A1(_10991_),
    .A2(\datamem.data_ram[12][7] ),
    .A3(_10984_),
    .B1(_10994_),
    .X(_02771_));
 sky130_fd_sc_hd__nor3_1 _25477_ (.A(_07808_),
    .B(_10043_),
    .C(_10600_),
    .Y(_10995_));
 sky130_fd_sc_hd__nor2_2 _25478_ (.A(_10780_),
    .B(net35),
    .Y(_10996_));
 sky130_fd_sc_hd__a22o_1 _25479_ (.A1(_10048_),
    .A2(net35),
    .B1(_10996_),
    .B2(\datamem.data_ram[41][0] ),
    .X(_02772_));
 sky130_fd_sc_hd__a22o_1 _25480_ (.A1(_10058_),
    .A2(net35),
    .B1(_10996_),
    .B2(\datamem.data_ram[41][1] ),
    .X(_02773_));
 sky130_fd_sc_hd__a22o_1 _25481_ (.A1(_10061_),
    .A2(net35),
    .B1(_10996_),
    .B2(\datamem.data_ram[41][2] ),
    .X(_02774_));
 sky130_fd_sc_hd__a22o_1 _25482_ (.A1(_10064_),
    .A2(net35),
    .B1(_10996_),
    .B2(\datamem.data_ram[41][3] ),
    .X(_02775_));
 sky130_fd_sc_hd__a22o_1 _25483_ (.A1(_10782_),
    .A2(net35),
    .B1(_10996_),
    .B2(\datamem.data_ram[41][4] ),
    .X(_02776_));
 sky130_fd_sc_hd__a22o_1 _25484_ (.A1(_10070_),
    .A2(net35),
    .B1(_10996_),
    .B2(\datamem.data_ram[41][5] ),
    .X(_02777_));
 sky130_fd_sc_hd__a22o_1 _25485_ (.A1(_10073_),
    .A2(_10995_),
    .B1(_10996_),
    .B2(\datamem.data_ram[41][6] ),
    .X(_02778_));
 sky130_fd_sc_hd__a22o_1 _25486_ (.A1(_10783_),
    .A2(net35),
    .B1(_10996_),
    .B2(\datamem.data_ram[41][7] ),
    .X(_02779_));
 sky130_fd_sc_hd__nor2_8 _25487_ (.A(_08151_),
    .B(net110),
    .Y(_10997_));
 sky130_fd_sc_hd__buf_8 _25488_ (.A(_10500_),
    .X(_10998_));
 sky130_fd_sc_hd__a21oi_4 _25489_ (.A1(_10570_),
    .A2(_10997_),
    .B1(_10998_),
    .Y(_10999_));
 sky130_fd_sc_hd__mux2_1 _25490_ (.A0(_10811_),
    .A1(\datamem.data_ram[9][24] ),
    .S(_10999_),
    .X(_11000_));
 sky130_fd_sc_hd__clkbuf_1 _25491_ (.A(_11000_),
    .X(_02780_));
 sky130_fd_sc_hd__mux2_1 _25492_ (.A0(_10814_),
    .A1(\datamem.data_ram[9][25] ),
    .S(_10999_),
    .X(_11001_));
 sky130_fd_sc_hd__clkbuf_1 _25493_ (.A(_11001_),
    .X(_02781_));
 sky130_fd_sc_hd__mux2_1 _25494_ (.A0(_10816_),
    .A1(\datamem.data_ram[9][26] ),
    .S(_10999_),
    .X(_11002_));
 sky130_fd_sc_hd__clkbuf_1 _25495_ (.A(_11002_),
    .X(_02782_));
 sky130_fd_sc_hd__mux2_1 _25496_ (.A0(_10818_),
    .A1(\datamem.data_ram[9][27] ),
    .S(_10999_),
    .X(_11003_));
 sky130_fd_sc_hd__clkbuf_1 _25497_ (.A(_11003_),
    .X(_02783_));
 sky130_fd_sc_hd__mux2_1 _25498_ (.A0(_10820_),
    .A1(\datamem.data_ram[9][28] ),
    .S(_10999_),
    .X(_11004_));
 sky130_fd_sc_hd__clkbuf_1 _25499_ (.A(_11004_),
    .X(_02784_));
 sky130_fd_sc_hd__mux2_1 _25500_ (.A0(_10822_),
    .A1(\datamem.data_ram[9][29] ),
    .S(_10999_),
    .X(_11005_));
 sky130_fd_sc_hd__clkbuf_1 _25501_ (.A(_11005_),
    .X(_02785_));
 sky130_fd_sc_hd__mux2_1 _25502_ (.A0(_10824_),
    .A1(\datamem.data_ram[9][30] ),
    .S(_10999_),
    .X(_11006_));
 sky130_fd_sc_hd__clkbuf_1 _25503_ (.A(_11006_),
    .X(_02786_));
 sky130_fd_sc_hd__mux2_1 _25504_ (.A0(_10826_),
    .A1(\datamem.data_ram[9][31] ),
    .S(_10999_),
    .X(_11007_));
 sky130_fd_sc_hd__clkbuf_1 _25505_ (.A(_11007_),
    .X(_02787_));
 sky130_fd_sc_hd__or3_1 _25506_ (.A(_07028_),
    .B(_10918_),
    .C(_10897_),
    .X(_11008_));
 sky130_fd_sc_hd__buf_2 _25507_ (.A(_11008_),
    .X(_11009_));
 sky130_fd_sc_hd__and3_2 _25508_ (.A(_09226_),
    .B(_10921_),
    .C(_10922_),
    .X(_11010_));
 sky130_fd_sc_hd__and2_1 _25509_ (.A(_10405_),
    .B(_11010_),
    .X(_11011_));
 sky130_fd_sc_hd__a31o_1 _25510_ (.A1(_10991_),
    .A2(\datamem.data_ram[38][0] ),
    .A3(_11009_),
    .B1(_11011_),
    .X(_02788_));
 sky130_fd_sc_hd__and2_1 _25511_ (.A(_10408_),
    .B(_11010_),
    .X(_11012_));
 sky130_fd_sc_hd__a31o_1 _25512_ (.A1(_10991_),
    .A2(\datamem.data_ram[38][1] ),
    .A3(_11009_),
    .B1(_11012_),
    .X(_02789_));
 sky130_fd_sc_hd__and2_1 _25513_ (.A(_10410_),
    .B(_11010_),
    .X(_11013_));
 sky130_fd_sc_hd__a31o_1 _25514_ (.A1(_10991_),
    .A2(\datamem.data_ram[38][2] ),
    .A3(_11009_),
    .B1(_11013_),
    .X(_02790_));
 sky130_fd_sc_hd__and2_1 _25515_ (.A(_10413_),
    .B(_11010_),
    .X(_11014_));
 sky130_fd_sc_hd__a31o_1 _25516_ (.A1(_10991_),
    .A2(\datamem.data_ram[38][3] ),
    .A3(_11009_),
    .B1(_11014_),
    .X(_02791_));
 sky130_fd_sc_hd__and2_1 _25517_ (.A(_10067_),
    .B(_11010_),
    .X(_11015_));
 sky130_fd_sc_hd__a31o_1 _25518_ (.A1(_10991_),
    .A2(\datamem.data_ram[38][4] ),
    .A3(_11009_),
    .B1(_11015_),
    .X(_02792_));
 sky130_fd_sc_hd__and2_1 _25519_ (.A(_10416_),
    .B(_11010_),
    .X(_11016_));
 sky130_fd_sc_hd__a31o_1 _25520_ (.A1(_10991_),
    .A2(\datamem.data_ram[38][5] ),
    .A3(_11009_),
    .B1(_11016_),
    .X(_02793_));
 sky130_fd_sc_hd__and2_1 _25521_ (.A(_10418_),
    .B(_11010_),
    .X(_11017_));
 sky130_fd_sc_hd__a31o_1 _25522_ (.A1(_10991_),
    .A2(\datamem.data_ram[38][6] ),
    .A3(_11009_),
    .B1(_11017_),
    .X(_02794_));
 sky130_fd_sc_hd__clkbuf_4 _25523_ (.A(_10055_),
    .X(_11018_));
 sky130_fd_sc_hd__and2_1 _25524_ (.A(_10076_),
    .B(_11010_),
    .X(_11019_));
 sky130_fd_sc_hd__a31o_1 _25525_ (.A1(_11018_),
    .A2(\datamem.data_ram[38][7] ),
    .A3(_11009_),
    .B1(_11019_),
    .X(_02795_));
 sky130_fd_sc_hd__nor2_4 _25526_ (.A(_08151_),
    .B(_09268_),
    .Y(_11020_));
 sky130_fd_sc_hd__a21oi_4 _25527_ (.A1(_10838_),
    .A2(_11020_),
    .B1(_10998_),
    .Y(_11021_));
 sky130_fd_sc_hd__mux2_1 _25528_ (.A0(_10724_),
    .A1(\datamem.data_ram[8][8] ),
    .S(net54),
    .X(_11022_));
 sky130_fd_sc_hd__clkbuf_1 _25529_ (.A(_11022_),
    .X(_02796_));
 sky130_fd_sc_hd__mux2_1 _25530_ (.A0(_10727_),
    .A1(\datamem.data_ram[8][9] ),
    .S(net54),
    .X(_11023_));
 sky130_fd_sc_hd__clkbuf_1 _25531_ (.A(_11023_),
    .X(_02797_));
 sky130_fd_sc_hd__mux2_1 _25532_ (.A0(_10729_),
    .A1(\datamem.data_ram[8][10] ),
    .S(net54),
    .X(_11024_));
 sky130_fd_sc_hd__clkbuf_1 _25533_ (.A(_11024_),
    .X(_02798_));
 sky130_fd_sc_hd__mux2_1 _25534_ (.A0(_10731_),
    .A1(\datamem.data_ram[8][11] ),
    .S(net54),
    .X(_11025_));
 sky130_fd_sc_hd__clkbuf_1 _25535_ (.A(_11025_),
    .X(_02799_));
 sky130_fd_sc_hd__mux2_1 _25536_ (.A0(_10733_),
    .A1(\datamem.data_ram[8][12] ),
    .S(net54),
    .X(_11026_));
 sky130_fd_sc_hd__clkbuf_1 _25537_ (.A(_11026_),
    .X(_02800_));
 sky130_fd_sc_hd__mux2_1 _25538_ (.A0(_10735_),
    .A1(\datamem.data_ram[8][13] ),
    .S(_11021_),
    .X(_11027_));
 sky130_fd_sc_hd__clkbuf_1 _25539_ (.A(_11027_),
    .X(_02801_));
 sky130_fd_sc_hd__mux2_1 _25540_ (.A0(_10737_),
    .A1(\datamem.data_ram[8][14] ),
    .S(_11021_),
    .X(_11028_));
 sky130_fd_sc_hd__clkbuf_1 _25541_ (.A(_11028_),
    .X(_02802_));
 sky130_fd_sc_hd__mux2_1 _25542_ (.A0(_10739_),
    .A1(\datamem.data_ram[8][15] ),
    .S(_11021_),
    .X(_11029_));
 sky130_fd_sc_hd__clkbuf_1 _25543_ (.A(_11029_),
    .X(_02803_));
 sky130_fd_sc_hd__a21oi_4 _25544_ (.A1(_10570_),
    .A2(_10960_),
    .B1(_10998_),
    .Y(_11030_));
 sky130_fd_sc_hd__mux2_1 _25545_ (.A0(_10751_),
    .A1(\datamem.data_ram[9][16] ),
    .S(_11030_),
    .X(_11031_));
 sky130_fd_sc_hd__clkbuf_1 _25546_ (.A(_11031_),
    .X(_02804_));
 sky130_fd_sc_hd__mux2_1 _25547_ (.A0(_10754_),
    .A1(\datamem.data_ram[9][17] ),
    .S(_11030_),
    .X(_11032_));
 sky130_fd_sc_hd__clkbuf_1 _25548_ (.A(_11032_),
    .X(_02805_));
 sky130_fd_sc_hd__mux2_1 _25549_ (.A0(_10756_),
    .A1(\datamem.data_ram[9][18] ),
    .S(_11030_),
    .X(_11033_));
 sky130_fd_sc_hd__clkbuf_1 _25550_ (.A(_11033_),
    .X(_02806_));
 sky130_fd_sc_hd__mux2_1 _25551_ (.A0(_10758_),
    .A1(\datamem.data_ram[9][19] ),
    .S(_11030_),
    .X(_11034_));
 sky130_fd_sc_hd__clkbuf_1 _25552_ (.A(_11034_),
    .X(_02807_));
 sky130_fd_sc_hd__mux2_1 _25553_ (.A0(_10760_),
    .A1(\datamem.data_ram[9][20] ),
    .S(_11030_),
    .X(_11035_));
 sky130_fd_sc_hd__clkbuf_1 _25554_ (.A(_11035_),
    .X(_02808_));
 sky130_fd_sc_hd__mux2_1 _25555_ (.A0(_10762_),
    .A1(\datamem.data_ram[9][21] ),
    .S(_11030_),
    .X(_11036_));
 sky130_fd_sc_hd__clkbuf_1 _25556_ (.A(_11036_),
    .X(_02809_));
 sky130_fd_sc_hd__mux2_1 _25557_ (.A0(_10764_),
    .A1(\datamem.data_ram[9][22] ),
    .S(_11030_),
    .X(_11037_));
 sky130_fd_sc_hd__clkbuf_1 _25558_ (.A(_11037_),
    .X(_02810_));
 sky130_fd_sc_hd__mux2_1 _25559_ (.A0(_10766_),
    .A1(\datamem.data_ram[9][23] ),
    .S(_11030_),
    .X(_11038_));
 sky130_fd_sc_hd__clkbuf_1 _25560_ (.A(_11038_),
    .X(_02811_));
 sky130_fd_sc_hd__nand2_4 _25561_ (.A(_09350_),
    .B(_10051_),
    .Y(_11039_));
 sky130_fd_sc_hd__or2_1 _25562_ (.A(_10946_),
    .B(_11039_),
    .X(_11040_));
 sky130_fd_sc_hd__buf_2 _25563_ (.A(_11040_),
    .X(_11041_));
 sky130_fd_sc_hd__nor2_2 _25564_ (.A(_10946_),
    .B(_11039_),
    .Y(_11042_));
 sky130_fd_sc_hd__and2_1 _25565_ (.A(_10405_),
    .B(_11042_),
    .X(_11043_));
 sky130_fd_sc_hd__a31o_1 _25566_ (.A1(_11018_),
    .A2(\datamem.data_ram[20][0] ),
    .A3(_11041_),
    .B1(_11043_),
    .X(_02812_));
 sky130_fd_sc_hd__and2_1 _25567_ (.A(_10408_),
    .B(_11042_),
    .X(_11044_));
 sky130_fd_sc_hd__a31o_1 _25568_ (.A1(_11018_),
    .A2(\datamem.data_ram[20][1] ),
    .A3(_11041_),
    .B1(_11044_),
    .X(_02813_));
 sky130_fd_sc_hd__and2_1 _25569_ (.A(_10410_),
    .B(_11042_),
    .X(_11045_));
 sky130_fd_sc_hd__a31o_1 _25570_ (.A1(_11018_),
    .A2(\datamem.data_ram[20][2] ),
    .A3(_11041_),
    .B1(_11045_),
    .X(_02814_));
 sky130_fd_sc_hd__and2_1 _25571_ (.A(_10413_),
    .B(_11042_),
    .X(_11046_));
 sky130_fd_sc_hd__a31o_1 _25572_ (.A1(_11018_),
    .A2(\datamem.data_ram[20][3] ),
    .A3(_11041_),
    .B1(_11046_),
    .X(_02815_));
 sky130_fd_sc_hd__clkbuf_4 _25573_ (.A(_10066_),
    .X(_11047_));
 sky130_fd_sc_hd__and2_1 _25574_ (.A(_11047_),
    .B(_11042_),
    .X(_11048_));
 sky130_fd_sc_hd__a31o_1 _25575_ (.A1(_11018_),
    .A2(\datamem.data_ram[20][4] ),
    .A3(_11041_),
    .B1(_11048_),
    .X(_02816_));
 sky130_fd_sc_hd__and2_1 _25576_ (.A(_10416_),
    .B(_11042_),
    .X(_11049_));
 sky130_fd_sc_hd__a31o_1 _25577_ (.A1(_11018_),
    .A2(\datamem.data_ram[20][5] ),
    .A3(_11041_),
    .B1(_11049_),
    .X(_02817_));
 sky130_fd_sc_hd__and2_1 _25578_ (.A(_10418_),
    .B(_11042_),
    .X(_11050_));
 sky130_fd_sc_hd__a31o_1 _25579_ (.A1(_11018_),
    .A2(\datamem.data_ram[20][6] ),
    .A3(_11041_),
    .B1(_11050_),
    .X(_02818_));
 sky130_fd_sc_hd__and2_1 _25580_ (.A(_10076_),
    .B(_11042_),
    .X(_11051_));
 sky130_fd_sc_hd__a31o_1 _25581_ (.A1(_11018_),
    .A2(\datamem.data_ram[20][7] ),
    .A3(_11041_),
    .B1(_11051_),
    .X(_02819_));
 sky130_fd_sc_hd__or3_1 _25582_ (.A(_07019_),
    .B(_10946_),
    .C(_10044_),
    .X(_11052_));
 sky130_fd_sc_hd__buf_2 _25583_ (.A(_11052_),
    .X(_11053_));
 sky130_fd_sc_hd__nor2_1 _25584_ (.A(_08124_),
    .B(_07177_),
    .Y(_11054_));
 sky130_fd_sc_hd__and3_2 _25585_ (.A(_09299_),
    .B(_11054_),
    .C(_10052_),
    .X(_11055_));
 sky130_fd_sc_hd__and2_1 _25586_ (.A(_10405_),
    .B(_11055_),
    .X(_11056_));
 sky130_fd_sc_hd__a31o_1 _25587_ (.A1(_11018_),
    .A2(\datamem.data_ram[21][0] ),
    .A3(_11053_),
    .B1(_11056_),
    .X(_02820_));
 sky130_fd_sc_hd__buf_2 _25588_ (.A(_10055_),
    .X(_11057_));
 sky130_fd_sc_hd__and2_1 _25589_ (.A(_10408_),
    .B(_11055_),
    .X(_11058_));
 sky130_fd_sc_hd__a31o_1 _25590_ (.A1(_11057_),
    .A2(\datamem.data_ram[21][1] ),
    .A3(_11053_),
    .B1(_11058_),
    .X(_02821_));
 sky130_fd_sc_hd__and2_1 _25591_ (.A(_10410_),
    .B(_11055_),
    .X(_11059_));
 sky130_fd_sc_hd__a31o_1 _25592_ (.A1(_11057_),
    .A2(\datamem.data_ram[21][2] ),
    .A3(_11053_),
    .B1(_11059_),
    .X(_02822_));
 sky130_fd_sc_hd__and2_1 _25593_ (.A(_10413_),
    .B(_11055_),
    .X(_11060_));
 sky130_fd_sc_hd__a31o_1 _25594_ (.A1(_11057_),
    .A2(\datamem.data_ram[21][3] ),
    .A3(_11053_),
    .B1(_11060_),
    .X(_02823_));
 sky130_fd_sc_hd__and2_1 _25595_ (.A(_11047_),
    .B(_11055_),
    .X(_11061_));
 sky130_fd_sc_hd__a31o_1 _25596_ (.A1(_11057_),
    .A2(\datamem.data_ram[21][4] ),
    .A3(_11053_),
    .B1(_11061_),
    .X(_02824_));
 sky130_fd_sc_hd__and2_1 _25597_ (.A(_10416_),
    .B(_11055_),
    .X(_11062_));
 sky130_fd_sc_hd__a31o_1 _25598_ (.A1(_11057_),
    .A2(\datamem.data_ram[21][5] ),
    .A3(_11053_),
    .B1(_11062_),
    .X(_02825_));
 sky130_fd_sc_hd__and2_1 _25599_ (.A(_10418_),
    .B(_11055_),
    .X(_11063_));
 sky130_fd_sc_hd__a31o_1 _25600_ (.A1(_11057_),
    .A2(\datamem.data_ram[21][6] ),
    .A3(_11053_),
    .B1(_11063_),
    .X(_02826_));
 sky130_fd_sc_hd__clkbuf_4 _25601_ (.A(_10075_),
    .X(_11064_));
 sky130_fd_sc_hd__and2_1 _25602_ (.A(_11064_),
    .B(_11055_),
    .X(_11065_));
 sky130_fd_sc_hd__a31o_1 _25603_ (.A1(_11057_),
    .A2(\datamem.data_ram[21][7] ),
    .A3(_11053_),
    .B1(_11065_),
    .X(_02827_));
 sky130_fd_sc_hd__a21oi_1 _25604_ (.A1(_10570_),
    .A2(_11020_),
    .B1(_10998_),
    .Y(_11066_));
 sky130_fd_sc_hd__mux2_1 _25605_ (.A0(_10724_),
    .A1(\datamem.data_ram[9][8] ),
    .S(net53),
    .X(_11067_));
 sky130_fd_sc_hd__clkbuf_1 _25606_ (.A(_11067_),
    .X(_02828_));
 sky130_fd_sc_hd__mux2_1 _25607_ (.A0(_10727_),
    .A1(\datamem.data_ram[9][9] ),
    .S(net53),
    .X(_11068_));
 sky130_fd_sc_hd__clkbuf_1 _25608_ (.A(_11068_),
    .X(_02829_));
 sky130_fd_sc_hd__mux2_1 _25609_ (.A0(_10729_),
    .A1(\datamem.data_ram[9][10] ),
    .S(net53),
    .X(_11069_));
 sky130_fd_sc_hd__clkbuf_1 _25610_ (.A(_11069_),
    .X(_02830_));
 sky130_fd_sc_hd__mux2_1 _25611_ (.A0(_10731_),
    .A1(\datamem.data_ram[9][11] ),
    .S(net53),
    .X(_11070_));
 sky130_fd_sc_hd__clkbuf_1 _25612_ (.A(_11070_),
    .X(_02831_));
 sky130_fd_sc_hd__mux2_1 _25613_ (.A0(_10733_),
    .A1(\datamem.data_ram[9][12] ),
    .S(net53),
    .X(_11071_));
 sky130_fd_sc_hd__clkbuf_1 _25614_ (.A(_11071_),
    .X(_02832_));
 sky130_fd_sc_hd__mux2_1 _25615_ (.A0(_10735_),
    .A1(\datamem.data_ram[9][13] ),
    .S(net53),
    .X(_11072_));
 sky130_fd_sc_hd__clkbuf_1 _25616_ (.A(_11072_),
    .X(_02833_));
 sky130_fd_sc_hd__mux2_1 _25617_ (.A0(_10737_),
    .A1(\datamem.data_ram[9][14] ),
    .S(net53),
    .X(_11073_));
 sky130_fd_sc_hd__clkbuf_1 _25618_ (.A(_11073_),
    .X(_02834_));
 sky130_fd_sc_hd__mux2_1 _25619_ (.A0(_10739_),
    .A1(\datamem.data_ram[9][15] ),
    .S(net53),
    .X(_11074_));
 sky130_fd_sc_hd__clkbuf_1 _25620_ (.A(_11074_),
    .X(_02835_));
 sky130_fd_sc_hd__nand2_8 _25621_ (.A(_10141_),
    .B(_10051_),
    .Y(_11075_));
 sky130_fd_sc_hd__or2_1 _25622_ (.A(_10946_),
    .B(_11075_),
    .X(_11076_));
 sky130_fd_sc_hd__buf_2 _25623_ (.A(_11076_),
    .X(_11077_));
 sky130_fd_sc_hd__clkbuf_4 _25624_ (.A(_10047_),
    .X(_11078_));
 sky130_fd_sc_hd__nor2_2 _25625_ (.A(_10946_),
    .B(_11075_),
    .Y(_11079_));
 sky130_fd_sc_hd__and2_1 _25626_ (.A(_11078_),
    .B(_11079_),
    .X(_11080_));
 sky130_fd_sc_hd__a31o_1 _25627_ (.A1(_11057_),
    .A2(\datamem.data_ram[19][0] ),
    .A3(_11077_),
    .B1(_11080_),
    .X(_02836_));
 sky130_fd_sc_hd__clkbuf_4 _25628_ (.A(_10057_),
    .X(_11081_));
 sky130_fd_sc_hd__and2_1 _25629_ (.A(_11081_),
    .B(_11079_),
    .X(_11082_));
 sky130_fd_sc_hd__a31o_1 _25630_ (.A1(_11057_),
    .A2(\datamem.data_ram[19][1] ),
    .A3(_11077_),
    .B1(_11082_),
    .X(_02837_));
 sky130_fd_sc_hd__clkbuf_4 _25631_ (.A(_10060_),
    .X(_11083_));
 sky130_fd_sc_hd__and2_1 _25632_ (.A(_11083_),
    .B(_11079_),
    .X(_11084_));
 sky130_fd_sc_hd__a31o_1 _25633_ (.A1(_11057_),
    .A2(\datamem.data_ram[19][2] ),
    .A3(_11077_),
    .B1(_11084_),
    .X(_02838_));
 sky130_fd_sc_hd__buf_2 _25634_ (.A(_10055_),
    .X(_11085_));
 sky130_fd_sc_hd__clkbuf_4 _25635_ (.A(_10063_),
    .X(_11086_));
 sky130_fd_sc_hd__and2_1 _25636_ (.A(_11086_),
    .B(_11079_),
    .X(_11087_));
 sky130_fd_sc_hd__a31o_1 _25637_ (.A1(_11085_),
    .A2(\datamem.data_ram[19][3] ),
    .A3(_11077_),
    .B1(_11087_),
    .X(_02839_));
 sky130_fd_sc_hd__and2_1 _25638_ (.A(_11047_),
    .B(_11079_),
    .X(_11088_));
 sky130_fd_sc_hd__a31o_1 _25639_ (.A1(_11085_),
    .A2(\datamem.data_ram[19][4] ),
    .A3(_11077_),
    .B1(_11088_),
    .X(_02840_));
 sky130_fd_sc_hd__clkbuf_4 _25640_ (.A(_10069_),
    .X(_11089_));
 sky130_fd_sc_hd__and2_1 _25641_ (.A(_11089_),
    .B(_11079_),
    .X(_11090_));
 sky130_fd_sc_hd__a31o_1 _25642_ (.A1(_11085_),
    .A2(\datamem.data_ram[19][5] ),
    .A3(_11077_),
    .B1(_11090_),
    .X(_02841_));
 sky130_fd_sc_hd__clkbuf_4 _25643_ (.A(_10072_),
    .X(_11091_));
 sky130_fd_sc_hd__and2_1 _25644_ (.A(_11091_),
    .B(_11079_),
    .X(_11092_));
 sky130_fd_sc_hd__a31o_1 _25645_ (.A1(_11085_),
    .A2(\datamem.data_ram[19][6] ),
    .A3(_11077_),
    .B1(_11092_),
    .X(_02842_));
 sky130_fd_sc_hd__and2_1 _25646_ (.A(_11064_),
    .B(_11079_),
    .X(_11093_));
 sky130_fd_sc_hd__a31o_1 _25647_ (.A1(_11085_),
    .A2(\datamem.data_ram[19][7] ),
    .A3(_11077_),
    .B1(_11093_),
    .X(_02843_));
 sky130_fd_sc_hd__nor2_2 _25648_ (.A(_10600_),
    .B(_11075_),
    .Y(_11094_));
 sky130_fd_sc_hd__nor2_2 _25649_ (.A(_10780_),
    .B(_11094_),
    .Y(_11095_));
 sky130_fd_sc_hd__a22o_1 _25650_ (.A1(_10048_),
    .A2(_11094_),
    .B1(_11095_),
    .B2(\datamem.data_ram[43][0] ),
    .X(_02844_));
 sky130_fd_sc_hd__a22o_1 _25651_ (.A1(_10058_),
    .A2(_11094_),
    .B1(_11095_),
    .B2(\datamem.data_ram[43][1] ),
    .X(_02845_));
 sky130_fd_sc_hd__a22o_1 _25652_ (.A1(_10061_),
    .A2(_11094_),
    .B1(_11095_),
    .B2(\datamem.data_ram[43][2] ),
    .X(_02846_));
 sky130_fd_sc_hd__a22o_1 _25653_ (.A1(_10064_),
    .A2(_11094_),
    .B1(_11095_),
    .B2(\datamem.data_ram[43][3] ),
    .X(_02847_));
 sky130_fd_sc_hd__a22o_1 _25654_ (.A1(_10782_),
    .A2(_11094_),
    .B1(_11095_),
    .B2(\datamem.data_ram[43][4] ),
    .X(_02848_));
 sky130_fd_sc_hd__a22o_1 _25655_ (.A1(_10070_),
    .A2(_11094_),
    .B1(_11095_),
    .B2(\datamem.data_ram[43][5] ),
    .X(_02849_));
 sky130_fd_sc_hd__a22o_1 _25656_ (.A1(_10073_),
    .A2(_11094_),
    .B1(_11095_),
    .B2(\datamem.data_ram[43][6] ),
    .X(_02850_));
 sky130_fd_sc_hd__a22o_1 _25657_ (.A1(_10783_),
    .A2(_11094_),
    .B1(_11095_),
    .B2(\datamem.data_ram[43][7] ),
    .X(_02851_));
 sky130_fd_sc_hd__or3_1 _25658_ (.A(_07077_),
    .B(_10918_),
    .C(_10897_),
    .X(_11096_));
 sky130_fd_sc_hd__clkbuf_2 _25659_ (.A(_11096_),
    .X(_11097_));
 sky130_fd_sc_hd__and3_2 _25660_ (.A(_10142_),
    .B(_10921_),
    .C(_10922_),
    .X(_11098_));
 sky130_fd_sc_hd__and2_1 _25661_ (.A(_11078_),
    .B(_11098_),
    .X(_11099_));
 sky130_fd_sc_hd__a31o_1 _25662_ (.A1(_11085_),
    .A2(\datamem.data_ram[35][0] ),
    .A3(_11097_),
    .B1(_11099_),
    .X(_02852_));
 sky130_fd_sc_hd__and2_1 _25663_ (.A(_11081_),
    .B(_11098_),
    .X(_11100_));
 sky130_fd_sc_hd__a31o_1 _25664_ (.A1(_11085_),
    .A2(\datamem.data_ram[35][1] ),
    .A3(_11097_),
    .B1(_11100_),
    .X(_02853_));
 sky130_fd_sc_hd__and2_1 _25665_ (.A(_11083_),
    .B(_11098_),
    .X(_11101_));
 sky130_fd_sc_hd__a31o_1 _25666_ (.A1(_11085_),
    .A2(\datamem.data_ram[35][2] ),
    .A3(_11097_),
    .B1(_11101_),
    .X(_02854_));
 sky130_fd_sc_hd__and2_1 _25667_ (.A(_11086_),
    .B(_11098_),
    .X(_11102_));
 sky130_fd_sc_hd__a31o_1 _25668_ (.A1(_11085_),
    .A2(\datamem.data_ram[35][3] ),
    .A3(_11097_),
    .B1(_11102_),
    .X(_02855_));
 sky130_fd_sc_hd__and2_1 _25669_ (.A(_11047_),
    .B(_11098_),
    .X(_11103_));
 sky130_fd_sc_hd__a31o_1 _25670_ (.A1(_11085_),
    .A2(\datamem.data_ram[35][4] ),
    .A3(_11097_),
    .B1(_11103_),
    .X(_02856_));
 sky130_fd_sc_hd__buf_2 _25671_ (.A(_06587_),
    .X(_11104_));
 sky130_fd_sc_hd__clkbuf_4 _25672_ (.A(_11104_),
    .X(_11105_));
 sky130_fd_sc_hd__and2_1 _25673_ (.A(_11089_),
    .B(_11098_),
    .X(_11106_));
 sky130_fd_sc_hd__a31o_1 _25674_ (.A1(_11105_),
    .A2(\datamem.data_ram[35][5] ),
    .A3(_11097_),
    .B1(_11106_),
    .X(_02857_));
 sky130_fd_sc_hd__and2_1 _25675_ (.A(_11091_),
    .B(_11098_),
    .X(_11107_));
 sky130_fd_sc_hd__a31o_1 _25676_ (.A1(_11105_),
    .A2(\datamem.data_ram[35][6] ),
    .A3(_11097_),
    .B1(_11107_),
    .X(_02858_));
 sky130_fd_sc_hd__and2_1 _25677_ (.A(_11064_),
    .B(_11098_),
    .X(_11108_));
 sky130_fd_sc_hd__a31o_1 _25678_ (.A1(_11105_),
    .A2(\datamem.data_ram[35][7] ),
    .A3(_11097_),
    .B1(_11108_),
    .X(_02859_));
 sky130_fd_sc_hd__buf_2 _25679_ (.A(_08125_),
    .X(_11109_));
 sky130_fd_sc_hd__or3_1 _25680_ (.A(_07808_),
    .B(_11109_),
    .C(_10044_),
    .X(_11110_));
 sky130_fd_sc_hd__clkbuf_2 _25681_ (.A(_11110_),
    .X(_11111_));
 sky130_fd_sc_hd__nor2_1 _25682_ (.A(_07131_),
    .B(_07177_),
    .Y(_11112_));
 sky130_fd_sc_hd__and3_2 _25683_ (.A(_10268_),
    .B(_11112_),
    .C(_10052_),
    .X(_11113_));
 sky130_fd_sc_hd__and2_1 _25684_ (.A(_11078_),
    .B(_11113_),
    .X(_11114_));
 sky130_fd_sc_hd__a31o_1 _25685_ (.A1(_11105_),
    .A2(\datamem.data_ram[25][0] ),
    .A3(_11111_),
    .B1(_11114_),
    .X(_02860_));
 sky130_fd_sc_hd__and2_1 _25686_ (.A(_11081_),
    .B(_11113_),
    .X(_11115_));
 sky130_fd_sc_hd__a31o_1 _25687_ (.A1(_11105_),
    .A2(\datamem.data_ram[25][1] ),
    .A3(_11111_),
    .B1(_11115_),
    .X(_02861_));
 sky130_fd_sc_hd__and2_1 _25688_ (.A(_11083_),
    .B(_11113_),
    .X(_11116_));
 sky130_fd_sc_hd__a31o_1 _25689_ (.A1(_11105_),
    .A2(\datamem.data_ram[25][2] ),
    .A3(_11111_),
    .B1(_11116_),
    .X(_02862_));
 sky130_fd_sc_hd__and2_1 _25690_ (.A(_11086_),
    .B(_11113_),
    .X(_11117_));
 sky130_fd_sc_hd__a31o_1 _25691_ (.A1(_11105_),
    .A2(\datamem.data_ram[25][3] ),
    .A3(_11111_),
    .B1(_11117_),
    .X(_02863_));
 sky130_fd_sc_hd__and2_1 _25692_ (.A(_11047_),
    .B(_11113_),
    .X(_11118_));
 sky130_fd_sc_hd__a31o_1 _25693_ (.A1(_11105_),
    .A2(\datamem.data_ram[25][4] ),
    .A3(_11111_),
    .B1(_11118_),
    .X(_02864_));
 sky130_fd_sc_hd__and2_1 _25694_ (.A(_11089_),
    .B(_11113_),
    .X(_11119_));
 sky130_fd_sc_hd__a31o_1 _25695_ (.A1(_11105_),
    .A2(\datamem.data_ram[25][5] ),
    .A3(_11111_),
    .B1(_11119_),
    .X(_02865_));
 sky130_fd_sc_hd__and2_1 _25696_ (.A(_11091_),
    .B(_11113_),
    .X(_11120_));
 sky130_fd_sc_hd__a31o_1 _25697_ (.A1(_11105_),
    .A2(\datamem.data_ram[25][6] ),
    .A3(_11111_),
    .B1(_11120_),
    .X(_02866_));
 sky130_fd_sc_hd__clkbuf_4 _25698_ (.A(_11104_),
    .X(_11121_));
 sky130_fd_sc_hd__and2_1 _25699_ (.A(_11064_),
    .B(_11113_),
    .X(_11122_));
 sky130_fd_sc_hd__a31o_1 _25700_ (.A1(_11121_),
    .A2(\datamem.data_ram[25][7] ),
    .A3(_11111_),
    .B1(_11122_),
    .X(_02867_));
 sky130_fd_sc_hd__nor2_8 _25701_ (.A(_08144_),
    .B(net109),
    .Y(_11123_));
 sky130_fd_sc_hd__a21oi_4 _25702_ (.A1(_10542_),
    .A2(_11123_),
    .B1(_10998_),
    .Y(_11124_));
 sky130_fd_sc_hd__mux2_1 _25703_ (.A0(_10811_),
    .A1(\datamem.data_ram[4][24] ),
    .S(_11124_),
    .X(_11125_));
 sky130_fd_sc_hd__clkbuf_1 _25704_ (.A(_11125_),
    .X(_02868_));
 sky130_fd_sc_hd__mux2_1 _25705_ (.A0(_10814_),
    .A1(\datamem.data_ram[4][25] ),
    .S(_11124_),
    .X(_11126_));
 sky130_fd_sc_hd__clkbuf_1 _25706_ (.A(_11126_),
    .X(_02869_));
 sky130_fd_sc_hd__mux2_1 _25707_ (.A0(_10816_),
    .A1(\datamem.data_ram[4][26] ),
    .S(_11124_),
    .X(_11127_));
 sky130_fd_sc_hd__clkbuf_1 _25708_ (.A(_11127_),
    .X(_02870_));
 sky130_fd_sc_hd__mux2_1 _25709_ (.A0(_10818_),
    .A1(\datamem.data_ram[4][27] ),
    .S(_11124_),
    .X(_11128_));
 sky130_fd_sc_hd__clkbuf_1 _25710_ (.A(_11128_),
    .X(_02871_));
 sky130_fd_sc_hd__mux2_1 _25711_ (.A0(_10820_),
    .A1(\datamem.data_ram[4][28] ),
    .S(_11124_),
    .X(_11129_));
 sky130_fd_sc_hd__clkbuf_1 _25712_ (.A(_11129_),
    .X(_02872_));
 sky130_fd_sc_hd__mux2_1 _25713_ (.A0(_10822_),
    .A1(\datamem.data_ram[4][29] ),
    .S(_11124_),
    .X(_11130_));
 sky130_fd_sc_hd__clkbuf_1 _25714_ (.A(_11130_),
    .X(_02873_));
 sky130_fd_sc_hd__mux2_1 _25715_ (.A0(_10824_),
    .A1(\datamem.data_ram[4][30] ),
    .S(_11124_),
    .X(_11131_));
 sky130_fd_sc_hd__clkbuf_1 _25716_ (.A(_11131_),
    .X(_02874_));
 sky130_fd_sc_hd__mux2_1 _25717_ (.A0(_10826_),
    .A1(\datamem.data_ram[4][31] ),
    .S(_11124_),
    .X(_11132_));
 sky130_fd_sc_hd__clkbuf_1 _25718_ (.A(_11132_),
    .X(_02875_));
 sky130_fd_sc_hd__a21oi_4 _25719_ (.A1(_10113_),
    .A2(_11123_),
    .B1(_10998_),
    .Y(_11133_));
 sky130_fd_sc_hd__mux2_1 _25720_ (.A0(_10811_),
    .A1(\datamem.data_ram[5][24] ),
    .S(_11133_),
    .X(_11134_));
 sky130_fd_sc_hd__clkbuf_1 _25721_ (.A(_11134_),
    .X(_02876_));
 sky130_fd_sc_hd__mux2_1 _25722_ (.A0(_10814_),
    .A1(\datamem.data_ram[5][25] ),
    .S(_11133_),
    .X(_11135_));
 sky130_fd_sc_hd__clkbuf_1 _25723_ (.A(_11135_),
    .X(_02877_));
 sky130_fd_sc_hd__mux2_1 _25724_ (.A0(_10816_),
    .A1(\datamem.data_ram[5][26] ),
    .S(_11133_),
    .X(_11136_));
 sky130_fd_sc_hd__clkbuf_1 _25725_ (.A(_11136_),
    .X(_02878_));
 sky130_fd_sc_hd__mux2_1 _25726_ (.A0(_10818_),
    .A1(\datamem.data_ram[5][27] ),
    .S(_11133_),
    .X(_11137_));
 sky130_fd_sc_hd__clkbuf_1 _25727_ (.A(_11137_),
    .X(_02879_));
 sky130_fd_sc_hd__mux2_1 _25728_ (.A0(_10820_),
    .A1(\datamem.data_ram[5][28] ),
    .S(_11133_),
    .X(_11138_));
 sky130_fd_sc_hd__clkbuf_1 _25729_ (.A(_11138_),
    .X(_02880_));
 sky130_fd_sc_hd__mux2_1 _25730_ (.A0(_10822_),
    .A1(\datamem.data_ram[5][29] ),
    .S(_11133_),
    .X(_11139_));
 sky130_fd_sc_hd__clkbuf_1 _25731_ (.A(_11139_),
    .X(_02881_));
 sky130_fd_sc_hd__mux2_1 _25732_ (.A0(_10824_),
    .A1(\datamem.data_ram[5][30] ),
    .S(_11133_),
    .X(_11140_));
 sky130_fd_sc_hd__clkbuf_1 _25733_ (.A(_11140_),
    .X(_02882_));
 sky130_fd_sc_hd__mux2_1 _25734_ (.A0(_10826_),
    .A1(\datamem.data_ram[5][31] ),
    .S(_11133_),
    .X(_11141_));
 sky130_fd_sc_hd__clkbuf_1 _25735_ (.A(_11141_),
    .X(_02883_));
 sky130_fd_sc_hd__clkbuf_4 _25736_ (.A(_08598_),
    .X(_11142_));
 sky130_fd_sc_hd__clkbuf_4 _25737_ (.A(_11142_),
    .X(_11143_));
 sky130_fd_sc_hd__clkbuf_4 _25738_ (.A(_11143_),
    .X(_11144_));
 sky130_fd_sc_hd__and2_1 _25739_ (.A(_08620_),
    .B(_08621_),
    .X(_11145_));
 sky130_fd_sc_hd__clkbuf_4 _25740_ (.A(_11145_),
    .X(_11146_));
 sky130_fd_sc_hd__clkbuf_4 _25741_ (.A(_11146_),
    .X(_11147_));
 sky130_fd_sc_hd__nand2_1 _25742_ (.A(_13328_),
    .B(_11142_),
    .Y(_11148_));
 sky130_fd_sc_hd__o211a_1 _25743_ (.A1(\rvcpu.dp.plfd.PCPlus4D[2] ),
    .A2(_11144_),
    .B1(_11147_),
    .C1(_11148_),
    .X(_02884_));
 sky130_fd_sc_hd__buf_2 _25744_ (.A(_08598_),
    .X(_11149_));
 sky130_fd_sc_hd__nand2_1 _25745_ (.A(_13391_),
    .B(_11149_),
    .Y(_11150_));
 sky130_fd_sc_hd__o211a_1 _25746_ (.A1(\rvcpu.dp.plfd.PCPlus4D[3] ),
    .A2(_11144_),
    .B1(_11147_),
    .C1(_11150_),
    .X(_02885_));
 sky130_fd_sc_hd__o21a_1 _25747_ (.A1(_08588_),
    .A2(_08597_),
    .B1(\rvcpu.dp.hu.ResultSrcE0 ),
    .X(_11151_));
 sky130_fd_sc_hd__buf_2 _25748_ (.A(_11151_),
    .X(_11152_));
 sky130_fd_sc_hd__clkbuf_4 _25749_ (.A(_11152_),
    .X(_11153_));
 sky130_fd_sc_hd__nand2_1 _25750_ (.A(_13335_),
    .B(_13717_),
    .Y(_11154_));
 sky130_fd_sc_hd__clkbuf_2 _25751_ (.A(_08598_),
    .X(_11155_));
 sky130_fd_sc_hd__or2_1 _25752_ (.A(\rvcpu.dp.plfd.PCPlus4D[4] ),
    .B(_11155_),
    .X(_11156_));
 sky130_fd_sc_hd__o211a_1 _25753_ (.A1(_11153_),
    .A2(_11154_),
    .B1(_11156_),
    .C1(_11147_),
    .X(_02886_));
 sky130_fd_sc_hd__buf_4 _25754_ (.A(_11151_),
    .X(_11157_));
 sky130_fd_sc_hd__or3b_1 _25755_ (.A(_13865_),
    .B(_11157_),
    .C_N(_13758_),
    .X(_11158_));
 sky130_fd_sc_hd__o211a_1 _25756_ (.A1(\rvcpu.dp.plfd.PCPlus4D[5] ),
    .A2(_11144_),
    .B1(_11147_),
    .C1(_11158_),
    .X(_02887_));
 sky130_fd_sc_hd__nand2_1 _25757_ (.A(_13823_),
    .B(_13876_),
    .Y(_11159_));
 sky130_fd_sc_hd__or2_1 _25758_ (.A(_13823_),
    .B(_13876_),
    .X(_11160_));
 sky130_fd_sc_hd__a21o_1 _25759_ (.A1(_11159_),
    .A2(_11160_),
    .B1(_11152_),
    .X(_11161_));
 sky130_fd_sc_hd__o211a_1 _25760_ (.A1(\rvcpu.dp.plfd.PCPlus4D[6] ),
    .A2(_11144_),
    .B1(_11147_),
    .C1(_11161_),
    .X(_02888_));
 sky130_fd_sc_hd__a21oi_1 _25761_ (.A1(_13823_),
    .A2(_13876_),
    .B1(_13706_),
    .Y(_11162_));
 sky130_fd_sc_hd__a21o_1 _25762_ (.A1(_13463_),
    .A2(_13876_),
    .B1(_11162_),
    .X(_11163_));
 sky130_fd_sc_hd__nand2_1 _25763_ (.A(_11149_),
    .B(_11163_),
    .Y(_11164_));
 sky130_fd_sc_hd__o211a_1 _25764_ (.A1(\rvcpu.dp.plfd.PCPlus4D[7] ),
    .A2(_11144_),
    .B1(_11147_),
    .C1(_11164_),
    .X(_02889_));
 sky130_fd_sc_hd__nand2_1 _25765_ (.A(_13514_),
    .B(_13876_),
    .Y(_11165_));
 sky130_fd_sc_hd__a31o_1 _25766_ (.A1(_13463_),
    .A2(_13301_),
    .A3(_13294_),
    .B1(_13439_),
    .X(_11166_));
 sky130_fd_sc_hd__a21o_1 _25767_ (.A1(_11165_),
    .A2(_11166_),
    .B1(_11157_),
    .X(_11167_));
 sky130_fd_sc_hd__o211a_1 _25768_ (.A1(\rvcpu.dp.plfd.PCPlus4D[8] ),
    .A2(_11144_),
    .B1(_11147_),
    .C1(_11167_),
    .X(_02890_));
 sky130_fd_sc_hd__nor2_1 _25769_ (.A(_13538_),
    .B(_11165_),
    .Y(_11168_));
 sky130_fd_sc_hd__and3_1 _25770_ (.A(_13539_),
    .B(_08598_),
    .C(_11165_),
    .X(_11169_));
 sky130_fd_sc_hd__a21oi_1 _25771_ (.A1(_11149_),
    .A2(_11168_),
    .B1(_11169_),
    .Y(_11170_));
 sky130_fd_sc_hd__o211a_1 _25772_ (.A1(\rvcpu.dp.plfd.PCPlus4D[9] ),
    .A2(_11144_),
    .B1(_11147_),
    .C1(_11170_),
    .X(_02891_));
 sky130_fd_sc_hd__and2_1 _25773_ (.A(\rvcpu.dp.pcreg.q[10] ),
    .B(_11168_),
    .X(_11171_));
 sky130_fd_sc_hd__nor2_1 _25774_ (.A(\rvcpu.dp.pcreg.q[10] ),
    .B(_11168_),
    .Y(_11172_));
 sky130_fd_sc_hd__o21ai_1 _25775_ (.A1(_11171_),
    .A2(_11172_),
    .B1(_11149_),
    .Y(_11173_));
 sky130_fd_sc_hd__o211a_1 _25776_ (.A1(\rvcpu.dp.plfd.PCPlus4D[10] ),
    .A2(_11144_),
    .B1(_11147_),
    .C1(_11173_),
    .X(_02892_));
 sky130_fd_sc_hd__nand2_1 _25777_ (.A(\rvcpu.dp.pcreg.q[11] ),
    .B(_11171_),
    .Y(_11174_));
 sky130_fd_sc_hd__or2_1 _25778_ (.A(\rvcpu.dp.pcreg.q[11] ),
    .B(_11171_),
    .X(_11175_));
 sky130_fd_sc_hd__a21o_1 _25779_ (.A1(_11174_),
    .A2(_11175_),
    .B1(_11157_),
    .X(_11176_));
 sky130_fd_sc_hd__o211a_1 _25780_ (.A1(\rvcpu.dp.plfd.PCPlus4D[11] ),
    .A2(_11144_),
    .B1(_11147_),
    .C1(_11176_),
    .X(_02893_));
 sky130_fd_sc_hd__clkbuf_4 _25781_ (.A(_11146_),
    .X(_11177_));
 sky130_fd_sc_hd__and3_1 _25782_ (.A(\rvcpu.dp.pcreg.q[12] ),
    .B(\rvcpu.dp.pcreg.q[11] ),
    .C(_11171_),
    .X(_11178_));
 sky130_fd_sc_hd__a21oi_1 _25783_ (.A1(\rvcpu.dp.pcreg.q[11] ),
    .A2(_11171_),
    .B1(\rvcpu.dp.pcreg.q[12] ),
    .Y(_11179_));
 sky130_fd_sc_hd__o21ai_1 _25784_ (.A1(_11178_),
    .A2(_11179_),
    .B1(_11149_),
    .Y(_11180_));
 sky130_fd_sc_hd__o211a_1 _25785_ (.A1(\rvcpu.dp.plfd.PCPlus4D[12] ),
    .A2(_11144_),
    .B1(_11177_),
    .C1(_11180_),
    .X(_02894_));
 sky130_fd_sc_hd__clkbuf_4 _25786_ (.A(_11143_),
    .X(_11181_));
 sky130_fd_sc_hd__and2_1 _25787_ (.A(\rvcpu.dp.pcreg.q[13] ),
    .B(_11178_),
    .X(_11182_));
 sky130_fd_sc_hd__nor2_1 _25788_ (.A(\rvcpu.dp.pcreg.q[13] ),
    .B(_11178_),
    .Y(_11183_));
 sky130_fd_sc_hd__o21ai_1 _25789_ (.A1(_11182_),
    .A2(_11183_),
    .B1(_11149_),
    .Y(_11184_));
 sky130_fd_sc_hd__o211a_1 _25790_ (.A1(\rvcpu.dp.plfd.PCPlus4D[13] ),
    .A2(_11181_),
    .B1(_11177_),
    .C1(_11184_),
    .X(_02895_));
 sky130_fd_sc_hd__nand2_1 _25791_ (.A(\rvcpu.dp.pcreg.q[14] ),
    .B(_11182_),
    .Y(_11185_));
 sky130_fd_sc_hd__or2_1 _25792_ (.A(\rvcpu.dp.pcreg.q[14] ),
    .B(_11182_),
    .X(_11186_));
 sky130_fd_sc_hd__a21o_1 _25793_ (.A1(_11185_),
    .A2(_11186_),
    .B1(_11157_),
    .X(_11187_));
 sky130_fd_sc_hd__o211a_1 _25794_ (.A1(\rvcpu.dp.plfd.PCPlus4D[14] ),
    .A2(_11181_),
    .B1(_11177_),
    .C1(_11187_),
    .X(_02896_));
 sky130_fd_sc_hd__and3_1 _25795_ (.A(\rvcpu.dp.pcreg.q[15] ),
    .B(\rvcpu.dp.pcreg.q[14] ),
    .C(_11182_),
    .X(_11188_));
 sky130_fd_sc_hd__a21oi_1 _25796_ (.A1(\rvcpu.dp.pcreg.q[14] ),
    .A2(_11182_),
    .B1(\rvcpu.dp.pcreg.q[15] ),
    .Y(_11189_));
 sky130_fd_sc_hd__o21ai_1 _25797_ (.A1(_11188_),
    .A2(_11189_),
    .B1(_11149_),
    .Y(_11190_));
 sky130_fd_sc_hd__o211a_1 _25798_ (.A1(\rvcpu.dp.plfd.PCPlus4D[15] ),
    .A2(_11181_),
    .B1(_11177_),
    .C1(_11190_),
    .X(_02897_));
 sky130_fd_sc_hd__and2_1 _25799_ (.A(\rvcpu.dp.pcreg.q[16] ),
    .B(_11188_),
    .X(_11191_));
 sky130_fd_sc_hd__nor2_1 _25800_ (.A(\rvcpu.dp.pcreg.q[16] ),
    .B(_11188_),
    .Y(_11192_));
 sky130_fd_sc_hd__o21ai_1 _25801_ (.A1(_11191_),
    .A2(_11192_),
    .B1(_11149_),
    .Y(_11193_));
 sky130_fd_sc_hd__o211a_1 _25802_ (.A1(\rvcpu.dp.plfd.PCPlus4D[16] ),
    .A2(_11181_),
    .B1(_11177_),
    .C1(_11193_),
    .X(_02898_));
 sky130_fd_sc_hd__nand2_1 _25803_ (.A(\rvcpu.dp.pcreg.q[17] ),
    .B(_11191_),
    .Y(_11194_));
 sky130_fd_sc_hd__or2_1 _25804_ (.A(\rvcpu.dp.pcreg.q[17] ),
    .B(_11191_),
    .X(_11195_));
 sky130_fd_sc_hd__a21o_1 _25805_ (.A1(_11194_),
    .A2(_11195_),
    .B1(_11157_),
    .X(_11196_));
 sky130_fd_sc_hd__o211a_1 _25806_ (.A1(\rvcpu.dp.plfd.PCPlus4D[17] ),
    .A2(_11181_),
    .B1(_11177_),
    .C1(_11196_),
    .X(_02899_));
 sky130_fd_sc_hd__and3_1 _25807_ (.A(\rvcpu.dp.pcreg.q[18] ),
    .B(\rvcpu.dp.pcreg.q[17] ),
    .C(_11191_),
    .X(_11197_));
 sky130_fd_sc_hd__a21oi_1 _25808_ (.A1(\rvcpu.dp.pcreg.q[17] ),
    .A2(_11191_),
    .B1(\rvcpu.dp.pcreg.q[18] ),
    .Y(_11198_));
 sky130_fd_sc_hd__o21ai_1 _25809_ (.A1(_11197_),
    .A2(_11198_),
    .B1(_11149_),
    .Y(_11199_));
 sky130_fd_sc_hd__o211a_1 _25810_ (.A1(\rvcpu.dp.plfd.PCPlus4D[18] ),
    .A2(_11181_),
    .B1(_11177_),
    .C1(_11199_),
    .X(_02900_));
 sky130_fd_sc_hd__and2_1 _25811_ (.A(\rvcpu.dp.pcreg.q[19] ),
    .B(_11197_),
    .X(_11200_));
 sky130_fd_sc_hd__nor2_1 _25812_ (.A(\rvcpu.dp.pcreg.q[19] ),
    .B(_11197_),
    .Y(_11201_));
 sky130_fd_sc_hd__o21ai_1 _25813_ (.A1(_11200_),
    .A2(_11201_),
    .B1(_11149_),
    .Y(_11202_));
 sky130_fd_sc_hd__o211a_1 _25814_ (.A1(\rvcpu.dp.plfd.PCPlus4D[19] ),
    .A2(_11181_),
    .B1(_11177_),
    .C1(_11202_),
    .X(_02901_));
 sky130_fd_sc_hd__nand2_1 _25815_ (.A(\rvcpu.dp.pcreg.q[20] ),
    .B(_11200_),
    .Y(_11203_));
 sky130_fd_sc_hd__or2_1 _25816_ (.A(\rvcpu.dp.pcreg.q[20] ),
    .B(_11200_),
    .X(_11204_));
 sky130_fd_sc_hd__a21o_1 _25817_ (.A1(_11203_),
    .A2(_11204_),
    .B1(_11157_),
    .X(_11205_));
 sky130_fd_sc_hd__o211a_1 _25818_ (.A1(\rvcpu.dp.plfd.PCPlus4D[20] ),
    .A2(_11181_),
    .B1(_11177_),
    .C1(_11205_),
    .X(_02902_));
 sky130_fd_sc_hd__clkbuf_2 _25819_ (.A(_08620_),
    .X(_11206_));
 sky130_fd_sc_hd__clkbuf_2 _25820_ (.A(_08621_),
    .X(_11207_));
 sky130_fd_sc_hd__and3_1 _25821_ (.A(\rvcpu.dp.pcreg.q[21] ),
    .B(\rvcpu.dp.pcreg.q[20] ),
    .C(_11200_),
    .X(_11208_));
 sky130_fd_sc_hd__a21oi_1 _25822_ (.A1(\rvcpu.dp.pcreg.q[20] ),
    .A2(_11200_),
    .B1(\rvcpu.dp.pcreg.q[21] ),
    .Y(_11209_));
 sky130_fd_sc_hd__nor2_1 _25823_ (.A(_11208_),
    .B(_11209_),
    .Y(_11210_));
 sky130_fd_sc_hd__mux2_1 _25824_ (.A0(\rvcpu.dp.plfd.PCPlus4D[21] ),
    .A1(_11210_),
    .S(_11142_),
    .X(_11211_));
 sky130_fd_sc_hd__and3_1 _25825_ (.A(_11206_),
    .B(_11207_),
    .C(_11211_),
    .X(_11212_));
 sky130_fd_sc_hd__clkbuf_1 _25826_ (.A(_11212_),
    .X(_02903_));
 sky130_fd_sc_hd__and2_1 _25827_ (.A(\rvcpu.dp.pcreg.q[22] ),
    .B(_11208_),
    .X(_11213_));
 sky130_fd_sc_hd__nor2_1 _25828_ (.A(\rvcpu.dp.pcreg.q[22] ),
    .B(_11208_),
    .Y(_11214_));
 sky130_fd_sc_hd__nor2_1 _25829_ (.A(_11213_),
    .B(_11214_),
    .Y(_11215_));
 sky130_fd_sc_hd__mux2_1 _25830_ (.A0(\rvcpu.dp.plfd.PCPlus4D[22] ),
    .A1(_11215_),
    .S(_11142_),
    .X(_11216_));
 sky130_fd_sc_hd__and3_1 _25831_ (.A(_11206_),
    .B(_11207_),
    .C(_11216_),
    .X(_11217_));
 sky130_fd_sc_hd__clkbuf_1 _25832_ (.A(_11217_),
    .X(_02904_));
 sky130_fd_sc_hd__xor2_1 _25833_ (.A(\rvcpu.dp.pcreg.q[23] ),
    .B(_11213_),
    .X(_11218_));
 sky130_fd_sc_hd__mux2_1 _25834_ (.A0(\rvcpu.dp.plfd.PCPlus4D[23] ),
    .A1(_11218_),
    .S(_11142_),
    .X(_11219_));
 sky130_fd_sc_hd__and3_1 _25835_ (.A(_11206_),
    .B(_11207_),
    .C(_11219_),
    .X(_11220_));
 sky130_fd_sc_hd__clkbuf_1 _25836_ (.A(_11220_),
    .X(_02905_));
 sky130_fd_sc_hd__and3_1 _25837_ (.A(\rvcpu.dp.pcreg.q[24] ),
    .B(\rvcpu.dp.pcreg.q[23] ),
    .C(_11213_),
    .X(_11221_));
 sky130_fd_sc_hd__a21oi_1 _25838_ (.A1(\rvcpu.dp.pcreg.q[23] ),
    .A2(_11213_),
    .B1(\rvcpu.dp.pcreg.q[24] ),
    .Y(_11222_));
 sky130_fd_sc_hd__nor2_1 _25839_ (.A(_11221_),
    .B(_11222_),
    .Y(_11223_));
 sky130_fd_sc_hd__mux2_1 _25840_ (.A0(\rvcpu.dp.plfd.PCPlus4D[24] ),
    .A1(_11223_),
    .S(_11142_),
    .X(_11224_));
 sky130_fd_sc_hd__and3_1 _25841_ (.A(_11206_),
    .B(_11207_),
    .C(_11224_),
    .X(_11225_));
 sky130_fd_sc_hd__clkbuf_1 _25842_ (.A(_11225_),
    .X(_02906_));
 sky130_fd_sc_hd__and2_1 _25843_ (.A(\rvcpu.dp.pcreg.q[25] ),
    .B(_11221_),
    .X(_11226_));
 sky130_fd_sc_hd__nor2_1 _25844_ (.A(\rvcpu.dp.pcreg.q[25] ),
    .B(_11221_),
    .Y(_11227_));
 sky130_fd_sc_hd__nor2_1 _25845_ (.A(_11226_),
    .B(_11227_),
    .Y(_11228_));
 sky130_fd_sc_hd__mux2_1 _25846_ (.A0(\rvcpu.dp.plfd.PCPlus4D[25] ),
    .A1(_11228_),
    .S(_11142_),
    .X(_11229_));
 sky130_fd_sc_hd__and3_1 _25847_ (.A(_11206_),
    .B(_11207_),
    .C(_11229_),
    .X(_11230_));
 sky130_fd_sc_hd__clkbuf_1 _25848_ (.A(_11230_),
    .X(_02907_));
 sky130_fd_sc_hd__xor2_1 _25849_ (.A(\rvcpu.dp.pcreg.q[26] ),
    .B(_11226_),
    .X(_11231_));
 sky130_fd_sc_hd__mux2_1 _25850_ (.A0(\rvcpu.dp.plfd.PCPlus4D[26] ),
    .A1(_11231_),
    .S(_11142_),
    .X(_11232_));
 sky130_fd_sc_hd__and3_1 _25851_ (.A(_11206_),
    .B(_11207_),
    .C(_11232_),
    .X(_11233_));
 sky130_fd_sc_hd__clkbuf_1 _25852_ (.A(_11233_),
    .X(_02908_));
 sky130_fd_sc_hd__and3_1 _25853_ (.A(\rvcpu.dp.pcreg.q[27] ),
    .B(\rvcpu.dp.pcreg.q[26] ),
    .C(_11226_),
    .X(_11234_));
 sky130_fd_sc_hd__a21oi_1 _25854_ (.A1(\rvcpu.dp.pcreg.q[26] ),
    .A2(_11226_),
    .B1(\rvcpu.dp.pcreg.q[27] ),
    .Y(_11235_));
 sky130_fd_sc_hd__nor2_1 _25855_ (.A(_11234_),
    .B(_11235_),
    .Y(_11236_));
 sky130_fd_sc_hd__mux2_1 _25856_ (.A0(\rvcpu.dp.plfd.PCPlus4D[27] ),
    .A1(_11236_),
    .S(_08598_),
    .X(_11237_));
 sky130_fd_sc_hd__and3_1 _25857_ (.A(_11206_),
    .B(_11207_),
    .C(_11237_),
    .X(_11238_));
 sky130_fd_sc_hd__clkbuf_1 _25858_ (.A(_11238_),
    .X(_02909_));
 sky130_fd_sc_hd__and2_1 _25859_ (.A(\rvcpu.dp.pcreg.q[28] ),
    .B(_11234_),
    .X(_11239_));
 sky130_fd_sc_hd__nor2_1 _25860_ (.A(\rvcpu.dp.pcreg.q[28] ),
    .B(_11234_),
    .Y(_11240_));
 sky130_fd_sc_hd__nor2_1 _25861_ (.A(_11239_),
    .B(_11240_),
    .Y(_11241_));
 sky130_fd_sc_hd__mux2_1 _25862_ (.A0(\rvcpu.dp.plfd.PCPlus4D[28] ),
    .A1(_11241_),
    .S(_08598_),
    .X(_11242_));
 sky130_fd_sc_hd__and3_1 _25863_ (.A(_11206_),
    .B(_11207_),
    .C(_11242_),
    .X(_11243_));
 sky130_fd_sc_hd__clkbuf_1 _25864_ (.A(_11243_),
    .X(_02910_));
 sky130_fd_sc_hd__xor2_1 _25865_ (.A(\rvcpu.dp.pcreg.q[29] ),
    .B(_11239_),
    .X(_11244_));
 sky130_fd_sc_hd__mux2_1 _25866_ (.A0(\rvcpu.dp.plfd.PCPlus4D[29] ),
    .A1(_11244_),
    .S(_08598_),
    .X(_11245_));
 sky130_fd_sc_hd__and3_1 _25867_ (.A(_11206_),
    .B(_11207_),
    .C(_11245_),
    .X(_11246_));
 sky130_fd_sc_hd__clkbuf_1 _25868_ (.A(_11246_),
    .X(_02911_));
 sky130_fd_sc_hd__and3_1 _25869_ (.A(\rvcpu.dp.pcreg.q[30] ),
    .B(\rvcpu.dp.pcreg.q[29] ),
    .C(_11239_),
    .X(_11247_));
 sky130_fd_sc_hd__a21oi_1 _25870_ (.A1(\rvcpu.dp.pcreg.q[29] ),
    .A2(_11239_),
    .B1(\rvcpu.dp.pcreg.q[30] ),
    .Y(_11248_));
 sky130_fd_sc_hd__nor2_1 _25871_ (.A(_11247_),
    .B(_11248_),
    .Y(_11249_));
 sky130_fd_sc_hd__mux2_1 _25872_ (.A0(\rvcpu.dp.plfd.PCPlus4D[30] ),
    .A1(_11249_),
    .S(_08598_),
    .X(_11250_));
 sky130_fd_sc_hd__and3_1 _25873_ (.A(_11206_),
    .B(_11207_),
    .C(_11250_),
    .X(_11251_));
 sky130_fd_sc_hd__clkbuf_1 _25874_ (.A(_11251_),
    .X(_02912_));
 sky130_fd_sc_hd__inv_2 _25875_ (.A(\rvcpu.dp.pcreg.q[31] ),
    .Y(_11252_));
 sky130_fd_sc_hd__xnor2_1 _25876_ (.A(_11252_),
    .B(_11247_),
    .Y(_11253_));
 sky130_fd_sc_hd__mux2_1 _25877_ (.A0(\rvcpu.dp.plfd.PCPlus4D[31] ),
    .A1(_11253_),
    .S(_08598_),
    .X(_11254_));
 sky130_fd_sc_hd__and3_1 _25878_ (.A(_08620_),
    .B(_08621_),
    .C(_11254_),
    .X(_11255_));
 sky130_fd_sc_hd__clkbuf_1 _25879_ (.A(_11255_),
    .X(_02913_));
 sky130_fd_sc_hd__clkbuf_4 _25880_ (.A(_11153_),
    .X(_11256_));
 sky130_fd_sc_hd__or2_1 _25881_ (.A(\rvcpu.dp.plfd.PCD[0] ),
    .B(_11143_),
    .X(_11257_));
 sky130_fd_sc_hd__o211a_1 _25882_ (.A1(\rvcpu.dp.pcreg.q[0] ),
    .A2(_11256_),
    .B1(_11177_),
    .C1(_11257_),
    .X(_02914_));
 sky130_fd_sc_hd__buf_2 _25883_ (.A(_11146_),
    .X(_11258_));
 sky130_fd_sc_hd__or2_1 _25884_ (.A(\rvcpu.dp.plfd.PCD[1] ),
    .B(_11143_),
    .X(_11259_));
 sky130_fd_sc_hd__o211a_1 _25885_ (.A1(\rvcpu.dp.pcreg.q[1] ),
    .A2(_11256_),
    .B1(_11258_),
    .C1(_11259_),
    .X(_02915_));
 sky130_fd_sc_hd__nand2_1 _25886_ (.A(\rvcpu.dp.plfd.PCD[2] ),
    .B(_11153_),
    .Y(_11260_));
 sky130_fd_sc_hd__nand2_1 _25887_ (.A(_08620_),
    .B(_08621_),
    .Y(_11261_));
 sky130_fd_sc_hd__a21oi_1 _25888_ (.A1(_11148_),
    .A2(_11260_),
    .B1(_11261_),
    .Y(_02916_));
 sky130_fd_sc_hd__or2_1 _25889_ (.A(\rvcpu.dp.plfd.PCD[3] ),
    .B(_11143_),
    .X(_11262_));
 sky130_fd_sc_hd__o211a_1 _25890_ (.A1(_13665_),
    .A2(_11256_),
    .B1(_11258_),
    .C1(_11262_),
    .X(_02917_));
 sky130_fd_sc_hd__buf_2 _25891_ (.A(_11142_),
    .X(_11263_));
 sky130_fd_sc_hd__or2_1 _25892_ (.A(\rvcpu.dp.plfd.PCD[4] ),
    .B(_11263_),
    .X(_11264_));
 sky130_fd_sc_hd__o211a_1 _25893_ (.A1(_13387_),
    .A2(_11256_),
    .B1(_11258_),
    .C1(_11264_),
    .X(_02918_));
 sky130_fd_sc_hd__or2_1 _25894_ (.A(\rvcpu.dp.plfd.PCD[5] ),
    .B(_11263_),
    .X(_11265_));
 sky130_fd_sc_hd__o211a_1 _25895_ (.A1(_13682_),
    .A2(_11256_),
    .B1(_11258_),
    .C1(_11265_),
    .X(_02919_));
 sky130_fd_sc_hd__or2_1 _25896_ (.A(\rvcpu.dp.plfd.PCD[6] ),
    .B(_11263_),
    .X(_11266_));
 sky130_fd_sc_hd__o211a_1 _25897_ (.A1(_13823_),
    .A2(_11256_),
    .B1(_11258_),
    .C1(_11266_),
    .X(_02920_));
 sky130_fd_sc_hd__or2_1 _25898_ (.A(\rvcpu.dp.plfd.PCD[7] ),
    .B(_11263_),
    .X(_11267_));
 sky130_fd_sc_hd__o211a_1 _25899_ (.A1(_13706_),
    .A2(_11256_),
    .B1(_11258_),
    .C1(_11267_),
    .X(_02921_));
 sky130_fd_sc_hd__clkbuf_4 _25900_ (.A(_11155_),
    .X(_11268_));
 sky130_fd_sc_hd__nand2_1 _25901_ (.A(_13368_),
    .B(_11268_),
    .Y(_11269_));
 sky130_fd_sc_hd__o211a_1 _25902_ (.A1(\rvcpu.dp.plfd.PCD[8] ),
    .A2(_11181_),
    .B1(_11258_),
    .C1(_11269_),
    .X(_02922_));
 sky130_fd_sc_hd__nand2_1 _25903_ (.A(_13539_),
    .B(_11268_),
    .Y(_11270_));
 sky130_fd_sc_hd__o211a_1 _25904_ (.A1(\rvcpu.dp.plfd.PCD[9] ),
    .A2(_11181_),
    .B1(_11258_),
    .C1(_11270_),
    .X(_02923_));
 sky130_fd_sc_hd__or2_1 _25905_ (.A(\rvcpu.dp.plfd.PCD[10] ),
    .B(_11263_),
    .X(_11271_));
 sky130_fd_sc_hd__o211a_1 _25906_ (.A1(\rvcpu.dp.pcreg.q[10] ),
    .A2(_11256_),
    .B1(_11258_),
    .C1(_11271_),
    .X(_02924_));
 sky130_fd_sc_hd__or2_1 _25907_ (.A(\rvcpu.dp.plfd.PCD[11] ),
    .B(_11263_),
    .X(_11272_));
 sky130_fd_sc_hd__o211a_1 _25908_ (.A1(\rvcpu.dp.pcreg.q[11] ),
    .A2(_11256_),
    .B1(_11258_),
    .C1(_11272_),
    .X(_02925_));
 sky130_fd_sc_hd__buf_2 _25909_ (.A(_11146_),
    .X(_11273_));
 sky130_fd_sc_hd__or2_1 _25910_ (.A(\rvcpu.dp.plfd.PCD[12] ),
    .B(_11263_),
    .X(_11274_));
 sky130_fd_sc_hd__o211a_1 _25911_ (.A1(\rvcpu.dp.pcreg.q[12] ),
    .A2(_11256_),
    .B1(_11273_),
    .C1(_11274_),
    .X(_02926_));
 sky130_fd_sc_hd__buf_2 _25912_ (.A(_11153_),
    .X(_11275_));
 sky130_fd_sc_hd__or2_1 _25913_ (.A(\rvcpu.dp.plfd.PCD[13] ),
    .B(_11263_),
    .X(_11276_));
 sky130_fd_sc_hd__o211a_1 _25914_ (.A1(\rvcpu.dp.pcreg.q[13] ),
    .A2(_11275_),
    .B1(_11273_),
    .C1(_11276_),
    .X(_02927_));
 sky130_fd_sc_hd__or2_1 _25915_ (.A(\rvcpu.dp.plfd.PCD[14] ),
    .B(_11263_),
    .X(_11277_));
 sky130_fd_sc_hd__o211a_1 _25916_ (.A1(\rvcpu.dp.pcreg.q[14] ),
    .A2(_11275_),
    .B1(_11273_),
    .C1(_11277_),
    .X(_02928_));
 sky130_fd_sc_hd__or2_1 _25917_ (.A(\rvcpu.dp.plfd.PCD[15] ),
    .B(_11263_),
    .X(_11278_));
 sky130_fd_sc_hd__o211a_1 _25918_ (.A1(\rvcpu.dp.pcreg.q[15] ),
    .A2(_11275_),
    .B1(_11273_),
    .C1(_11278_),
    .X(_02929_));
 sky130_fd_sc_hd__clkbuf_2 _25919_ (.A(_11142_),
    .X(_11279_));
 sky130_fd_sc_hd__or2_1 _25920_ (.A(\rvcpu.dp.plfd.PCD[16] ),
    .B(_11279_),
    .X(_11280_));
 sky130_fd_sc_hd__o211a_1 _25921_ (.A1(\rvcpu.dp.pcreg.q[16] ),
    .A2(_11275_),
    .B1(_11273_),
    .C1(_11280_),
    .X(_02930_));
 sky130_fd_sc_hd__or2_1 _25922_ (.A(\rvcpu.dp.plfd.PCD[17] ),
    .B(_11279_),
    .X(_11281_));
 sky130_fd_sc_hd__o211a_1 _25923_ (.A1(\rvcpu.dp.pcreg.q[17] ),
    .A2(_11275_),
    .B1(_11273_),
    .C1(_11281_),
    .X(_02931_));
 sky130_fd_sc_hd__or2_1 _25924_ (.A(\rvcpu.dp.plfd.PCD[18] ),
    .B(_11279_),
    .X(_11282_));
 sky130_fd_sc_hd__o211a_1 _25925_ (.A1(\rvcpu.dp.pcreg.q[18] ),
    .A2(_11275_),
    .B1(_11273_),
    .C1(_11282_),
    .X(_02932_));
 sky130_fd_sc_hd__or2_1 _25926_ (.A(\rvcpu.dp.plfd.PCD[19] ),
    .B(_11279_),
    .X(_11283_));
 sky130_fd_sc_hd__o211a_1 _25927_ (.A1(\rvcpu.dp.pcreg.q[19] ),
    .A2(_11275_),
    .B1(_11273_),
    .C1(_11283_),
    .X(_02933_));
 sky130_fd_sc_hd__or2_1 _25928_ (.A(\rvcpu.dp.plfd.PCD[20] ),
    .B(_11279_),
    .X(_11284_));
 sky130_fd_sc_hd__o211a_1 _25929_ (.A1(\rvcpu.dp.pcreg.q[20] ),
    .A2(_11275_),
    .B1(_11273_),
    .C1(_11284_),
    .X(_02934_));
 sky130_fd_sc_hd__or2_1 _25930_ (.A(\rvcpu.dp.plfd.PCD[21] ),
    .B(_11279_),
    .X(_11285_));
 sky130_fd_sc_hd__o211a_1 _25931_ (.A1(\rvcpu.dp.pcreg.q[21] ),
    .A2(_11275_),
    .B1(_11273_),
    .C1(_11285_),
    .X(_02935_));
 sky130_fd_sc_hd__buf_2 _25932_ (.A(_11146_),
    .X(_11286_));
 sky130_fd_sc_hd__or2_1 _25933_ (.A(\rvcpu.dp.plfd.PCD[22] ),
    .B(_11279_),
    .X(_11287_));
 sky130_fd_sc_hd__o211a_1 _25934_ (.A1(\rvcpu.dp.pcreg.q[22] ),
    .A2(_11275_),
    .B1(_11286_),
    .C1(_11287_),
    .X(_02936_));
 sky130_fd_sc_hd__buf_2 _25935_ (.A(_11157_),
    .X(_11288_));
 sky130_fd_sc_hd__clkbuf_2 _25936_ (.A(_11288_),
    .X(_11289_));
 sky130_fd_sc_hd__clkbuf_4 _25937_ (.A(_11289_),
    .X(_11290_));
 sky130_fd_sc_hd__or2_1 _25938_ (.A(\rvcpu.dp.plfd.PCD[23] ),
    .B(_11279_),
    .X(_11291_));
 sky130_fd_sc_hd__o211a_1 _25939_ (.A1(\rvcpu.dp.pcreg.q[23] ),
    .A2(_11290_),
    .B1(_11286_),
    .C1(_11291_),
    .X(_02937_));
 sky130_fd_sc_hd__or2_1 _25940_ (.A(\rvcpu.dp.plfd.PCD[24] ),
    .B(_11279_),
    .X(_11292_));
 sky130_fd_sc_hd__o211a_1 _25941_ (.A1(\rvcpu.dp.pcreg.q[24] ),
    .A2(_11290_),
    .B1(_11286_),
    .C1(_11292_),
    .X(_02938_));
 sky130_fd_sc_hd__or2_1 _25942_ (.A(\rvcpu.dp.plfd.PCD[25] ),
    .B(_11279_),
    .X(_11293_));
 sky130_fd_sc_hd__o211a_1 _25943_ (.A1(\rvcpu.dp.pcreg.q[25] ),
    .A2(_11290_),
    .B1(_11286_),
    .C1(_11293_),
    .X(_02939_));
 sky130_fd_sc_hd__or2_1 _25944_ (.A(\rvcpu.dp.plfd.PCD[26] ),
    .B(_11155_),
    .X(_11294_));
 sky130_fd_sc_hd__o211a_1 _25945_ (.A1(\rvcpu.dp.pcreg.q[26] ),
    .A2(_11290_),
    .B1(_11286_),
    .C1(_11294_),
    .X(_02940_));
 sky130_fd_sc_hd__or2_1 _25946_ (.A(\rvcpu.dp.plfd.PCD[27] ),
    .B(_11155_),
    .X(_11295_));
 sky130_fd_sc_hd__o211a_1 _25947_ (.A1(\rvcpu.dp.pcreg.q[27] ),
    .A2(_11290_),
    .B1(_11286_),
    .C1(_11295_),
    .X(_02941_));
 sky130_fd_sc_hd__or2_1 _25948_ (.A(\rvcpu.dp.plfd.PCD[28] ),
    .B(_11155_),
    .X(_11296_));
 sky130_fd_sc_hd__o211a_1 _25949_ (.A1(\rvcpu.dp.pcreg.q[28] ),
    .A2(_11290_),
    .B1(_11286_),
    .C1(_11296_),
    .X(_02942_));
 sky130_fd_sc_hd__or2_1 _25950_ (.A(\rvcpu.dp.plfd.PCD[29] ),
    .B(_11155_),
    .X(_11297_));
 sky130_fd_sc_hd__o211a_1 _25951_ (.A1(\rvcpu.dp.pcreg.q[29] ),
    .A2(_11290_),
    .B1(_11286_),
    .C1(_11297_),
    .X(_02943_));
 sky130_fd_sc_hd__or2_1 _25952_ (.A(\rvcpu.dp.plfd.PCD[30] ),
    .B(_11155_),
    .X(_11298_));
 sky130_fd_sc_hd__o211a_1 _25953_ (.A1(\rvcpu.dp.pcreg.q[30] ),
    .A2(_11290_),
    .B1(_11286_),
    .C1(_11298_),
    .X(_02944_));
 sky130_fd_sc_hd__or2_1 _25954_ (.A(\rvcpu.dp.plfd.PCD[31] ),
    .B(_11155_),
    .X(_11299_));
 sky130_fd_sc_hd__o211a_1 _25955_ (.A1(\rvcpu.dp.pcreg.q[31] ),
    .A2(_11290_),
    .B1(_11286_),
    .C1(_11299_),
    .X(_02945_));
 sky130_fd_sc_hd__buf_2 _25956_ (.A(_11146_),
    .X(_11300_));
 sky130_fd_sc_hd__or2_1 _25957_ (.A(\rvcpu.dp.plfd.InstrD[0] ),
    .B(_11155_),
    .X(_11301_));
 sky130_fd_sc_hd__o211a_1 _25958_ (.A1(net13),
    .A2(_11290_),
    .B1(_11300_),
    .C1(_11301_),
    .X(_02946_));
 sky130_fd_sc_hd__buf_2 _25959_ (.A(_11143_),
    .X(_11302_));
 sky130_fd_sc_hd__or2_1 _25960_ (.A(net24),
    .B(_11289_),
    .X(_11303_));
 sky130_fd_sc_hd__o211a_1 _25961_ (.A1(\rvcpu.dp.plfd.InstrD[2] ),
    .A2(_11302_),
    .B1(_11300_),
    .C1(_11303_),
    .X(_02947_));
 sky130_fd_sc_hd__or2_1 _25962_ (.A(net27),
    .B(_11289_),
    .X(_11304_));
 sky130_fd_sc_hd__o211a_1 _25963_ (.A1(\rvcpu.dp.plfd.InstrD[3] ),
    .A2(_11302_),
    .B1(_11300_),
    .C1(_11304_),
    .X(_02948_));
 sky130_fd_sc_hd__or2_1 _25964_ (.A(\rvcpu.dp.plfd.InstrD[4] ),
    .B(_11155_),
    .X(_11305_));
 sky130_fd_sc_hd__o211a_1 _25965_ (.A1(net28),
    .A2(_11153_),
    .B1(_11300_),
    .C1(_11305_),
    .X(_02949_));
 sky130_fd_sc_hd__or2_1 _25966_ (.A(net29),
    .B(_11289_),
    .X(_11306_));
 sky130_fd_sc_hd__o211a_1 _25967_ (.A1(\rvcpu.c.ad.opb5 ),
    .A2(_11302_),
    .B1(_11300_),
    .C1(_11306_),
    .X(_02950_));
 sky130_fd_sc_hd__or2_1 _25968_ (.A(net30),
    .B(_11289_),
    .X(_11307_));
 sky130_fd_sc_hd__o211a_1 _25969_ (.A1(\rvcpu.dp.plfd.InstrD[6] ),
    .A2(_11302_),
    .B1(_11300_),
    .C1(_11307_),
    .X(_02951_));
 sky130_fd_sc_hd__or2_1 _25970_ (.A(net31),
    .B(_11289_),
    .X(_11308_));
 sky130_fd_sc_hd__o211a_1 _25971_ (.A1(\rvcpu.dp.plfd.InstrD[7] ),
    .A2(_11302_),
    .B1(_11300_),
    .C1(_11308_),
    .X(_02952_));
 sky130_fd_sc_hd__nand2_1 _25972_ (.A(_14002_),
    .B(_11268_),
    .Y(_11309_));
 sky130_fd_sc_hd__o211a_1 _25973_ (.A1(\rvcpu.dp.plfd.InstrD[8] ),
    .A2(_11302_),
    .B1(_11300_),
    .C1(_11309_),
    .X(_02953_));
 sky130_fd_sc_hd__or2_1 _25974_ (.A(net33),
    .B(_11289_),
    .X(_11310_));
 sky130_fd_sc_hd__o211a_1 _25975_ (.A1(\rvcpu.dp.plfd.InstrD[9] ),
    .A2(_11302_),
    .B1(_11300_),
    .C1(_11310_),
    .X(_02954_));
 sky130_fd_sc_hd__or2_1 _25976_ (.A(net3),
    .B(_11289_),
    .X(_11311_));
 sky130_fd_sc_hd__o211a_1 _25977_ (.A1(\rvcpu.dp.plfd.InstrD[10] ),
    .A2(_11302_),
    .B1(_11300_),
    .C1(_11311_),
    .X(_02955_));
 sky130_fd_sc_hd__buf_2 _25978_ (.A(_11146_),
    .X(_11312_));
 sky130_fd_sc_hd__nand2_1 _25979_ (.A(_13932_),
    .B(_11268_),
    .Y(_11313_));
 sky130_fd_sc_hd__o211a_1 _25980_ (.A1(\rvcpu.dp.plfd.InstrD[11] ),
    .A2(_11302_),
    .B1(_11312_),
    .C1(_11313_),
    .X(_02956_));
 sky130_fd_sc_hd__or2_1 _25981_ (.A(net5),
    .B(_11289_),
    .X(_11314_));
 sky130_fd_sc_hd__o211a_1 _25982_ (.A1(\rvcpu.dp.plfd.InstrD[12] ),
    .A2(_11302_),
    .B1(_11312_),
    .C1(_11314_),
    .X(_02957_));
 sky130_fd_sc_hd__buf_2 _25983_ (.A(_11143_),
    .X(_11315_));
 sky130_fd_sc_hd__nand2_1 _25984_ (.A(_13903_),
    .B(_11268_),
    .Y(_11316_));
 sky130_fd_sc_hd__o211a_1 _25985_ (.A1(\rvcpu.dp.plfd.InstrD[13] ),
    .A2(_11315_),
    .B1(_11312_),
    .C1(_11316_),
    .X(_02958_));
 sky130_fd_sc_hd__clkbuf_2 _25986_ (.A(_11157_),
    .X(_11317_));
 sky130_fd_sc_hd__or2_1 _25987_ (.A(net7),
    .B(_11317_),
    .X(_11318_));
 sky130_fd_sc_hd__o211a_1 _25988_ (.A1(\rvcpu.dp.plfd.InstrD[14] ),
    .A2(_11315_),
    .B1(_11312_),
    .C1(_11318_),
    .X(_02959_));
 sky130_fd_sc_hd__or2_1 _25989_ (.A(net8),
    .B(_11317_),
    .X(_11319_));
 sky130_fd_sc_hd__o211a_1 _25990_ (.A1(_08567_),
    .A2(_11315_),
    .B1(_11312_),
    .C1(_11319_),
    .X(_02960_));
 sky130_fd_sc_hd__or2_1 _25991_ (.A(net9),
    .B(_11317_),
    .X(_11320_));
 sky130_fd_sc_hd__o211a_1 _25992_ (.A1(_08570_),
    .A2(_11315_),
    .B1(_11312_),
    .C1(_11320_),
    .X(_02961_));
 sky130_fd_sc_hd__or2_1 _25993_ (.A(net10),
    .B(_11317_),
    .X(_11321_));
 sky130_fd_sc_hd__o211a_1 _25994_ (.A1(_08572_),
    .A2(_11315_),
    .B1(_11312_),
    .C1(_11321_),
    .X(_02962_));
 sky130_fd_sc_hd__or2_1 _25995_ (.A(net11),
    .B(_11317_),
    .X(_11322_));
 sky130_fd_sc_hd__o211a_1 _25996_ (.A1(_08513_),
    .A2(_11315_),
    .B1(_11312_),
    .C1(_11322_),
    .X(_02963_));
 sky130_fd_sc_hd__or2_1 _25997_ (.A(net12),
    .B(_11317_),
    .X(_11323_));
 sky130_fd_sc_hd__o211a_1 _25998_ (.A1(\rvcpu.dp.plfd.InstrD[19] ),
    .A2(_11315_),
    .B1(_11312_),
    .C1(_11323_),
    .X(_02964_));
 sky130_fd_sc_hd__or2_1 _25999_ (.A(net14),
    .B(_11317_),
    .X(_11324_));
 sky130_fd_sc_hd__o211a_1 _26000_ (.A1(_09478_),
    .A2(_11315_),
    .B1(_11312_),
    .C1(_11324_),
    .X(_02965_));
 sky130_fd_sc_hd__clkbuf_4 _26001_ (.A(_11146_),
    .X(_11325_));
 sky130_fd_sc_hd__or2_1 _26002_ (.A(net15),
    .B(_11317_),
    .X(_11326_));
 sky130_fd_sc_hd__o211a_1 _26003_ (.A1(_09479_),
    .A2(_11315_),
    .B1(_11325_),
    .C1(_11326_),
    .X(_02966_));
 sky130_fd_sc_hd__nand2_1 _26004_ (.A(_09476_),
    .B(_11153_),
    .Y(_11327_));
 sky130_fd_sc_hd__o211a_1 _26005_ (.A1(net16),
    .A2(_11153_),
    .B1(_11325_),
    .C1(_11327_),
    .X(_02967_));
 sky130_fd_sc_hd__or2_1 _26006_ (.A(net17),
    .B(_11317_),
    .X(_11328_));
 sky130_fd_sc_hd__o211a_1 _26007_ (.A1(_09457_),
    .A2(_11315_),
    .B1(_11325_),
    .C1(_11328_),
    .X(_02968_));
 sky130_fd_sc_hd__clkbuf_4 _26008_ (.A(_11143_),
    .X(_11329_));
 sky130_fd_sc_hd__or2_1 _26009_ (.A(net18),
    .B(_11317_),
    .X(_11330_));
 sky130_fd_sc_hd__o211a_1 _26010_ (.A1(\rvcpu.dp.plfd.InstrD[24] ),
    .A2(_11329_),
    .B1(_11325_),
    .C1(_11330_),
    .X(_02969_));
 sky130_fd_sc_hd__or2_1 _26011_ (.A(net19),
    .B(_11152_),
    .X(_11331_));
 sky130_fd_sc_hd__o211a_1 _26012_ (.A1(\rvcpu.dp.plfd.InstrD[25] ),
    .A2(_11329_),
    .B1(_11325_),
    .C1(_11331_),
    .X(_02970_));
 sky130_fd_sc_hd__or2_1 _26013_ (.A(net20),
    .B(_11152_),
    .X(_11332_));
 sky130_fd_sc_hd__o211a_1 _26014_ (.A1(\rvcpu.dp.plfd.InstrD[26] ),
    .A2(_11329_),
    .B1(_11325_),
    .C1(_11332_),
    .X(_02971_));
 sky130_fd_sc_hd__or2_1 _26015_ (.A(net21),
    .B(_11152_),
    .X(_11333_));
 sky130_fd_sc_hd__o211a_1 _26016_ (.A1(\rvcpu.dp.plfd.InstrD[27] ),
    .A2(_11329_),
    .B1(_11325_),
    .C1(_11333_),
    .X(_02972_));
 sky130_fd_sc_hd__or2_1 _26017_ (.A(net22),
    .B(_11152_),
    .X(_11334_));
 sky130_fd_sc_hd__o211a_1 _26018_ (.A1(\rvcpu.dp.plfd.InstrD[28] ),
    .A2(_11329_),
    .B1(_11325_),
    .C1(_11334_),
    .X(_02973_));
 sky130_fd_sc_hd__or2_1 _26019_ (.A(net23),
    .B(_11152_),
    .X(_11335_));
 sky130_fd_sc_hd__o211a_1 _26020_ (.A1(\rvcpu.dp.plfd.InstrD[29] ),
    .A2(_11329_),
    .B1(_11325_),
    .C1(_11335_),
    .X(_02974_));
 sky130_fd_sc_hd__or2_1 _26021_ (.A(net25),
    .B(_11152_),
    .X(_11336_));
 sky130_fd_sc_hd__o211a_1 _26022_ (.A1(\rvcpu.c.ad.funct7b5 ),
    .A2(_11329_),
    .B1(_11325_),
    .C1(_11336_),
    .X(_02975_));
 sky130_fd_sc_hd__or2_1 _26023_ (.A(net26),
    .B(_11152_),
    .X(_11337_));
 sky130_fd_sc_hd__o211a_1 _26024_ (.A1(\rvcpu.dp.plfd.InstrD[31] ),
    .A2(_11329_),
    .B1(_11146_),
    .C1(_11337_),
    .X(_02976_));
 sky130_fd_sc_hd__or2_1 _26025_ (.A(_11109_),
    .B(_10980_),
    .X(_11338_));
 sky130_fd_sc_hd__clkbuf_2 _26026_ (.A(_11338_),
    .X(_11339_));
 sky130_fd_sc_hd__nor2_1 _26027_ (.A(_11109_),
    .B(_10980_),
    .Y(_11340_));
 sky130_fd_sc_hd__and2_1 _26028_ (.A(_11078_),
    .B(_11340_),
    .X(_11341_));
 sky130_fd_sc_hd__a31o_1 _26029_ (.A1(_11121_),
    .A2(\datamem.data_ram[24][0] ),
    .A3(_11339_),
    .B1(_11341_),
    .X(_02977_));
 sky130_fd_sc_hd__and2_1 _26030_ (.A(_11081_),
    .B(_11340_),
    .X(_11342_));
 sky130_fd_sc_hd__a31o_1 _26031_ (.A1(_11121_),
    .A2(\datamem.data_ram[24][1] ),
    .A3(_11339_),
    .B1(_11342_),
    .X(_02978_));
 sky130_fd_sc_hd__and2_1 _26032_ (.A(_11083_),
    .B(_11340_),
    .X(_11343_));
 sky130_fd_sc_hd__a31o_1 _26033_ (.A1(_11121_),
    .A2(\datamem.data_ram[24][2] ),
    .A3(_11339_),
    .B1(_11343_),
    .X(_02979_));
 sky130_fd_sc_hd__and2_1 _26034_ (.A(_11086_),
    .B(_11340_),
    .X(_11344_));
 sky130_fd_sc_hd__a31o_1 _26035_ (.A1(_11121_),
    .A2(\datamem.data_ram[24][3] ),
    .A3(_11339_),
    .B1(_11344_),
    .X(_02980_));
 sky130_fd_sc_hd__and2_1 _26036_ (.A(_11047_),
    .B(_11340_),
    .X(_11345_));
 sky130_fd_sc_hd__a31o_1 _26037_ (.A1(_11121_),
    .A2(\datamem.data_ram[24][4] ),
    .A3(_11339_),
    .B1(_11345_),
    .X(_02981_));
 sky130_fd_sc_hd__and2_1 _26038_ (.A(_11089_),
    .B(_11340_),
    .X(_11346_));
 sky130_fd_sc_hd__a31o_1 _26039_ (.A1(_11121_),
    .A2(\datamem.data_ram[24][5] ),
    .A3(_11339_),
    .B1(_11346_),
    .X(_02982_));
 sky130_fd_sc_hd__and2_1 _26040_ (.A(_11091_),
    .B(_11340_),
    .X(_11347_));
 sky130_fd_sc_hd__a31o_1 _26041_ (.A1(_11121_),
    .A2(\datamem.data_ram[24][6] ),
    .A3(_11339_),
    .B1(_11347_),
    .X(_02983_));
 sky130_fd_sc_hd__and2_1 _26042_ (.A(_11064_),
    .B(_11340_),
    .X(_11348_));
 sky130_fd_sc_hd__a31o_1 _26043_ (.A1(_11121_),
    .A2(\datamem.data_ram[24][7] ),
    .A3(_11339_),
    .B1(_11348_),
    .X(_02984_));
 sky130_fd_sc_hd__or3_1 _26044_ (.A(_07203_),
    .B(_10918_),
    .C(_10897_),
    .X(_11349_));
 sky130_fd_sc_hd__clkbuf_2 _26045_ (.A(_11349_),
    .X(_11350_));
 sky130_fd_sc_hd__and3_2 _26046_ (.A(_10209_),
    .B(_10921_),
    .C(_10922_),
    .X(_11351_));
 sky130_fd_sc_hd__and2_1 _26047_ (.A(_11078_),
    .B(_11351_),
    .X(_11352_));
 sky130_fd_sc_hd__a31o_1 _26048_ (.A1(_11121_),
    .A2(\datamem.data_ram[34][0] ),
    .A3(_11350_),
    .B1(_11352_),
    .X(_02985_));
 sky130_fd_sc_hd__clkbuf_4 _26049_ (.A(_11104_),
    .X(_11353_));
 sky130_fd_sc_hd__and2_1 _26050_ (.A(_11081_),
    .B(_11351_),
    .X(_11354_));
 sky130_fd_sc_hd__a31o_1 _26051_ (.A1(_11353_),
    .A2(\datamem.data_ram[34][1] ),
    .A3(_11350_),
    .B1(_11354_),
    .X(_02986_));
 sky130_fd_sc_hd__and2_1 _26052_ (.A(_11083_),
    .B(_11351_),
    .X(_11355_));
 sky130_fd_sc_hd__a31o_1 _26053_ (.A1(_11353_),
    .A2(\datamem.data_ram[34][2] ),
    .A3(_11350_),
    .B1(_11355_),
    .X(_02987_));
 sky130_fd_sc_hd__and2_1 _26054_ (.A(_11086_),
    .B(_11351_),
    .X(_11356_));
 sky130_fd_sc_hd__a31o_1 _26055_ (.A1(_11353_),
    .A2(\datamem.data_ram[34][3] ),
    .A3(_11350_),
    .B1(_11356_),
    .X(_02988_));
 sky130_fd_sc_hd__and2_1 _26056_ (.A(_11047_),
    .B(_11351_),
    .X(_11357_));
 sky130_fd_sc_hd__a31o_1 _26057_ (.A1(_11353_),
    .A2(\datamem.data_ram[34][4] ),
    .A3(_11350_),
    .B1(_11357_),
    .X(_02989_));
 sky130_fd_sc_hd__and2_1 _26058_ (.A(_11089_),
    .B(_11351_),
    .X(_11358_));
 sky130_fd_sc_hd__a31o_1 _26059_ (.A1(_11353_),
    .A2(\datamem.data_ram[34][5] ),
    .A3(_11350_),
    .B1(_11358_),
    .X(_02990_));
 sky130_fd_sc_hd__and2_1 _26060_ (.A(_11091_),
    .B(_11351_),
    .X(_11359_));
 sky130_fd_sc_hd__a31o_1 _26061_ (.A1(_11353_),
    .A2(\datamem.data_ram[34][6] ),
    .A3(_11350_),
    .B1(_11359_),
    .X(_02991_));
 sky130_fd_sc_hd__and2_1 _26062_ (.A(_11064_),
    .B(_11351_),
    .X(_11360_));
 sky130_fd_sc_hd__a31o_1 _26063_ (.A1(_11353_),
    .A2(\datamem.data_ram[34][7] ),
    .A3(_11350_),
    .B1(_11360_),
    .X(_02992_));
 sky130_fd_sc_hd__and2_1 _26064_ (.A(\rvcpu.c.ad.opb5 ),
    .B(_06572_),
    .X(_11361_));
 sky130_fd_sc_hd__clkbuf_2 _26065_ (.A(_08622_),
    .X(_11362_));
 sky130_fd_sc_hd__and3b_1 _26066_ (.A_N(\rvcpu.dp.plfd.InstrD[6] ),
    .B(_11361_),
    .C(_11362_),
    .X(_11363_));
 sky130_fd_sc_hd__buf_2 _26067_ (.A(_11363_),
    .X(_02993_));
 sky130_fd_sc_hd__and2_1 _26068_ (.A(\rvcpu.dp.plfd.InstrD[12] ),
    .B(_08622_),
    .X(_11364_));
 sky130_fd_sc_hd__buf_1 _26069_ (.A(_11364_),
    .X(_03029_));
 sky130_fd_sc_hd__and4_1 _26070_ (.A(_06568_),
    .B(\rvcpu.dp.plfd.InstrD[13] ),
    .C(_06567_),
    .D(_03029_),
    .X(_11365_));
 sky130_fd_sc_hd__clkbuf_1 _26071_ (.A(_11365_),
    .X(_02994_));
 sky130_fd_sc_hd__and3b_1 _26072_ (.A_N(\rvcpu.dp.plfd.InstrD[4] ),
    .B(\rvcpu.c.ad.opb5 ),
    .C(\rvcpu.dp.plfd.InstrD[6] ),
    .X(_11366_));
 sky130_fd_sc_hd__and4b_1 _26073_ (.A_N(\rvcpu.dp.plfd.InstrD[3] ),
    .B(\rvcpu.dp.plfd.InstrD[2] ),
    .C(\rvcpu.dp.plfd.InstrD[0] ),
    .D(_11366_),
    .X(_11367_));
 sky130_fd_sc_hd__and2_1 _26074_ (.A(_08622_),
    .B(_11367_),
    .X(_11368_));
 sky130_fd_sc_hd__clkbuf_1 _26075_ (.A(_11368_),
    .X(_02995_));
 sky130_fd_sc_hd__and4_1 _26076_ (.A(\rvcpu.dp.plfd.InstrD[3] ),
    .B(\rvcpu.dp.plfd.InstrD[2] ),
    .C(\rvcpu.dp.plfd.InstrD[0] ),
    .D(_11366_),
    .X(_11369_));
 sky130_fd_sc_hd__and2_1 _26077_ (.A(_08622_),
    .B(_11369_),
    .X(_11370_));
 sky130_fd_sc_hd__clkbuf_1 _26078_ (.A(_11370_),
    .X(_02996_));
 sky130_fd_sc_hd__clkbuf_4 _26079_ (.A(_11362_),
    .X(_11371_));
 sky130_fd_sc_hd__clkbuf_4 _26080_ (.A(_11371_),
    .X(_11372_));
 sky130_fd_sc_hd__and2_1 _26081_ (.A(_06573_),
    .B(_11372_),
    .X(_11373_));
 sky130_fd_sc_hd__clkbuf_1 _26082_ (.A(_11373_),
    .X(_02997_));
 sky130_fd_sc_hd__inv_2 _26083_ (.A(\rvcpu.c.ad.opb5 ),
    .Y(_11374_));
 sky130_fd_sc_hd__and3b_1 _26084_ (.A_N(\rvcpu.dp.plfd.InstrD[6] ),
    .B(_11374_),
    .C(_06572_),
    .X(_11375_));
 sky130_fd_sc_hd__nand2_1 _26085_ (.A(\rvcpu.dp.plfd.InstrD[2] ),
    .B(\rvcpu.dp.plfd.InstrD[0] ),
    .Y(_11376_));
 sky130_fd_sc_hd__nor4b_1 _26086_ (.A(\rvcpu.dp.plfd.InstrD[6] ),
    .B(\rvcpu.dp.plfd.InstrD[3] ),
    .C(_11376_),
    .D_N(\rvcpu.dp.plfd.InstrD[4] ),
    .Y(_11377_));
 sky130_fd_sc_hd__or2_1 _26087_ (.A(_11369_),
    .B(net116),
    .X(_11378_));
 sky130_fd_sc_hd__clkbuf_4 _26088_ (.A(_11378_),
    .X(_11379_));
 sky130_fd_sc_hd__o41a_1 _26089_ (.A1(_06567_),
    .A2(_11367_),
    .A3(_11375_),
    .A4(_11379_),
    .B1(_11372_),
    .X(_02998_));
 sky130_fd_sc_hd__and2_1 _26090_ (.A(\rvcpu.dp.plfd.PCPlus4D[2] ),
    .B(_11372_),
    .X(_11380_));
 sky130_fd_sc_hd__clkbuf_1 _26091_ (.A(_11380_),
    .X(_02999_));
 sky130_fd_sc_hd__and2_1 _26092_ (.A(\rvcpu.dp.plfd.PCPlus4D[3] ),
    .B(_11372_),
    .X(_11381_));
 sky130_fd_sc_hd__clkbuf_1 _26093_ (.A(_11381_),
    .X(_03000_));
 sky130_fd_sc_hd__and2_1 _26094_ (.A(\rvcpu.dp.plfd.PCPlus4D[4] ),
    .B(_11372_),
    .X(_11382_));
 sky130_fd_sc_hd__clkbuf_1 _26095_ (.A(_11382_),
    .X(_03001_));
 sky130_fd_sc_hd__and2_1 _26096_ (.A(\rvcpu.dp.plfd.PCPlus4D[5] ),
    .B(_11372_),
    .X(_11383_));
 sky130_fd_sc_hd__clkbuf_1 _26097_ (.A(_11383_),
    .X(_03002_));
 sky130_fd_sc_hd__and2_1 _26098_ (.A(\rvcpu.dp.plfd.PCPlus4D[6] ),
    .B(_11372_),
    .X(_11384_));
 sky130_fd_sc_hd__clkbuf_1 _26099_ (.A(_11384_),
    .X(_03003_));
 sky130_fd_sc_hd__and2_1 _26100_ (.A(\rvcpu.dp.plfd.PCPlus4D[7] ),
    .B(_11372_),
    .X(_11385_));
 sky130_fd_sc_hd__clkbuf_1 _26101_ (.A(_11385_),
    .X(_03004_));
 sky130_fd_sc_hd__buf_2 _26102_ (.A(_11371_),
    .X(_11386_));
 sky130_fd_sc_hd__and2_1 _26103_ (.A(\rvcpu.dp.plfd.PCPlus4D[8] ),
    .B(_11386_),
    .X(_11387_));
 sky130_fd_sc_hd__clkbuf_1 _26104_ (.A(_11387_),
    .X(_03005_));
 sky130_fd_sc_hd__and2_1 _26105_ (.A(\rvcpu.dp.plfd.PCPlus4D[9] ),
    .B(_11386_),
    .X(_11388_));
 sky130_fd_sc_hd__clkbuf_1 _26106_ (.A(_11388_),
    .X(_03006_));
 sky130_fd_sc_hd__and2_1 _26107_ (.A(\rvcpu.dp.plfd.PCPlus4D[10] ),
    .B(_11386_),
    .X(_11389_));
 sky130_fd_sc_hd__clkbuf_1 _26108_ (.A(_11389_),
    .X(_03007_));
 sky130_fd_sc_hd__and2_1 _26109_ (.A(\rvcpu.dp.plfd.PCPlus4D[11] ),
    .B(_11386_),
    .X(_11390_));
 sky130_fd_sc_hd__clkbuf_1 _26110_ (.A(_11390_),
    .X(_03008_));
 sky130_fd_sc_hd__and2_1 _26111_ (.A(\rvcpu.dp.plfd.PCPlus4D[12] ),
    .B(_11386_),
    .X(_11391_));
 sky130_fd_sc_hd__clkbuf_1 _26112_ (.A(_11391_),
    .X(_03009_));
 sky130_fd_sc_hd__and2_1 _26113_ (.A(\rvcpu.dp.plfd.PCPlus4D[13] ),
    .B(_11386_),
    .X(_11392_));
 sky130_fd_sc_hd__clkbuf_1 _26114_ (.A(_11392_),
    .X(_03010_));
 sky130_fd_sc_hd__and2_1 _26115_ (.A(\rvcpu.dp.plfd.PCPlus4D[14] ),
    .B(_11386_),
    .X(_11393_));
 sky130_fd_sc_hd__clkbuf_1 _26116_ (.A(_11393_),
    .X(_03011_));
 sky130_fd_sc_hd__and2_1 _26117_ (.A(\rvcpu.dp.plfd.PCPlus4D[15] ),
    .B(_11386_),
    .X(_11394_));
 sky130_fd_sc_hd__clkbuf_1 _26118_ (.A(_11394_),
    .X(_03012_));
 sky130_fd_sc_hd__and2_1 _26119_ (.A(\rvcpu.dp.plfd.PCPlus4D[16] ),
    .B(_11386_),
    .X(_11395_));
 sky130_fd_sc_hd__clkbuf_1 _26120_ (.A(_11395_),
    .X(_03013_));
 sky130_fd_sc_hd__and2_1 _26121_ (.A(\rvcpu.dp.plfd.PCPlus4D[17] ),
    .B(_11386_),
    .X(_11396_));
 sky130_fd_sc_hd__clkbuf_1 _26122_ (.A(_11396_),
    .X(_03014_));
 sky130_fd_sc_hd__clkbuf_2 _26123_ (.A(_11371_),
    .X(_11397_));
 sky130_fd_sc_hd__and2_1 _26124_ (.A(\rvcpu.dp.plfd.PCPlus4D[18] ),
    .B(_11397_),
    .X(_11398_));
 sky130_fd_sc_hd__clkbuf_1 _26125_ (.A(_11398_),
    .X(_03015_));
 sky130_fd_sc_hd__and2_1 _26126_ (.A(\rvcpu.dp.plfd.PCPlus4D[19] ),
    .B(_11397_),
    .X(_11399_));
 sky130_fd_sc_hd__clkbuf_1 _26127_ (.A(_11399_),
    .X(_03016_));
 sky130_fd_sc_hd__and2_1 _26128_ (.A(\rvcpu.dp.plfd.PCPlus4D[20] ),
    .B(_11397_),
    .X(_11400_));
 sky130_fd_sc_hd__clkbuf_1 _26129_ (.A(_11400_),
    .X(_03017_));
 sky130_fd_sc_hd__and2_1 _26130_ (.A(\rvcpu.dp.plfd.PCPlus4D[21] ),
    .B(_11397_),
    .X(_11401_));
 sky130_fd_sc_hd__clkbuf_1 _26131_ (.A(_11401_),
    .X(_03018_));
 sky130_fd_sc_hd__and2_1 _26132_ (.A(\rvcpu.dp.plfd.PCPlus4D[22] ),
    .B(_11397_),
    .X(_11402_));
 sky130_fd_sc_hd__clkbuf_1 _26133_ (.A(_11402_),
    .X(_03019_));
 sky130_fd_sc_hd__and2_1 _26134_ (.A(\rvcpu.dp.plfd.PCPlus4D[23] ),
    .B(_11397_),
    .X(_11403_));
 sky130_fd_sc_hd__clkbuf_1 _26135_ (.A(_11403_),
    .X(_03020_));
 sky130_fd_sc_hd__and2_1 _26136_ (.A(\rvcpu.dp.plfd.PCPlus4D[24] ),
    .B(_11397_),
    .X(_11404_));
 sky130_fd_sc_hd__clkbuf_1 _26137_ (.A(_11404_),
    .X(_03021_));
 sky130_fd_sc_hd__and2_1 _26138_ (.A(\rvcpu.dp.plfd.PCPlus4D[25] ),
    .B(_11397_),
    .X(_11405_));
 sky130_fd_sc_hd__clkbuf_1 _26139_ (.A(_11405_),
    .X(_03022_));
 sky130_fd_sc_hd__and2_1 _26140_ (.A(\rvcpu.dp.plfd.PCPlus4D[26] ),
    .B(_11397_),
    .X(_11406_));
 sky130_fd_sc_hd__clkbuf_1 _26141_ (.A(_11406_),
    .X(_03023_));
 sky130_fd_sc_hd__and2_1 _26142_ (.A(\rvcpu.dp.plfd.PCPlus4D[27] ),
    .B(_11397_),
    .X(_11407_));
 sky130_fd_sc_hd__clkbuf_1 _26143_ (.A(_11407_),
    .X(_03024_));
 sky130_fd_sc_hd__clkbuf_2 _26144_ (.A(_11371_),
    .X(_11408_));
 sky130_fd_sc_hd__and2_1 _26145_ (.A(\rvcpu.dp.plfd.PCPlus4D[28] ),
    .B(_11408_),
    .X(_11409_));
 sky130_fd_sc_hd__clkbuf_1 _26146_ (.A(_11409_),
    .X(_03025_));
 sky130_fd_sc_hd__and2_1 _26147_ (.A(\rvcpu.dp.plfd.PCPlus4D[29] ),
    .B(_11408_),
    .X(_11410_));
 sky130_fd_sc_hd__clkbuf_1 _26148_ (.A(_11410_),
    .X(_03026_));
 sky130_fd_sc_hd__and2_1 _26149_ (.A(\rvcpu.dp.plfd.PCPlus4D[30] ),
    .B(_11408_),
    .X(_11411_));
 sky130_fd_sc_hd__clkbuf_1 _26150_ (.A(_11411_),
    .X(_03027_));
 sky130_fd_sc_hd__and2_1 _26151_ (.A(\rvcpu.dp.plfd.PCPlus4D[31] ),
    .B(_11408_),
    .X(_11412_));
 sky130_fd_sc_hd__clkbuf_1 _26152_ (.A(_11412_),
    .X(_03028_));
 sky130_fd_sc_hd__buf_2 _26153_ (.A(_08622_),
    .X(_11413_));
 sky130_fd_sc_hd__and2_1 _26154_ (.A(\rvcpu.dp.plfd.InstrD[13] ),
    .B(_11413_),
    .X(_11414_));
 sky130_fd_sc_hd__clkbuf_1 _26155_ (.A(_11414_),
    .X(_03030_));
 sky130_fd_sc_hd__and2_1 _26156_ (.A(\rvcpu.dp.plfd.InstrD[14] ),
    .B(_11413_),
    .X(_11415_));
 sky130_fd_sc_hd__clkbuf_1 _26157_ (.A(_11415_),
    .X(_03031_));
 sky130_fd_sc_hd__and2_1 _26158_ (.A(\rvcpu.dp.plfd.InstrD[7] ),
    .B(_11408_),
    .X(_11416_));
 sky130_fd_sc_hd__clkbuf_1 _26159_ (.A(_11416_),
    .X(_03032_));
 sky130_fd_sc_hd__and2_1 _26160_ (.A(\rvcpu.dp.plfd.InstrD[8] ),
    .B(_11408_),
    .X(_11417_));
 sky130_fd_sc_hd__clkbuf_1 _26161_ (.A(_11417_),
    .X(_03033_));
 sky130_fd_sc_hd__and2_1 _26162_ (.A(\rvcpu.dp.plfd.InstrD[9] ),
    .B(_11408_),
    .X(_11418_));
 sky130_fd_sc_hd__clkbuf_1 _26163_ (.A(_11418_),
    .X(_03034_));
 sky130_fd_sc_hd__and2_1 _26164_ (.A(\rvcpu.dp.plfd.InstrD[10] ),
    .B(_11408_),
    .X(_11419_));
 sky130_fd_sc_hd__clkbuf_1 _26165_ (.A(_11419_),
    .X(_03035_));
 sky130_fd_sc_hd__and2_1 _26166_ (.A(\rvcpu.dp.plfd.InstrD[11] ),
    .B(_11408_),
    .X(_11420_));
 sky130_fd_sc_hd__clkbuf_1 _26167_ (.A(_11420_),
    .X(_03036_));
 sky130_fd_sc_hd__and2_1 _26168_ (.A(_09478_),
    .B(_11362_),
    .X(_11421_));
 sky130_fd_sc_hd__clkbuf_1 _26169_ (.A(_11421_),
    .X(_03037_));
 sky130_fd_sc_hd__and2_1 _26170_ (.A(_09479_),
    .B(_11362_),
    .X(_11422_));
 sky130_fd_sc_hd__clkbuf_1 _26171_ (.A(_11422_),
    .X(_03038_));
 sky130_fd_sc_hd__and2_1 _26172_ (.A(_09482_),
    .B(_11362_),
    .X(_11423_));
 sky130_fd_sc_hd__clkbuf_1 _26173_ (.A(_11423_),
    .X(_03039_));
 sky130_fd_sc_hd__and2_1 _26174_ (.A(_09457_),
    .B(_11362_),
    .X(_11424_));
 sky130_fd_sc_hd__clkbuf_1 _26175_ (.A(_11424_),
    .X(_03040_));
 sky130_fd_sc_hd__and2_1 _26176_ (.A(\rvcpu.dp.plfd.InstrD[24] ),
    .B(_11362_),
    .X(_11425_));
 sky130_fd_sc_hd__clkbuf_1 _26177_ (.A(_11425_),
    .X(_03041_));
 sky130_fd_sc_hd__and2_1 _26178_ (.A(_08567_),
    .B(_11413_),
    .X(_11426_));
 sky130_fd_sc_hd__clkbuf_1 _26179_ (.A(_11426_),
    .X(_03042_));
 sky130_fd_sc_hd__and2_1 _26180_ (.A(_08570_),
    .B(_11413_),
    .X(_11427_));
 sky130_fd_sc_hd__clkbuf_1 _26181_ (.A(_11427_),
    .X(_03043_));
 sky130_fd_sc_hd__and2_1 _26182_ (.A(_08572_),
    .B(_11413_),
    .X(_11428_));
 sky130_fd_sc_hd__clkbuf_1 _26183_ (.A(_11428_),
    .X(_03044_));
 sky130_fd_sc_hd__and2_1 _26184_ (.A(_08513_),
    .B(_11413_),
    .X(_11429_));
 sky130_fd_sc_hd__clkbuf_1 _26185_ (.A(_11429_),
    .X(_03045_));
 sky130_fd_sc_hd__and2_1 _26186_ (.A(\rvcpu.dp.plfd.InstrD[19] ),
    .B(_11362_),
    .X(_11430_));
 sky130_fd_sc_hd__clkbuf_1 _26187_ (.A(_11430_),
    .X(_03046_));
 sky130_fd_sc_hd__and2_1 _26188_ (.A(\rvcpu.ALUControl[0] ),
    .B(_11408_),
    .X(_11431_));
 sky130_fd_sc_hd__clkbuf_1 _26189_ (.A(_11431_),
    .X(_03047_));
 sky130_fd_sc_hd__clkbuf_4 _26190_ (.A(_11413_),
    .X(_11432_));
 sky130_fd_sc_hd__and2_1 _26191_ (.A(\rvcpu.ALUControl[1] ),
    .B(_11432_),
    .X(_11433_));
 sky130_fd_sc_hd__clkbuf_1 _26192_ (.A(_11433_),
    .X(_03048_));
 sky130_fd_sc_hd__and2_1 _26193_ (.A(\rvcpu.ALUControl[2] ),
    .B(_11432_),
    .X(_11434_));
 sky130_fd_sc_hd__clkbuf_1 _26194_ (.A(_11434_),
    .X(_03049_));
 sky130_fd_sc_hd__and2_1 _26195_ (.A(\rvcpu.ALUControl[3] ),
    .B(_11432_),
    .X(_11435_));
 sky130_fd_sc_hd__clkbuf_1 _26196_ (.A(_11435_),
    .X(_03050_));
 sky130_fd_sc_hd__clkbuf_2 _26197_ (.A(_11413_),
    .X(_11436_));
 sky130_fd_sc_hd__and3_1 _26198_ (.A(\rvcpu.c.ad.opb5 ),
    .B(_11436_),
    .C(_11377_),
    .X(_11437_));
 sky130_fd_sc_hd__clkbuf_1 _26199_ (.A(_11437_),
    .X(_03051_));
 sky130_fd_sc_hd__clkbuf_2 _26200_ (.A(net116),
    .X(_11438_));
 sky130_fd_sc_hd__o21a_1 _26201_ (.A1(_11375_),
    .A2(_11438_),
    .B1(_11372_),
    .X(_03052_));
 sky130_fd_sc_hd__and2_1 _26202_ (.A(_11362_),
    .B(net116),
    .X(_11439_));
 sky130_fd_sc_hd__or3_1 _26203_ (.A(_02995_),
    .B(_02996_),
    .C(_11439_),
    .X(_11440_));
 sky130_fd_sc_hd__buf_1 _26204_ (.A(_11440_),
    .X(_03053_));
 sky130_fd_sc_hd__nor2_1 _26205_ (.A(_11361_),
    .B(_11379_),
    .Y(_11441_));
 sky130_fd_sc_hd__a22o_1 _26206_ (.A1(\rvcpu.dp.plfd.InstrD[7] ),
    .A2(_02993_),
    .B1(_03037_),
    .B2(_11441_),
    .X(_03054_));
 sky130_fd_sc_hd__and2_1 _26207_ (.A(_11361_),
    .B(_11371_),
    .X(_11442_));
 sky130_fd_sc_hd__or2_1 _26208_ (.A(_11369_),
    .B(_11441_),
    .X(_11443_));
 sky130_fd_sc_hd__a22o_1 _26209_ (.A1(\rvcpu.dp.plfd.InstrD[8] ),
    .A2(_11442_),
    .B1(_03038_),
    .B2(_11443_),
    .X(_03055_));
 sky130_fd_sc_hd__a22o_1 _26210_ (.A1(\rvcpu.dp.plfd.InstrD[9] ),
    .A2(_11442_),
    .B1(_03039_),
    .B2(_11443_),
    .X(_03056_));
 sky130_fd_sc_hd__a22o_1 _26211_ (.A1(\rvcpu.dp.plfd.InstrD[10] ),
    .A2(_11442_),
    .B1(_03040_),
    .B2(_11443_),
    .X(_03057_));
 sky130_fd_sc_hd__a22o_1 _26212_ (.A1(\rvcpu.dp.plfd.InstrD[11] ),
    .A2(_11442_),
    .B1(_03041_),
    .B2(_11443_),
    .X(_03058_));
 sky130_fd_sc_hd__or4b_2 _26213_ (.A(\rvcpu.dp.plfd.InstrD[6] ),
    .B(\rvcpu.dp.plfd.InstrD[3] ),
    .C(_11376_),
    .D_N(\rvcpu.dp.plfd.InstrD[4] ),
    .X(_11444_));
 sky130_fd_sc_hd__and3_1 _26214_ (.A(\rvcpu.dp.plfd.InstrD[25] ),
    .B(_11436_),
    .C(_11444_),
    .X(_11445_));
 sky130_fd_sc_hd__clkbuf_1 _26215_ (.A(_11445_),
    .X(_03059_));
 sky130_fd_sc_hd__and3_1 _26216_ (.A(\rvcpu.dp.plfd.InstrD[26] ),
    .B(_11436_),
    .C(_11444_),
    .X(_11446_));
 sky130_fd_sc_hd__clkbuf_1 _26217_ (.A(_11446_),
    .X(_03060_));
 sky130_fd_sc_hd__and3_1 _26218_ (.A(\rvcpu.dp.plfd.InstrD[27] ),
    .B(_11436_),
    .C(_11444_),
    .X(_11447_));
 sky130_fd_sc_hd__clkbuf_1 _26219_ (.A(_11447_),
    .X(_03061_));
 sky130_fd_sc_hd__and3_1 _26220_ (.A(\rvcpu.dp.plfd.InstrD[28] ),
    .B(_11436_),
    .C(_11444_),
    .X(_11448_));
 sky130_fd_sc_hd__clkbuf_1 _26221_ (.A(_11448_),
    .X(_03062_));
 sky130_fd_sc_hd__and3_1 _26222_ (.A(\rvcpu.dp.plfd.InstrD[29] ),
    .B(_11371_),
    .C(_11444_),
    .X(_11449_));
 sky130_fd_sc_hd__clkbuf_1 _26223_ (.A(_11449_),
    .X(_03063_));
 sky130_fd_sc_hd__and3_1 _26224_ (.A(\rvcpu.c.ad.funct7b5 ),
    .B(_11371_),
    .C(_11444_),
    .X(_11450_));
 sky130_fd_sc_hd__clkbuf_1 _26225_ (.A(_11450_),
    .X(_03064_));
 sky130_fd_sc_hd__nand2_1 _26226_ (.A(\rvcpu.dp.plfd.InstrD[6] ),
    .B(_11361_),
    .Y(_11451_));
 sky130_fd_sc_hd__inv_2 _26227_ (.A(_11378_),
    .Y(_11452_));
 sky130_fd_sc_hd__and3_1 _26228_ (.A(\rvcpu.dp.plfd.InstrD[31] ),
    .B(_11362_),
    .C(_11452_),
    .X(_11453_));
 sky130_fd_sc_hd__buf_2 _26229_ (.A(_11453_),
    .X(_11454_));
 sky130_fd_sc_hd__and3_1 _26230_ (.A(_09478_),
    .B(_11371_),
    .C(_11369_),
    .X(_11455_));
 sky130_fd_sc_hd__and3_1 _26231_ (.A(\rvcpu.dp.plfd.InstrD[7] ),
    .B(_06573_),
    .C(_11371_),
    .X(_11456_));
 sky130_fd_sc_hd__a211o_1 _26232_ (.A1(_11451_),
    .A2(_11454_),
    .B1(_11455_),
    .C1(_11456_),
    .X(_03065_));
 sky130_fd_sc_hd__a21o_1 _26233_ (.A1(_03029_),
    .A2(_11379_),
    .B1(_11454_),
    .X(_03066_));
 sky130_fd_sc_hd__a21o_1 _26234_ (.A1(_11379_),
    .A2(_03030_),
    .B1(_11454_),
    .X(_03067_));
 sky130_fd_sc_hd__a21o_1 _26235_ (.A1(_11379_),
    .A2(_03031_),
    .B1(_11454_),
    .X(_03068_));
 sky130_fd_sc_hd__a21o_1 _26236_ (.A1(_11379_),
    .A2(_03042_),
    .B1(_11454_),
    .X(_03069_));
 sky130_fd_sc_hd__a21o_1 _26237_ (.A1(_11379_),
    .A2(_03043_),
    .B1(_11454_),
    .X(_03070_));
 sky130_fd_sc_hd__a21o_1 _26238_ (.A1(_11379_),
    .A2(_03044_),
    .B1(_11454_),
    .X(_03071_));
 sky130_fd_sc_hd__a21o_1 _26239_ (.A1(_11379_),
    .A2(_03045_),
    .B1(_11454_),
    .X(_03072_));
 sky130_fd_sc_hd__a21o_1 _26240_ (.A1(_11379_),
    .A2(_03046_),
    .B1(_11454_),
    .X(_03073_));
 sky130_fd_sc_hd__nand2_1 _26241_ (.A(\rvcpu.dp.plfd.InstrD[31] ),
    .B(_11371_),
    .Y(_11457_));
 sky130_fd_sc_hd__clkbuf_2 _26242_ (.A(_11457_),
    .X(_11458_));
 sky130_fd_sc_hd__clkbuf_2 _26243_ (.A(_11439_),
    .X(_11459_));
 sky130_fd_sc_hd__a2bb2o_1 _26244_ (.A1_N(_11438_),
    .A2_N(_11458_),
    .B1(_11459_),
    .B2(_09478_),
    .X(_03074_));
 sky130_fd_sc_hd__a2bb2o_1 _26245_ (.A1_N(_11438_),
    .A2_N(_11458_),
    .B1(_11459_),
    .B2(_09479_),
    .X(_03075_));
 sky130_fd_sc_hd__a2bb2o_1 _26246_ (.A1_N(_11438_),
    .A2_N(_11458_),
    .B1(_11459_),
    .B2(_09482_),
    .X(_03076_));
 sky130_fd_sc_hd__a2bb2o_1 _26247_ (.A1_N(_11438_),
    .A2_N(_11458_),
    .B1(_11459_),
    .B2(_09457_),
    .X(_03077_));
 sky130_fd_sc_hd__a2bb2o_1 _26248_ (.A1_N(_11438_),
    .A2_N(_11458_),
    .B1(_11459_),
    .B2(\rvcpu.dp.plfd.InstrD[24] ),
    .X(_03078_));
 sky130_fd_sc_hd__a2bb2o_1 _26249_ (.A1_N(_11438_),
    .A2_N(_11458_),
    .B1(_11459_),
    .B2(\rvcpu.dp.plfd.InstrD[25] ),
    .X(_03079_));
 sky130_fd_sc_hd__a2bb2o_1 _26250_ (.A1_N(_11438_),
    .A2_N(_11458_),
    .B1(_11459_),
    .B2(\rvcpu.dp.plfd.InstrD[26] ),
    .X(_03080_));
 sky130_fd_sc_hd__a2bb2o_1 _26251_ (.A1_N(_11438_),
    .A2_N(_11458_),
    .B1(_11459_),
    .B2(\rvcpu.dp.plfd.InstrD[27] ),
    .X(_03081_));
 sky130_fd_sc_hd__a2bb2o_1 _26252_ (.A1_N(_11438_),
    .A2_N(_11458_),
    .B1(_11459_),
    .B2(\rvcpu.dp.plfd.InstrD[28] ),
    .X(_03082_));
 sky130_fd_sc_hd__a2bb2o_1 _26253_ (.A1_N(net116),
    .A2_N(_11457_),
    .B1(_11459_),
    .B2(\rvcpu.dp.plfd.InstrD[29] ),
    .X(_03083_));
 sky130_fd_sc_hd__a2bb2o_1 _26254_ (.A1_N(net116),
    .A2_N(_11457_),
    .B1(_11439_),
    .B2(\rvcpu.c.ad.funct7b5 ),
    .X(_03084_));
 sky130_fd_sc_hd__inv_2 _26255_ (.A(_11458_),
    .Y(_03085_));
 sky130_fd_sc_hd__and2_1 _26256_ (.A(\rvcpu.dp.plfd.PCD[0] ),
    .B(_11432_),
    .X(_11460_));
 sky130_fd_sc_hd__clkbuf_1 _26257_ (.A(_11460_),
    .X(_03086_));
 sky130_fd_sc_hd__and2_1 _26258_ (.A(\rvcpu.dp.plfd.PCD[1] ),
    .B(_11432_),
    .X(_11461_));
 sky130_fd_sc_hd__clkbuf_1 _26259_ (.A(_11461_),
    .X(_03087_));
 sky130_fd_sc_hd__and2_1 _26260_ (.A(\rvcpu.dp.plfd.PCD[2] ),
    .B(_11432_),
    .X(_11462_));
 sky130_fd_sc_hd__clkbuf_1 _26261_ (.A(_11462_),
    .X(_03088_));
 sky130_fd_sc_hd__and2_1 _26262_ (.A(\rvcpu.dp.plfd.PCD[3] ),
    .B(_11432_),
    .X(_11463_));
 sky130_fd_sc_hd__clkbuf_1 _26263_ (.A(_11463_),
    .X(_03089_));
 sky130_fd_sc_hd__and2_1 _26264_ (.A(\rvcpu.dp.plfd.PCD[4] ),
    .B(_11432_),
    .X(_11464_));
 sky130_fd_sc_hd__clkbuf_1 _26265_ (.A(_11464_),
    .X(_03090_));
 sky130_fd_sc_hd__and2_1 _26266_ (.A(\rvcpu.dp.plfd.PCD[5] ),
    .B(_11432_),
    .X(_11465_));
 sky130_fd_sc_hd__clkbuf_1 _26267_ (.A(_11465_),
    .X(_03091_));
 sky130_fd_sc_hd__and2_1 _26268_ (.A(\rvcpu.dp.plfd.PCD[6] ),
    .B(_11432_),
    .X(_11466_));
 sky130_fd_sc_hd__clkbuf_1 _26269_ (.A(_11466_),
    .X(_03092_));
 sky130_fd_sc_hd__buf_2 _26270_ (.A(_11413_),
    .X(_11467_));
 sky130_fd_sc_hd__and2_1 _26271_ (.A(\rvcpu.dp.plfd.PCD[7] ),
    .B(_11467_),
    .X(_11468_));
 sky130_fd_sc_hd__clkbuf_1 _26272_ (.A(_11468_),
    .X(_03093_));
 sky130_fd_sc_hd__and2_1 _26273_ (.A(\rvcpu.dp.plfd.PCD[8] ),
    .B(_11467_),
    .X(_11469_));
 sky130_fd_sc_hd__clkbuf_1 _26274_ (.A(_11469_),
    .X(_03094_));
 sky130_fd_sc_hd__and2_1 _26275_ (.A(\rvcpu.dp.plfd.PCD[9] ),
    .B(_11467_),
    .X(_11470_));
 sky130_fd_sc_hd__clkbuf_1 _26276_ (.A(_11470_),
    .X(_03095_));
 sky130_fd_sc_hd__and2_1 _26277_ (.A(\rvcpu.dp.plfd.PCD[10] ),
    .B(_11467_),
    .X(_11471_));
 sky130_fd_sc_hd__clkbuf_1 _26278_ (.A(_11471_),
    .X(_03096_));
 sky130_fd_sc_hd__and2_1 _26279_ (.A(\rvcpu.dp.plfd.PCD[11] ),
    .B(_11467_),
    .X(_11472_));
 sky130_fd_sc_hd__clkbuf_1 _26280_ (.A(_11472_),
    .X(_03097_));
 sky130_fd_sc_hd__and2_1 _26281_ (.A(\rvcpu.dp.plfd.PCD[12] ),
    .B(_11467_),
    .X(_11473_));
 sky130_fd_sc_hd__clkbuf_1 _26282_ (.A(_11473_),
    .X(_03098_));
 sky130_fd_sc_hd__and2_1 _26283_ (.A(\rvcpu.dp.plfd.PCD[13] ),
    .B(_11467_),
    .X(_11474_));
 sky130_fd_sc_hd__clkbuf_1 _26284_ (.A(_11474_),
    .X(_03099_));
 sky130_fd_sc_hd__and2_1 _26285_ (.A(\rvcpu.dp.plfd.PCD[14] ),
    .B(_11467_),
    .X(_11475_));
 sky130_fd_sc_hd__clkbuf_1 _26286_ (.A(_11475_),
    .X(_03100_));
 sky130_fd_sc_hd__and2_1 _26287_ (.A(\rvcpu.dp.plfd.PCD[15] ),
    .B(_11467_),
    .X(_11476_));
 sky130_fd_sc_hd__clkbuf_1 _26288_ (.A(_11476_),
    .X(_03101_));
 sky130_fd_sc_hd__and2_1 _26289_ (.A(\rvcpu.dp.plfd.PCD[16] ),
    .B(_11467_),
    .X(_11477_));
 sky130_fd_sc_hd__clkbuf_1 _26290_ (.A(_11477_),
    .X(_03102_));
 sky130_fd_sc_hd__buf_2 _26291_ (.A(_11413_),
    .X(_11478_));
 sky130_fd_sc_hd__and2_1 _26292_ (.A(\rvcpu.dp.plfd.PCD[17] ),
    .B(_11478_),
    .X(_11479_));
 sky130_fd_sc_hd__clkbuf_1 _26293_ (.A(_11479_),
    .X(_03103_));
 sky130_fd_sc_hd__and2_1 _26294_ (.A(\rvcpu.dp.plfd.PCD[18] ),
    .B(_11478_),
    .X(_11480_));
 sky130_fd_sc_hd__clkbuf_1 _26295_ (.A(_11480_),
    .X(_03104_));
 sky130_fd_sc_hd__and2_1 _26296_ (.A(\rvcpu.dp.plfd.PCD[19] ),
    .B(_11478_),
    .X(_11481_));
 sky130_fd_sc_hd__clkbuf_1 _26297_ (.A(_11481_),
    .X(_03105_));
 sky130_fd_sc_hd__and2_1 _26298_ (.A(\rvcpu.dp.plfd.PCD[20] ),
    .B(_11478_),
    .X(_11482_));
 sky130_fd_sc_hd__clkbuf_1 _26299_ (.A(_11482_),
    .X(_03106_));
 sky130_fd_sc_hd__and2_1 _26300_ (.A(\rvcpu.dp.plfd.PCD[21] ),
    .B(_11478_),
    .X(_11483_));
 sky130_fd_sc_hd__clkbuf_1 _26301_ (.A(_11483_),
    .X(_03107_));
 sky130_fd_sc_hd__and2_1 _26302_ (.A(\rvcpu.dp.plfd.PCD[22] ),
    .B(_11478_),
    .X(_11484_));
 sky130_fd_sc_hd__clkbuf_1 _26303_ (.A(_11484_),
    .X(_03108_));
 sky130_fd_sc_hd__and2_1 _26304_ (.A(\rvcpu.dp.plfd.PCD[23] ),
    .B(_11478_),
    .X(_11485_));
 sky130_fd_sc_hd__clkbuf_1 _26305_ (.A(_11485_),
    .X(_03109_));
 sky130_fd_sc_hd__and2_1 _26306_ (.A(\rvcpu.dp.plfd.PCD[24] ),
    .B(_11478_),
    .X(_11486_));
 sky130_fd_sc_hd__clkbuf_1 _26307_ (.A(_11486_),
    .X(_03110_));
 sky130_fd_sc_hd__and2_1 _26308_ (.A(\rvcpu.dp.plfd.PCD[25] ),
    .B(_11478_),
    .X(_11487_));
 sky130_fd_sc_hd__clkbuf_1 _26309_ (.A(_11487_),
    .X(_03111_));
 sky130_fd_sc_hd__and2_1 _26310_ (.A(\rvcpu.dp.plfd.PCD[26] ),
    .B(_11478_),
    .X(_11488_));
 sky130_fd_sc_hd__clkbuf_1 _26311_ (.A(_11488_),
    .X(_03112_));
 sky130_fd_sc_hd__and2_1 _26312_ (.A(\rvcpu.dp.plfd.PCD[27] ),
    .B(_11436_),
    .X(_11489_));
 sky130_fd_sc_hd__clkbuf_1 _26313_ (.A(_11489_),
    .X(_03113_));
 sky130_fd_sc_hd__and2_1 _26314_ (.A(\rvcpu.dp.plfd.PCD[28] ),
    .B(_11436_),
    .X(_11490_));
 sky130_fd_sc_hd__clkbuf_1 _26315_ (.A(_11490_),
    .X(_03114_));
 sky130_fd_sc_hd__and2_1 _26316_ (.A(\rvcpu.dp.plfd.PCD[29] ),
    .B(_11436_),
    .X(_11491_));
 sky130_fd_sc_hd__clkbuf_1 _26317_ (.A(_11491_),
    .X(_03115_));
 sky130_fd_sc_hd__and2_1 _26318_ (.A(\rvcpu.dp.plfd.PCD[30] ),
    .B(_11436_),
    .X(_11492_));
 sky130_fd_sc_hd__clkbuf_1 _26319_ (.A(_11492_),
    .X(_03116_));
 sky130_fd_sc_hd__and2_1 _26320_ (.A(\rvcpu.dp.plfd.PCD[31] ),
    .B(_11436_),
    .X(_11493_));
 sky130_fd_sc_hd__clkbuf_1 _26321_ (.A(_11493_),
    .X(_03117_));
 sky130_fd_sc_hd__buf_2 _26322_ (.A(_10043_),
    .X(_11494_));
 sky130_fd_sc_hd__or3_1 _26323_ (.A(_07791_),
    .B(_10932_),
    .C(_11494_),
    .X(_11495_));
 sky130_fd_sc_hd__clkbuf_2 _26324_ (.A(_11495_),
    .X(_11496_));
 sky130_fd_sc_hd__and3_2 _26325_ (.A(_10325_),
    .B(_10935_),
    .C(_10052_),
    .X(_11497_));
 sky130_fd_sc_hd__and2_1 _26326_ (.A(_11078_),
    .B(_11497_),
    .X(_11498_));
 sky130_fd_sc_hd__a31o_1 _26327_ (.A1(_11353_),
    .A2(\datamem.data_ram[15][0] ),
    .A3(_11496_),
    .B1(_11498_),
    .X(_03118_));
 sky130_fd_sc_hd__and2_1 _26328_ (.A(_11081_),
    .B(_11497_),
    .X(_11499_));
 sky130_fd_sc_hd__a31o_1 _26329_ (.A1(_11353_),
    .A2(\datamem.data_ram[15][1] ),
    .A3(_11496_),
    .B1(_11499_),
    .X(_03119_));
 sky130_fd_sc_hd__and2_1 _26330_ (.A(_11083_),
    .B(_11497_),
    .X(_11500_));
 sky130_fd_sc_hd__a31o_1 _26331_ (.A1(_11353_),
    .A2(\datamem.data_ram[15][2] ),
    .A3(_11496_),
    .B1(_11500_),
    .X(_03120_));
 sky130_fd_sc_hd__buf_2 _26332_ (.A(_11104_),
    .X(_11501_));
 sky130_fd_sc_hd__and2_1 _26333_ (.A(_11086_),
    .B(_11497_),
    .X(_11502_));
 sky130_fd_sc_hd__a31o_1 _26334_ (.A1(_11501_),
    .A2(\datamem.data_ram[15][3] ),
    .A3(_11496_),
    .B1(_11502_),
    .X(_03121_));
 sky130_fd_sc_hd__and2_1 _26335_ (.A(_11047_),
    .B(_11497_),
    .X(_11503_));
 sky130_fd_sc_hd__a31o_1 _26336_ (.A1(_11501_),
    .A2(\datamem.data_ram[15][4] ),
    .A3(_11496_),
    .B1(_11503_),
    .X(_03122_));
 sky130_fd_sc_hd__and2_1 _26337_ (.A(_11089_),
    .B(_11497_),
    .X(_11504_));
 sky130_fd_sc_hd__a31o_1 _26338_ (.A1(_11501_),
    .A2(\datamem.data_ram[15][5] ),
    .A3(_11496_),
    .B1(_11504_),
    .X(_03123_));
 sky130_fd_sc_hd__and2_1 _26339_ (.A(_11091_),
    .B(_11497_),
    .X(_11505_));
 sky130_fd_sc_hd__a31o_1 _26340_ (.A1(_11501_),
    .A2(\datamem.data_ram[15][6] ),
    .A3(_11496_),
    .B1(_11505_),
    .X(_03124_));
 sky130_fd_sc_hd__and2_1 _26341_ (.A(_11064_),
    .B(_11497_),
    .X(_11506_));
 sky130_fd_sc_hd__a31o_1 _26342_ (.A1(_11501_),
    .A2(\datamem.data_ram[15][7] ),
    .A3(_11496_),
    .B1(_11506_),
    .X(_03125_));
 sky130_fd_sc_hd__nor2_4 _26343_ (.A(_11039_),
    .B(_10600_),
    .Y(_11507_));
 sky130_fd_sc_hd__nor2_2 _26344_ (.A(_10780_),
    .B(_11507_),
    .Y(_11508_));
 sky130_fd_sc_hd__a22o_1 _26345_ (.A1(_10048_),
    .A2(_11507_),
    .B1(_11508_),
    .B2(\datamem.data_ram[44][0] ),
    .X(_03126_));
 sky130_fd_sc_hd__a22o_1 _26346_ (.A1(_10058_),
    .A2(_11507_),
    .B1(_11508_),
    .B2(\datamem.data_ram[44][1] ),
    .X(_03127_));
 sky130_fd_sc_hd__a22o_1 _26347_ (.A1(_10061_),
    .A2(_11507_),
    .B1(_11508_),
    .B2(\datamem.data_ram[44][2] ),
    .X(_03128_));
 sky130_fd_sc_hd__a22o_1 _26348_ (.A1(_10064_),
    .A2(_11507_),
    .B1(_11508_),
    .B2(\datamem.data_ram[44][3] ),
    .X(_03129_));
 sky130_fd_sc_hd__a22o_1 _26349_ (.A1(_10782_),
    .A2(_11507_),
    .B1(_11508_),
    .B2(\datamem.data_ram[44][4] ),
    .X(_03130_));
 sky130_fd_sc_hd__a22o_1 _26350_ (.A1(_10070_),
    .A2(_11507_),
    .B1(_11508_),
    .B2(\datamem.data_ram[44][5] ),
    .X(_03131_));
 sky130_fd_sc_hd__a22o_1 _26351_ (.A1(_10073_),
    .A2(_11507_),
    .B1(_11508_),
    .B2(\datamem.data_ram[44][6] ),
    .X(_03132_));
 sky130_fd_sc_hd__a22o_1 _26352_ (.A1(_10783_),
    .A2(_11507_),
    .B1(_11508_),
    .B2(\datamem.data_ram[44][7] ),
    .X(_03133_));
 sky130_fd_sc_hd__or3_1 _26353_ (.A(_07028_),
    .B(_10932_),
    .C(_11494_),
    .X(_11509_));
 sky130_fd_sc_hd__clkbuf_2 _26354_ (.A(_11509_),
    .X(_11510_));
 sky130_fd_sc_hd__and3_2 _26355_ (.A(_09226_),
    .B(_10935_),
    .C(_10052_),
    .X(_11511_));
 sky130_fd_sc_hd__and2_1 _26356_ (.A(_11078_),
    .B(_11511_),
    .X(_11512_));
 sky130_fd_sc_hd__a31o_1 _26357_ (.A1(_11501_),
    .A2(\datamem.data_ram[14][0] ),
    .A3(_11510_),
    .B1(_11512_),
    .X(_03134_));
 sky130_fd_sc_hd__and2_1 _26358_ (.A(_11081_),
    .B(_11511_),
    .X(_11513_));
 sky130_fd_sc_hd__a31o_1 _26359_ (.A1(_11501_),
    .A2(\datamem.data_ram[14][1] ),
    .A3(_11510_),
    .B1(_11513_),
    .X(_03135_));
 sky130_fd_sc_hd__and2_1 _26360_ (.A(_11083_),
    .B(_11511_),
    .X(_11514_));
 sky130_fd_sc_hd__a31o_1 _26361_ (.A1(_11501_),
    .A2(\datamem.data_ram[14][2] ),
    .A3(_11510_),
    .B1(_11514_),
    .X(_03136_));
 sky130_fd_sc_hd__and2_1 _26362_ (.A(_11086_),
    .B(_11511_),
    .X(_11515_));
 sky130_fd_sc_hd__a31o_1 _26363_ (.A1(_11501_),
    .A2(\datamem.data_ram[14][3] ),
    .A3(_11510_),
    .B1(_11515_),
    .X(_03137_));
 sky130_fd_sc_hd__and2_1 _26364_ (.A(_11047_),
    .B(_11511_),
    .X(_11516_));
 sky130_fd_sc_hd__a31o_1 _26365_ (.A1(_11501_),
    .A2(\datamem.data_ram[14][4] ),
    .A3(_11510_),
    .B1(_11516_),
    .X(_03138_));
 sky130_fd_sc_hd__buf_2 _26366_ (.A(_11104_),
    .X(_11517_));
 sky130_fd_sc_hd__and2_1 _26367_ (.A(_11089_),
    .B(_11511_),
    .X(_11518_));
 sky130_fd_sc_hd__a31o_1 _26368_ (.A1(_11517_),
    .A2(\datamem.data_ram[14][5] ),
    .A3(_11510_),
    .B1(_11518_),
    .X(_03139_));
 sky130_fd_sc_hd__and2_1 _26369_ (.A(_11091_),
    .B(_11511_),
    .X(_11519_));
 sky130_fd_sc_hd__a31o_1 _26370_ (.A1(_11517_),
    .A2(\datamem.data_ram[14][6] ),
    .A3(_11510_),
    .B1(_11519_),
    .X(_03140_));
 sky130_fd_sc_hd__and2_1 _26371_ (.A(_11064_),
    .B(_11511_),
    .X(_11520_));
 sky130_fd_sc_hd__a31o_1 _26372_ (.A1(_11517_),
    .A2(\datamem.data_ram[14][7] ),
    .A3(_11510_),
    .B1(_11520_),
    .X(_03141_));
 sky130_fd_sc_hd__a21oi_1 _26373_ (.A1(_08620_),
    .A2(_08621_),
    .B1(\rvcpu.dp.plde.JalrE ),
    .Y(_11521_));
 sky130_fd_sc_hd__buf_2 _26374_ (.A(_11521_),
    .X(_11522_));
 sky130_fd_sc_hd__and2_1 _26375_ (.A(_06365_),
    .B(_11522_),
    .X(_11523_));
 sky130_fd_sc_hd__clkbuf_4 _26376_ (.A(\rvcpu.dp.plde.JalrE ),
    .X(_11524_));
 sky130_fd_sc_hd__a21o_1 _26377_ (.A1(_08620_),
    .A2(_08621_),
    .B1(_11151_),
    .X(_11525_));
 sky130_fd_sc_hd__buf_2 _26378_ (.A(_11525_),
    .X(_11526_));
 sky130_fd_sc_hd__a22o_1 _26379_ (.A1(_11524_),
    .A2(\rvcpu.ALUResultE[2] ),
    .B1(_11148_),
    .B2(_11526_),
    .X(_11527_));
 sky130_fd_sc_hd__o221a_1 _26380_ (.A1(_13328_),
    .A2(_11268_),
    .B1(_11523_),
    .B2(_11527_),
    .C1(_10041_),
    .X(_03142_));
 sky130_fd_sc_hd__a22o_1 _26381_ (.A1(_11524_),
    .A2(\rvcpu.ALUResultE[3] ),
    .B1(_06371_),
    .B2(_11522_),
    .X(_11528_));
 sky130_fd_sc_hd__clkbuf_4 _26382_ (.A(_11525_),
    .X(_11529_));
 sky130_fd_sc_hd__and2_1 _26383_ (.A(_11150_),
    .B(_11529_),
    .X(_11530_));
 sky130_fd_sc_hd__o221a_1 _26384_ (.A1(_13665_),
    .A2(_11268_),
    .B1(_11528_),
    .B2(_11530_),
    .C1(_10041_),
    .X(_03143_));
 sky130_fd_sc_hd__a31o_1 _26385_ (.A1(_08620_),
    .A2(_08621_),
    .A3(_11154_),
    .B1(_11157_),
    .X(_11531_));
 sky130_fd_sc_hd__a221o_1 _26386_ (.A1(_11524_),
    .A2(\rvcpu.ALUResultE[4] ),
    .B1(_06377_),
    .B2(_11522_),
    .C1(_11531_),
    .X(_11532_));
 sky130_fd_sc_hd__clkbuf_4 _26387_ (.A(_06587_),
    .X(_11533_));
 sky130_fd_sc_hd__clkbuf_4 _26388_ (.A(_11533_),
    .X(_11534_));
 sky130_fd_sc_hd__o211a_1 _26389_ (.A1(_13387_),
    .A2(_11329_),
    .B1(_11532_),
    .C1(_11534_),
    .X(_03144_));
 sky130_fd_sc_hd__buf_2 _26390_ (.A(\rvcpu.dp.plde.JalrE ),
    .X(_11535_));
 sky130_fd_sc_hd__and2_1 _26391_ (.A(_11535_),
    .B(\rvcpu.ALUResultE[5] ),
    .X(_11536_));
 sky130_fd_sc_hd__a221o_1 _26392_ (.A1(_06384_),
    .A2(_11522_),
    .B1(_11526_),
    .B2(_11158_),
    .C1(_11536_),
    .X(_11537_));
 sky130_fd_sc_hd__o211a_1 _26393_ (.A1(_13682_),
    .A2(_11329_),
    .B1(_11537_),
    .C1(_11534_),
    .X(_03145_));
 sky130_fd_sc_hd__nand2_1 _26394_ (.A(_11161_),
    .B(_11526_),
    .Y(_11538_));
 sky130_fd_sc_hd__clkbuf_4 _26395_ (.A(_11521_),
    .X(_11539_));
 sky130_fd_sc_hd__clkbuf_4 _26396_ (.A(_11539_),
    .X(_11540_));
 sky130_fd_sc_hd__a22oi_1 _26397_ (.A1(_11524_),
    .A2(\rvcpu.ALUResultE[6] ),
    .B1(_06392_),
    .B2(_11540_),
    .Y(_11541_));
 sky130_fd_sc_hd__a221oi_1 _26398_ (.A1(_13517_),
    .A2(_11153_),
    .B1(_11538_),
    .B2(_11541_),
    .C1(_10780_),
    .Y(_03146_));
 sky130_fd_sc_hd__clkbuf_4 _26399_ (.A(_11143_),
    .X(_11542_));
 sky130_fd_sc_hd__and2_1 _26400_ (.A(_11535_),
    .B(\rvcpu.ALUResultE[7] ),
    .X(_11543_));
 sky130_fd_sc_hd__a221o_1 _26401_ (.A1(_06398_),
    .A2(_11522_),
    .B1(_11526_),
    .B2(_11164_),
    .C1(_11543_),
    .X(_11544_));
 sky130_fd_sc_hd__o211a_1 _26402_ (.A1(_13706_),
    .A2(_11542_),
    .B1(_11544_),
    .C1(_11534_),
    .X(_03147_));
 sky130_fd_sc_hd__clkbuf_2 _26403_ (.A(\rvcpu.dp.plde.JalrE ),
    .X(_11545_));
 sky130_fd_sc_hd__and2_1 _26404_ (.A(_11545_),
    .B(\rvcpu.ALUResultE[8] ),
    .X(_11546_));
 sky130_fd_sc_hd__a221o_1 _26405_ (.A1(_06404_),
    .A2(_11522_),
    .B1(_11526_),
    .B2(_11167_),
    .C1(_11546_),
    .X(_11547_));
 sky130_fd_sc_hd__o211a_1 _26406_ (.A1(_13439_),
    .A2(_11542_),
    .B1(_11547_),
    .C1(_11534_),
    .X(_03148_));
 sky130_fd_sc_hd__nand2_1 _26407_ (.A(_06411_),
    .B(_11540_),
    .Y(_11548_));
 sky130_fd_sc_hd__nand2_1 _26408_ (.A(_11524_),
    .B(\rvcpu.ALUResultE[9] ),
    .Y(_11549_));
 sky130_fd_sc_hd__nand2_1 _26409_ (.A(_11170_),
    .B(_11526_),
    .Y(_11550_));
 sky130_fd_sc_hd__a21o_1 _26410_ (.A1(_13539_),
    .A2(_11152_),
    .B1(_10780_),
    .X(_11551_));
 sky130_fd_sc_hd__a31oi_1 _26411_ (.A1(_11548_),
    .A2(_11549_),
    .A3(_11550_),
    .B1(_11551_),
    .Y(_03149_));
 sky130_fd_sc_hd__and2_1 _26412_ (.A(_06418_),
    .B(_11522_),
    .X(_11552_));
 sky130_fd_sc_hd__a22o_1 _26413_ (.A1(_11524_),
    .A2(\rvcpu.ALUResultE[10] ),
    .B1(_11173_),
    .B2(_11526_),
    .X(_11553_));
 sky130_fd_sc_hd__o221a_1 _26414_ (.A1(\rvcpu.dp.pcreg.q[10] ),
    .A2(_11268_),
    .B1(_11552_),
    .B2(_11553_),
    .C1(_10041_),
    .X(_03150_));
 sky130_fd_sc_hd__and2_1 _26415_ (.A(_11545_),
    .B(\rvcpu.ALUResultE[11] ),
    .X(_11554_));
 sky130_fd_sc_hd__a221o_1 _26416_ (.A1(_06425_),
    .A2(_11539_),
    .B1(_11529_),
    .B2(_11176_),
    .C1(_11554_),
    .X(_11555_));
 sky130_fd_sc_hd__o211a_1 _26417_ (.A1(\rvcpu.dp.pcreg.q[11] ),
    .A2(_11542_),
    .B1(_11555_),
    .C1(_11534_),
    .X(_03151_));
 sky130_fd_sc_hd__and2_1 _26418_ (.A(_11545_),
    .B(\rvcpu.ALUResultE[12] ),
    .X(_11556_));
 sky130_fd_sc_hd__a221o_1 _26419_ (.A1(_06432_),
    .A2(_11539_),
    .B1(_11529_),
    .B2(_11180_),
    .C1(_11556_),
    .X(_11557_));
 sky130_fd_sc_hd__o211a_1 _26420_ (.A1(\rvcpu.dp.pcreg.q[12] ),
    .A2(_11542_),
    .B1(_11557_),
    .C1(_11534_),
    .X(_03152_));
 sky130_fd_sc_hd__and2_1 _26421_ (.A(_11545_),
    .B(\rvcpu.ALUResultE[13] ),
    .X(_11558_));
 sky130_fd_sc_hd__a221o_1 _26422_ (.A1(_06438_),
    .A2(_11539_),
    .B1(_11529_),
    .B2(_11184_),
    .C1(_11558_),
    .X(_11559_));
 sky130_fd_sc_hd__o211a_1 _26423_ (.A1(\rvcpu.dp.pcreg.q[13] ),
    .A2(_11542_),
    .B1(_11559_),
    .C1(_11534_),
    .X(_03153_));
 sky130_fd_sc_hd__and2_1 _26424_ (.A(_11545_),
    .B(\rvcpu.ALUResultE[14] ),
    .X(_11560_));
 sky130_fd_sc_hd__a221o_1 _26425_ (.A1(_06447_),
    .A2(_11539_),
    .B1(_11529_),
    .B2(_11187_),
    .C1(_11560_),
    .X(_11561_));
 sky130_fd_sc_hd__o211a_1 _26426_ (.A1(\rvcpu.dp.pcreg.q[14] ),
    .A2(_11542_),
    .B1(_11561_),
    .C1(_11534_),
    .X(_03154_));
 sky130_fd_sc_hd__and2_1 _26427_ (.A(_11545_),
    .B(\rvcpu.ALUResultE[15] ),
    .X(_11562_));
 sky130_fd_sc_hd__a221o_1 _26428_ (.A1(_06453_),
    .A2(_11539_),
    .B1(_11529_),
    .B2(_11190_),
    .C1(_11562_),
    .X(_11563_));
 sky130_fd_sc_hd__o211a_1 _26429_ (.A1(\rvcpu.dp.pcreg.q[15] ),
    .A2(_11542_),
    .B1(_11563_),
    .C1(_11534_),
    .X(_03155_));
 sky130_fd_sc_hd__and2_1 _26430_ (.A(_06461_),
    .B(_11522_),
    .X(_11564_));
 sky130_fd_sc_hd__a22o_1 _26431_ (.A1(_11524_),
    .A2(\rvcpu.ALUResultE[16] ),
    .B1(_11193_),
    .B2(_11526_),
    .X(_11565_));
 sky130_fd_sc_hd__o221a_1 _26432_ (.A1(\rvcpu.dp.pcreg.q[16] ),
    .A2(_11268_),
    .B1(_11564_),
    .B2(_11565_),
    .C1(_10041_),
    .X(_03156_));
 sky130_fd_sc_hd__and2_1 _26433_ (.A(_11545_),
    .B(\rvcpu.ALUResultE[17] ),
    .X(_11566_));
 sky130_fd_sc_hd__a221o_1 _26434_ (.A1(_06468_),
    .A2(_11539_),
    .B1(_11529_),
    .B2(_11196_),
    .C1(_11566_),
    .X(_11567_));
 sky130_fd_sc_hd__o211a_1 _26435_ (.A1(\rvcpu.dp.pcreg.q[17] ),
    .A2(_11542_),
    .B1(_11567_),
    .C1(_11534_),
    .X(_03157_));
 sky130_fd_sc_hd__and2_1 _26436_ (.A(_11545_),
    .B(\rvcpu.ALUResultE[18] ),
    .X(_11568_));
 sky130_fd_sc_hd__a221o_1 _26437_ (.A1(_06478_),
    .A2(_11539_),
    .B1(_11529_),
    .B2(_11199_),
    .C1(_11568_),
    .X(_11569_));
 sky130_fd_sc_hd__buf_2 _26438_ (.A(_11533_),
    .X(_11570_));
 sky130_fd_sc_hd__o211a_1 _26439_ (.A1(\rvcpu.dp.pcreg.q[18] ),
    .A2(_11542_),
    .B1(_11569_),
    .C1(_11570_),
    .X(_03158_));
 sky130_fd_sc_hd__and2_1 _26440_ (.A(_11545_),
    .B(\rvcpu.ALUResultE[19] ),
    .X(_11571_));
 sky130_fd_sc_hd__a221o_1 _26441_ (.A1(_06484_),
    .A2(_11539_),
    .B1(_11529_),
    .B2(_11202_),
    .C1(_11571_),
    .X(_11572_));
 sky130_fd_sc_hd__o211a_1 _26442_ (.A1(\rvcpu.dp.pcreg.q[19] ),
    .A2(_11542_),
    .B1(_11572_),
    .C1(_11570_),
    .X(_03159_));
 sky130_fd_sc_hd__clkbuf_4 _26443_ (.A(_11143_),
    .X(_11573_));
 sky130_fd_sc_hd__and2_1 _26444_ (.A(_11545_),
    .B(\rvcpu.ALUResultE[20] ),
    .X(_11574_));
 sky130_fd_sc_hd__a221o_1 _26445_ (.A1(_06492_),
    .A2(_11539_),
    .B1(_11529_),
    .B2(_11205_),
    .C1(_11574_),
    .X(_11575_));
 sky130_fd_sc_hd__o211a_1 _26446_ (.A1(\rvcpu.dp.pcreg.q[20] ),
    .A2(_11573_),
    .B1(_11575_),
    .C1(_11570_),
    .X(_03160_));
 sky130_fd_sc_hd__buf_2 _26447_ (.A(_11145_),
    .X(_11576_));
 sky130_fd_sc_hd__a21o_1 _26448_ (.A1(_11524_),
    .A2(\rvcpu.ALUResultE[21] ),
    .B1(_11288_),
    .X(_11577_));
 sky130_fd_sc_hd__a221o_1 _26449_ (.A1(_11576_),
    .A2(_11210_),
    .B1(_11540_),
    .B2(_06499_),
    .C1(_11577_),
    .X(_11578_));
 sky130_fd_sc_hd__o211a_1 _26450_ (.A1(\rvcpu.dp.pcreg.q[21] ),
    .A2(_11573_),
    .B1(_11578_),
    .C1(_11570_),
    .X(_03161_));
 sky130_fd_sc_hd__a21o_1 _26451_ (.A1(_11524_),
    .A2(\rvcpu.ALUResultE[22] ),
    .B1(_11288_),
    .X(_11579_));
 sky130_fd_sc_hd__a221o_1 _26452_ (.A1(_11576_),
    .A2(_11215_),
    .B1(_11540_),
    .B2(_06505_),
    .C1(_11579_),
    .X(_11580_));
 sky130_fd_sc_hd__o211a_1 _26453_ (.A1(\rvcpu.dp.pcreg.q[22] ),
    .A2(_11573_),
    .B1(_11580_),
    .C1(_11570_),
    .X(_03162_));
 sky130_fd_sc_hd__a21o_1 _26454_ (.A1(_11535_),
    .A2(\rvcpu.ALUResultE[23] ),
    .B1(_11288_),
    .X(_11581_));
 sky130_fd_sc_hd__a221o_1 _26455_ (.A1(_11576_),
    .A2(_11218_),
    .B1(_11540_),
    .B2(_06512_),
    .C1(_11581_),
    .X(_11582_));
 sky130_fd_sc_hd__o211a_1 _26456_ (.A1(\rvcpu.dp.pcreg.q[23] ),
    .A2(_11573_),
    .B1(_11582_),
    .C1(_11570_),
    .X(_03163_));
 sky130_fd_sc_hd__a21o_1 _26457_ (.A1(_11535_),
    .A2(\rvcpu.ALUResultE[24] ),
    .B1(_11288_),
    .X(_11583_));
 sky130_fd_sc_hd__a221o_1 _26458_ (.A1(_11576_),
    .A2(_11223_),
    .B1(_11540_),
    .B2(_06518_),
    .C1(_11583_),
    .X(_11584_));
 sky130_fd_sc_hd__o211a_1 _26459_ (.A1(\rvcpu.dp.pcreg.q[24] ),
    .A2(_11573_),
    .B1(_11584_),
    .C1(_11570_),
    .X(_03164_));
 sky130_fd_sc_hd__a21o_1 _26460_ (.A1(_11535_),
    .A2(\rvcpu.ALUResultE[25] ),
    .B1(_11288_),
    .X(_11585_));
 sky130_fd_sc_hd__a221o_1 _26461_ (.A1(_11576_),
    .A2(_11228_),
    .B1(_11540_),
    .B2(_06525_),
    .C1(_11585_),
    .X(_11586_));
 sky130_fd_sc_hd__o211a_1 _26462_ (.A1(\rvcpu.dp.pcreg.q[25] ),
    .A2(_11573_),
    .B1(_11586_),
    .C1(_11570_),
    .X(_03165_));
 sky130_fd_sc_hd__a21o_1 _26463_ (.A1(_11535_),
    .A2(\rvcpu.ALUResultE[26] ),
    .B1(_11288_),
    .X(_11587_));
 sky130_fd_sc_hd__a221o_1 _26464_ (.A1(_11576_),
    .A2(_11231_),
    .B1(_11540_),
    .B2(_06531_),
    .C1(_11587_),
    .X(_11588_));
 sky130_fd_sc_hd__o211a_1 _26465_ (.A1(\rvcpu.dp.pcreg.q[26] ),
    .A2(_11573_),
    .B1(_11588_),
    .C1(_11570_),
    .X(_03166_));
 sky130_fd_sc_hd__a21o_1 _26466_ (.A1(_11535_),
    .A2(\rvcpu.ALUResultE[27] ),
    .B1(_11288_),
    .X(_11589_));
 sky130_fd_sc_hd__a221o_1 _26467_ (.A1(_11576_),
    .A2(_11236_),
    .B1(_11540_),
    .B2(_06538_),
    .C1(_11589_),
    .X(_11590_));
 sky130_fd_sc_hd__o211a_1 _26468_ (.A1(\rvcpu.dp.pcreg.q[27] ),
    .A2(_11573_),
    .B1(_11590_),
    .C1(_11570_),
    .X(_03167_));
 sky130_fd_sc_hd__a21o_1 _26469_ (.A1(_11535_),
    .A2(\rvcpu.ALUResultE[28] ),
    .B1(_11288_),
    .X(_11591_));
 sky130_fd_sc_hd__a221o_1 _26470_ (.A1(_11576_),
    .A2(_11241_),
    .B1(_11540_),
    .B2(_06545_),
    .C1(_11591_),
    .X(_11592_));
 sky130_fd_sc_hd__o211a_1 _26471_ (.A1(\rvcpu.dp.pcreg.q[28] ),
    .A2(_11573_),
    .B1(_11592_),
    .C1(_10041_),
    .X(_03168_));
 sky130_fd_sc_hd__a21o_1 _26472_ (.A1(_11535_),
    .A2(\rvcpu.ALUResultE[29] ),
    .B1(_11288_),
    .X(_11593_));
 sky130_fd_sc_hd__a221o_1 _26473_ (.A1(_11576_),
    .A2(_11244_),
    .B1(_11522_),
    .B2(_06551_),
    .C1(_11593_),
    .X(_11594_));
 sky130_fd_sc_hd__o211a_1 _26474_ (.A1(\rvcpu.dp.pcreg.q[29] ),
    .A2(_11573_),
    .B1(_11594_),
    .C1(_10041_),
    .X(_03169_));
 sky130_fd_sc_hd__a21o_1 _26475_ (.A1(_11535_),
    .A2(\rvcpu.ALUResultE[30] ),
    .B1(_11157_),
    .X(_11595_));
 sky130_fd_sc_hd__a221o_1 _26476_ (.A1(_11576_),
    .A2(_11249_),
    .B1(_11522_),
    .B2(_06558_),
    .C1(_11595_),
    .X(_11596_));
 sky130_fd_sc_hd__o211a_1 _26477_ (.A1(\rvcpu.dp.pcreg.q[30] ),
    .A2(_11268_),
    .B1(_11596_),
    .C1(_10041_),
    .X(_03170_));
 sky130_fd_sc_hd__a21o_1 _26478_ (.A1(_08620_),
    .A2(_08621_),
    .B1(_06562_),
    .X(_11597_));
 sky130_fd_sc_hd__inv_2 _26479_ (.A(\rvcpu.dp.plde.JalrE ),
    .Y(_11598_));
 sky130_fd_sc_hd__o211ai_1 _26480_ (.A1(_11261_),
    .A2(_11253_),
    .B1(_11597_),
    .C1(_11598_),
    .Y(_11599_));
 sky130_fd_sc_hd__a21oi_1 _26481_ (.A1(_11524_),
    .A2(\rvcpu.ALUResultE[31] ),
    .B1(_11289_),
    .Y(_11600_));
 sky130_fd_sc_hd__a221oi_1 _26482_ (.A1(_11252_),
    .A2(_11153_),
    .B1(_11599_),
    .B2(_11600_),
    .C1(_10780_),
    .Y(_03171_));
 sky130_fd_sc_hd__inv_2 _26483_ (.A(_10267_),
    .Y(_00996_));
 sky130_fd_sc_hd__inv_2 _26484_ (.A(_10267_),
    .Y(_00997_));
 sky130_fd_sc_hd__inv_2 _26485_ (.A(_10267_),
    .Y(_00998_));
 sky130_fd_sc_hd__inv_2 _26486_ (.A(_10267_),
    .Y(_00999_));
 sky130_fd_sc_hd__inv_2 _26487_ (.A(_10267_),
    .Y(_01000_));
 sky130_fd_sc_hd__inv_2 _26488_ (.A(_10267_),
    .Y(_01001_));
 sky130_fd_sc_hd__inv_2 _26489_ (.A(_10267_),
    .Y(_01002_));
 sky130_fd_sc_hd__inv_2 _26490_ (.A(_10267_),
    .Y(_01003_));
 sky130_fd_sc_hd__buf_1 _26491_ (.A(_10079_),
    .X(_11601_));
 sky130_fd_sc_hd__inv_2 _26492_ (.A(_11601_),
    .Y(_01004_));
 sky130_fd_sc_hd__inv_2 _26493_ (.A(_11601_),
    .Y(_01005_));
 sky130_fd_sc_hd__inv_2 _26494_ (.A(_11601_),
    .Y(_01006_));
 sky130_fd_sc_hd__inv_2 _26495_ (.A(_11601_),
    .Y(_01007_));
 sky130_fd_sc_hd__inv_2 _26496_ (.A(_11601_),
    .Y(_01008_));
 sky130_fd_sc_hd__inv_2 _26497_ (.A(_11601_),
    .Y(_01009_));
 sky130_fd_sc_hd__inv_2 _26498_ (.A(_11601_),
    .Y(_01010_));
 sky130_fd_sc_hd__inv_2 _26499_ (.A(_11601_),
    .Y(_01011_));
 sky130_fd_sc_hd__inv_2 _26500_ (.A(_11601_),
    .Y(_01012_));
 sky130_fd_sc_hd__inv_2 _26501_ (.A(_11601_),
    .Y(_01013_));
 sky130_fd_sc_hd__buf_1 _26502_ (.A(_10079_),
    .X(_11602_));
 sky130_fd_sc_hd__inv_2 _26503_ (.A(_11602_),
    .Y(_01014_));
 sky130_fd_sc_hd__inv_2 _26504_ (.A(_11602_),
    .Y(_01015_));
 sky130_fd_sc_hd__inv_2 _26505_ (.A(_11602_),
    .Y(_01016_));
 sky130_fd_sc_hd__inv_2 _26506_ (.A(_11602_),
    .Y(_01017_));
 sky130_fd_sc_hd__inv_2 _26507_ (.A(_11602_),
    .Y(_01018_));
 sky130_fd_sc_hd__inv_2 _26508_ (.A(_11602_),
    .Y(_01019_));
 sky130_fd_sc_hd__inv_2 _26509_ (.A(_11602_),
    .Y(_01020_));
 sky130_fd_sc_hd__inv_2 _26510_ (.A(_11602_),
    .Y(_01021_));
 sky130_fd_sc_hd__inv_2 _26511_ (.A(_11602_),
    .Y(_01022_));
 sky130_fd_sc_hd__inv_2 _26512_ (.A(_11602_),
    .Y(_01023_));
 sky130_fd_sc_hd__inv_2 _26513_ (.A(_10080_),
    .Y(_01024_));
 sky130_fd_sc_hd__inv_2 _26514_ (.A(_10080_),
    .Y(_01025_));
 sky130_fd_sc_hd__inv_2 _26515_ (.A(_10080_),
    .Y(_01026_));
 sky130_fd_sc_hd__inv_2 _26516_ (.A(_10080_),
    .Y(_01027_));
 sky130_fd_sc_hd__nand2_4 _26517_ (.A(_07132_),
    .B(_10050_),
    .Y(_11603_));
 sky130_fd_sc_hd__nor2_4 _26518_ (.A(_11603_),
    .B(_10600_),
    .Y(_11604_));
 sky130_fd_sc_hd__nor2_2 _26519_ (.A(_10780_),
    .B(_11604_),
    .Y(_11605_));
 sky130_fd_sc_hd__a22o_1 _26520_ (.A1(_10048_),
    .A2(_11604_),
    .B1(_11605_),
    .B2(\datamem.data_ram[45][0] ),
    .X(_03204_));
 sky130_fd_sc_hd__a22o_1 _26521_ (.A1(_10058_),
    .A2(_11604_),
    .B1(_11605_),
    .B2(\datamem.data_ram[45][1] ),
    .X(_03205_));
 sky130_fd_sc_hd__a22o_1 _26522_ (.A1(_10061_),
    .A2(_11604_),
    .B1(_11605_),
    .B2(\datamem.data_ram[45][2] ),
    .X(_03206_));
 sky130_fd_sc_hd__a22o_1 _26523_ (.A1(_10064_),
    .A2(_11604_),
    .B1(_11605_),
    .B2(\datamem.data_ram[45][3] ),
    .X(_03207_));
 sky130_fd_sc_hd__a22o_1 _26524_ (.A1(_10782_),
    .A2(_11604_),
    .B1(_11605_),
    .B2(\datamem.data_ram[45][4] ),
    .X(_03208_));
 sky130_fd_sc_hd__a22o_1 _26525_ (.A1(_10070_),
    .A2(_11604_),
    .B1(_11605_),
    .B2(\datamem.data_ram[45][5] ),
    .X(_03209_));
 sky130_fd_sc_hd__a22o_1 _26526_ (.A1(_10073_),
    .A2(_11604_),
    .B1(_11605_),
    .B2(\datamem.data_ram[45][6] ),
    .X(_03210_));
 sky130_fd_sc_hd__a22o_1 _26527_ (.A1(_10783_),
    .A2(_11604_),
    .B1(_11605_),
    .B2(\datamem.data_ram[45][7] ),
    .X(_03211_));
 sky130_fd_sc_hd__a211o_1 _26528_ (.A1(_11374_),
    .A2(_06567_),
    .B1(_11367_),
    .C1(_11375_),
    .X(_11606_));
 sky130_fd_sc_hd__a21o_1 _26529_ (.A1(_11372_),
    .A2(_11606_),
    .B1(_02993_),
    .X(_03212_));
 sky130_fd_sc_hd__or3_1 _26530_ (.A(_07203_),
    .B(_10946_),
    .C(_11494_),
    .X(_11607_));
 sky130_fd_sc_hd__clkbuf_2 _26531_ (.A(_11607_),
    .X(_11608_));
 sky130_fd_sc_hd__clkbuf_4 _26532_ (.A(_10051_),
    .X(_11609_));
 sky130_fd_sc_hd__and3_1 _26533_ (.A(_10209_),
    .B(_11054_),
    .C(_11609_),
    .X(_11610_));
 sky130_fd_sc_hd__and2_1 _26534_ (.A(_11078_),
    .B(_11610_),
    .X(_11611_));
 sky130_fd_sc_hd__a31o_1 _26535_ (.A1(_11517_),
    .A2(\datamem.data_ram[18][0] ),
    .A3(_11608_),
    .B1(_11611_),
    .X(_03213_));
 sky130_fd_sc_hd__and2_1 _26536_ (.A(_11081_),
    .B(_11610_),
    .X(_11612_));
 sky130_fd_sc_hd__a31o_1 _26537_ (.A1(_11517_),
    .A2(\datamem.data_ram[18][1] ),
    .A3(_11608_),
    .B1(_11612_),
    .X(_03214_));
 sky130_fd_sc_hd__and2_1 _26538_ (.A(_11083_),
    .B(_11610_),
    .X(_11613_));
 sky130_fd_sc_hd__a31o_1 _26539_ (.A1(_11517_),
    .A2(\datamem.data_ram[18][2] ),
    .A3(_11608_),
    .B1(_11613_),
    .X(_03215_));
 sky130_fd_sc_hd__and2_1 _26540_ (.A(_11086_),
    .B(_11610_),
    .X(_11614_));
 sky130_fd_sc_hd__a31o_1 _26541_ (.A1(_11517_),
    .A2(\datamem.data_ram[18][3] ),
    .A3(_11608_),
    .B1(_11614_),
    .X(_03216_));
 sky130_fd_sc_hd__and2_1 _26542_ (.A(_11047_),
    .B(_11610_),
    .X(_11615_));
 sky130_fd_sc_hd__a31o_1 _26543_ (.A1(_11517_),
    .A2(\datamem.data_ram[18][4] ),
    .A3(_11608_),
    .B1(_11615_),
    .X(_03217_));
 sky130_fd_sc_hd__and2_1 _26544_ (.A(_11089_),
    .B(_11610_),
    .X(_11616_));
 sky130_fd_sc_hd__a31o_1 _26545_ (.A1(_11517_),
    .A2(\datamem.data_ram[18][5] ),
    .A3(_11608_),
    .B1(_11616_),
    .X(_03218_));
 sky130_fd_sc_hd__and2_1 _26546_ (.A(_11091_),
    .B(_11610_),
    .X(_11617_));
 sky130_fd_sc_hd__a31o_1 _26547_ (.A1(_11517_),
    .A2(\datamem.data_ram[18][6] ),
    .A3(_11608_),
    .B1(_11617_),
    .X(_03219_));
 sky130_fd_sc_hd__clkbuf_4 _26548_ (.A(_11104_),
    .X(_11618_));
 sky130_fd_sc_hd__and2_1 _26549_ (.A(_11064_),
    .B(_11610_),
    .X(_11619_));
 sky130_fd_sc_hd__a31o_1 _26550_ (.A1(_11618_),
    .A2(\datamem.data_ram[18][7] ),
    .A3(_11608_),
    .B1(_11619_),
    .X(_03220_));
 sky130_fd_sc_hd__a21oi_4 _26551_ (.A1(_10570_),
    .A2(_11123_),
    .B1(_10998_),
    .Y(_11620_));
 sky130_fd_sc_hd__mux2_1 _26552_ (.A0(_10811_),
    .A1(\datamem.data_ram[1][24] ),
    .S(_11620_),
    .X(_11621_));
 sky130_fd_sc_hd__clkbuf_1 _26553_ (.A(_11621_),
    .X(_03221_));
 sky130_fd_sc_hd__mux2_1 _26554_ (.A0(_10814_),
    .A1(\datamem.data_ram[1][25] ),
    .S(_11620_),
    .X(_11622_));
 sky130_fd_sc_hd__clkbuf_1 _26555_ (.A(_11622_),
    .X(_03222_));
 sky130_fd_sc_hd__mux2_1 _26556_ (.A0(_10816_),
    .A1(\datamem.data_ram[1][26] ),
    .S(_11620_),
    .X(_11623_));
 sky130_fd_sc_hd__clkbuf_1 _26557_ (.A(_11623_),
    .X(_03223_));
 sky130_fd_sc_hd__mux2_1 _26558_ (.A0(_10818_),
    .A1(\datamem.data_ram[1][27] ),
    .S(_11620_),
    .X(_11624_));
 sky130_fd_sc_hd__clkbuf_1 _26559_ (.A(_11624_),
    .X(_03224_));
 sky130_fd_sc_hd__mux2_1 _26560_ (.A0(_10820_),
    .A1(\datamem.data_ram[1][28] ),
    .S(_11620_),
    .X(_11625_));
 sky130_fd_sc_hd__clkbuf_1 _26561_ (.A(_11625_),
    .X(_03225_));
 sky130_fd_sc_hd__mux2_1 _26562_ (.A0(_10822_),
    .A1(\datamem.data_ram[1][29] ),
    .S(_11620_),
    .X(_11626_));
 sky130_fd_sc_hd__clkbuf_1 _26563_ (.A(_11626_),
    .X(_03226_));
 sky130_fd_sc_hd__mux2_1 _26564_ (.A0(_10824_),
    .A1(\datamem.data_ram[1][30] ),
    .S(_11620_),
    .X(_11627_));
 sky130_fd_sc_hd__clkbuf_1 _26565_ (.A(_11627_),
    .X(_03227_));
 sky130_fd_sc_hd__mux2_1 _26566_ (.A0(_10826_),
    .A1(\datamem.data_ram[1][31] ),
    .S(_11620_),
    .X(_11628_));
 sky130_fd_sc_hd__clkbuf_1 _26567_ (.A(_11628_),
    .X(_03228_));
 sky130_fd_sc_hd__a21oi_4 _26568_ (.A1(_10668_),
    .A2(_10092_),
    .B1(_10998_),
    .Y(_11629_));
 sky130_fd_sc_hd__mux2_1 _26569_ (.A0(_10724_),
    .A1(\datamem.data_ram[6][8] ),
    .S(_11629_),
    .X(_11630_));
 sky130_fd_sc_hd__clkbuf_1 _26570_ (.A(_11630_),
    .X(_03229_));
 sky130_fd_sc_hd__mux2_1 _26571_ (.A0(_10727_),
    .A1(\datamem.data_ram[6][9] ),
    .S(_11629_),
    .X(_11631_));
 sky130_fd_sc_hd__clkbuf_1 _26572_ (.A(_11631_),
    .X(_03230_));
 sky130_fd_sc_hd__mux2_1 _26573_ (.A0(_10729_),
    .A1(\datamem.data_ram[6][10] ),
    .S(_11629_),
    .X(_11632_));
 sky130_fd_sc_hd__clkbuf_1 _26574_ (.A(_11632_),
    .X(_03231_));
 sky130_fd_sc_hd__mux2_1 _26575_ (.A0(_10731_),
    .A1(\datamem.data_ram[6][11] ),
    .S(_11629_),
    .X(_11633_));
 sky130_fd_sc_hd__clkbuf_1 _26576_ (.A(_11633_),
    .X(_03232_));
 sky130_fd_sc_hd__mux2_1 _26577_ (.A0(_10733_),
    .A1(\datamem.data_ram[6][12] ),
    .S(_11629_),
    .X(_11634_));
 sky130_fd_sc_hd__clkbuf_1 _26578_ (.A(_11634_),
    .X(_03233_));
 sky130_fd_sc_hd__mux2_1 _26579_ (.A0(_10735_),
    .A1(\datamem.data_ram[6][13] ),
    .S(_11629_),
    .X(_11635_));
 sky130_fd_sc_hd__clkbuf_1 _26580_ (.A(_11635_),
    .X(_03234_));
 sky130_fd_sc_hd__mux2_1 _26581_ (.A0(_10737_),
    .A1(\datamem.data_ram[6][14] ),
    .S(_11629_),
    .X(_11636_));
 sky130_fd_sc_hd__clkbuf_1 _26582_ (.A(_11636_),
    .X(_03235_));
 sky130_fd_sc_hd__mux2_1 _26583_ (.A0(_10739_),
    .A1(\datamem.data_ram[6][15] ),
    .S(_11629_),
    .X(_11637_));
 sky130_fd_sc_hd__clkbuf_1 _26584_ (.A(_11637_),
    .X(_03236_));
 sky130_fd_sc_hd__or3_1 _26585_ (.A(_07191_),
    .B(_10932_),
    .C(_11494_),
    .X(_11638_));
 sky130_fd_sc_hd__buf_2 _26586_ (.A(_11638_),
    .X(_11639_));
 sky130_fd_sc_hd__and3_2 _26587_ (.A(_10297_),
    .B(_10935_),
    .C(_11609_),
    .X(_11640_));
 sky130_fd_sc_hd__and2_1 _26588_ (.A(_11078_),
    .B(_11640_),
    .X(_11641_));
 sky130_fd_sc_hd__a31o_1 _26589_ (.A1(_11618_),
    .A2(\datamem.data_ram[8][0] ),
    .A3(_11639_),
    .B1(_11641_),
    .X(_03237_));
 sky130_fd_sc_hd__and2_1 _26590_ (.A(_11081_),
    .B(_11640_),
    .X(_11642_));
 sky130_fd_sc_hd__a31o_1 _26591_ (.A1(_11618_),
    .A2(\datamem.data_ram[8][1] ),
    .A3(_11639_),
    .B1(_11642_),
    .X(_03238_));
 sky130_fd_sc_hd__and2_1 _26592_ (.A(_11083_),
    .B(_11640_),
    .X(_11643_));
 sky130_fd_sc_hd__a31o_1 _26593_ (.A1(_11618_),
    .A2(\datamem.data_ram[8][2] ),
    .A3(_11639_),
    .B1(_11643_),
    .X(_03239_));
 sky130_fd_sc_hd__and2_1 _26594_ (.A(_11086_),
    .B(_11640_),
    .X(_11644_));
 sky130_fd_sc_hd__a31o_1 _26595_ (.A1(_11618_),
    .A2(\datamem.data_ram[8][3] ),
    .A3(_11639_),
    .B1(_11644_),
    .X(_03240_));
 sky130_fd_sc_hd__clkbuf_4 _26596_ (.A(_10066_),
    .X(_11645_));
 sky130_fd_sc_hd__and2_1 _26597_ (.A(_11645_),
    .B(_11640_),
    .X(_11646_));
 sky130_fd_sc_hd__a31o_1 _26598_ (.A1(_11618_),
    .A2(\datamem.data_ram[8][4] ),
    .A3(_11639_),
    .B1(_11646_),
    .X(_03241_));
 sky130_fd_sc_hd__and2_1 _26599_ (.A(_11089_),
    .B(_11640_),
    .X(_11647_));
 sky130_fd_sc_hd__a31o_1 _26600_ (.A1(_11618_),
    .A2(\datamem.data_ram[8][5] ),
    .A3(_11639_),
    .B1(_11647_),
    .X(_03242_));
 sky130_fd_sc_hd__and2_1 _26601_ (.A(_11091_),
    .B(_11640_),
    .X(_11648_));
 sky130_fd_sc_hd__a31o_1 _26602_ (.A1(_11618_),
    .A2(\datamem.data_ram[8][6] ),
    .A3(_11639_),
    .B1(_11648_),
    .X(_03243_));
 sky130_fd_sc_hd__and2_1 _26603_ (.A(_11064_),
    .B(_11640_),
    .X(_11649_));
 sky130_fd_sc_hd__a31o_1 _26604_ (.A1(_11618_),
    .A2(\datamem.data_ram[8][7] ),
    .A3(_11639_),
    .B1(_11649_),
    .X(_03244_));
 sky130_fd_sc_hd__a21oi_4 _26605_ (.A1(_10520_),
    .A2(_11123_),
    .B1(_10998_),
    .Y(_11650_));
 sky130_fd_sc_hd__mux2_1 _26606_ (.A0(_10811_),
    .A1(\datamem.data_ram[2][24] ),
    .S(_11650_),
    .X(_11651_));
 sky130_fd_sc_hd__clkbuf_1 _26607_ (.A(_11651_),
    .X(_03245_));
 sky130_fd_sc_hd__mux2_1 _26608_ (.A0(_10814_),
    .A1(\datamem.data_ram[2][25] ),
    .S(_11650_),
    .X(_11652_));
 sky130_fd_sc_hd__clkbuf_1 _26609_ (.A(_11652_),
    .X(_03246_));
 sky130_fd_sc_hd__mux2_1 _26610_ (.A0(_10816_),
    .A1(\datamem.data_ram[2][26] ),
    .S(_11650_),
    .X(_11653_));
 sky130_fd_sc_hd__clkbuf_1 _26611_ (.A(_11653_),
    .X(_03247_));
 sky130_fd_sc_hd__mux2_1 _26612_ (.A0(_10818_),
    .A1(\datamem.data_ram[2][27] ),
    .S(_11650_),
    .X(_11654_));
 sky130_fd_sc_hd__clkbuf_1 _26613_ (.A(_11654_),
    .X(_03248_));
 sky130_fd_sc_hd__mux2_1 _26614_ (.A0(_10820_),
    .A1(\datamem.data_ram[2][28] ),
    .S(_11650_),
    .X(_11655_));
 sky130_fd_sc_hd__clkbuf_1 _26615_ (.A(_11655_),
    .X(_03249_));
 sky130_fd_sc_hd__mux2_1 _26616_ (.A0(_10822_),
    .A1(\datamem.data_ram[2][29] ),
    .S(_11650_),
    .X(_11656_));
 sky130_fd_sc_hd__clkbuf_1 _26617_ (.A(_11656_),
    .X(_03250_));
 sky130_fd_sc_hd__mux2_1 _26618_ (.A0(_10824_),
    .A1(\datamem.data_ram[2][30] ),
    .S(_11650_),
    .X(_11657_));
 sky130_fd_sc_hd__clkbuf_1 _26619_ (.A(_11657_),
    .X(_03251_));
 sky130_fd_sc_hd__mux2_1 _26620_ (.A0(_10826_),
    .A1(\datamem.data_ram[2][31] ),
    .S(_11650_),
    .X(_11658_));
 sky130_fd_sc_hd__clkbuf_1 _26621_ (.A(_11658_),
    .X(_03252_));
 sky130_fd_sc_hd__nor2_4 _26622_ (.A(_10600_),
    .B(_10947_),
    .Y(_11659_));
 sky130_fd_sc_hd__nor2_2 _26623_ (.A(_09231_),
    .B(_11659_),
    .Y(_11660_));
 sky130_fd_sc_hd__a22o_1 _26624_ (.A1(_10048_),
    .A2(_11659_),
    .B1(_11660_),
    .B2(\datamem.data_ram[46][0] ),
    .X(_03253_));
 sky130_fd_sc_hd__a22o_1 _26625_ (.A1(_10058_),
    .A2(_11659_),
    .B1(_11660_),
    .B2(\datamem.data_ram[46][1] ),
    .X(_03254_));
 sky130_fd_sc_hd__a22o_1 _26626_ (.A1(_10061_),
    .A2(_11659_),
    .B1(_11660_),
    .B2(\datamem.data_ram[46][2] ),
    .X(_03255_));
 sky130_fd_sc_hd__a22o_1 _26627_ (.A1(_10064_),
    .A2(_11659_),
    .B1(_11660_),
    .B2(\datamem.data_ram[46][3] ),
    .X(_03256_));
 sky130_fd_sc_hd__a22o_1 _26628_ (.A1(_10782_),
    .A2(_11659_),
    .B1(_11660_),
    .B2(\datamem.data_ram[46][4] ),
    .X(_03257_));
 sky130_fd_sc_hd__a22o_1 _26629_ (.A1(_10070_),
    .A2(_11659_),
    .B1(_11660_),
    .B2(\datamem.data_ram[46][5] ),
    .X(_03258_));
 sky130_fd_sc_hd__a22o_1 _26630_ (.A1(_10073_),
    .A2(_11659_),
    .B1(_11660_),
    .B2(\datamem.data_ram[46][6] ),
    .X(_03259_));
 sky130_fd_sc_hd__a22o_1 _26631_ (.A1(_10783_),
    .A2(_11659_),
    .B1(_11660_),
    .B2(\datamem.data_ram[46][7] ),
    .X(_03260_));
 sky130_fd_sc_hd__or3_1 _26632_ (.A(_07808_),
    .B(_10946_),
    .C(_11494_),
    .X(_11661_));
 sky130_fd_sc_hd__clkbuf_2 _26633_ (.A(_11661_),
    .X(_11662_));
 sky130_fd_sc_hd__and3_1 _26634_ (.A(_10268_),
    .B(_11054_),
    .C(_11609_),
    .X(_11663_));
 sky130_fd_sc_hd__and2_1 _26635_ (.A(_11078_),
    .B(_11663_),
    .X(_11664_));
 sky130_fd_sc_hd__a31o_1 _26636_ (.A1(_11618_),
    .A2(\datamem.data_ram[17][0] ),
    .A3(_11662_),
    .B1(_11664_),
    .X(_03261_));
 sky130_fd_sc_hd__buf_2 _26637_ (.A(_11104_),
    .X(_11665_));
 sky130_fd_sc_hd__and2_1 _26638_ (.A(_11081_),
    .B(_11663_),
    .X(_11666_));
 sky130_fd_sc_hd__a31o_1 _26639_ (.A1(_11665_),
    .A2(\datamem.data_ram[17][1] ),
    .A3(_11662_),
    .B1(_11666_),
    .X(_03262_));
 sky130_fd_sc_hd__and2_1 _26640_ (.A(_11083_),
    .B(_11663_),
    .X(_11667_));
 sky130_fd_sc_hd__a31o_1 _26641_ (.A1(_11665_),
    .A2(\datamem.data_ram[17][2] ),
    .A3(_11662_),
    .B1(_11667_),
    .X(_03263_));
 sky130_fd_sc_hd__and2_1 _26642_ (.A(_11086_),
    .B(_11663_),
    .X(_11668_));
 sky130_fd_sc_hd__a31o_1 _26643_ (.A1(_11665_),
    .A2(\datamem.data_ram[17][3] ),
    .A3(_11662_),
    .B1(_11668_),
    .X(_03264_));
 sky130_fd_sc_hd__and2_1 _26644_ (.A(_11645_),
    .B(_11663_),
    .X(_11669_));
 sky130_fd_sc_hd__a31o_1 _26645_ (.A1(_11665_),
    .A2(\datamem.data_ram[17][4] ),
    .A3(_11662_),
    .B1(_11669_),
    .X(_03265_));
 sky130_fd_sc_hd__and2_1 _26646_ (.A(_11089_),
    .B(_11663_),
    .X(_11670_));
 sky130_fd_sc_hd__a31o_1 _26647_ (.A1(_11665_),
    .A2(\datamem.data_ram[17][5] ),
    .A3(_11662_),
    .B1(_11670_),
    .X(_03266_));
 sky130_fd_sc_hd__and2_1 _26648_ (.A(_11091_),
    .B(_11663_),
    .X(_11671_));
 sky130_fd_sc_hd__a31o_1 _26649_ (.A1(_11665_),
    .A2(\datamem.data_ram[17][6] ),
    .A3(_11662_),
    .B1(_11671_),
    .X(_03267_));
 sky130_fd_sc_hd__buf_2 _26650_ (.A(_10075_),
    .X(_11672_));
 sky130_fd_sc_hd__and2_1 _26651_ (.A(_11672_),
    .B(_11663_),
    .X(_11673_));
 sky130_fd_sc_hd__a31o_1 _26652_ (.A1(_11665_),
    .A2(\datamem.data_ram[17][7] ),
    .A3(_11662_),
    .B1(_11673_),
    .X(_03268_));
 sky130_fd_sc_hd__or3_1 _26653_ (.A(_07808_),
    .B(_10932_),
    .C(_11494_),
    .X(_11674_));
 sky130_fd_sc_hd__clkbuf_2 _26654_ (.A(_11674_),
    .X(_11675_));
 sky130_fd_sc_hd__buf_2 _26655_ (.A(_10047_),
    .X(_11676_));
 sky130_fd_sc_hd__and3_2 _26656_ (.A(_10268_),
    .B(_10935_),
    .C(_11609_),
    .X(_11677_));
 sky130_fd_sc_hd__and2_1 _26657_ (.A(_11676_),
    .B(_11677_),
    .X(_11678_));
 sky130_fd_sc_hd__a31o_1 _26658_ (.A1(_11665_),
    .A2(\datamem.data_ram[9][0] ),
    .A3(_11675_),
    .B1(_11678_),
    .X(_03269_));
 sky130_fd_sc_hd__buf_2 _26659_ (.A(_10057_),
    .X(_11679_));
 sky130_fd_sc_hd__and2_1 _26660_ (.A(_11679_),
    .B(_11677_),
    .X(_11680_));
 sky130_fd_sc_hd__a31o_1 _26661_ (.A1(_11665_),
    .A2(\datamem.data_ram[9][1] ),
    .A3(_11675_),
    .B1(_11680_),
    .X(_03270_));
 sky130_fd_sc_hd__clkbuf_4 _26662_ (.A(_10060_),
    .X(_11681_));
 sky130_fd_sc_hd__and2_1 _26663_ (.A(_11681_),
    .B(_11677_),
    .X(_11682_));
 sky130_fd_sc_hd__a31o_1 _26664_ (.A1(_11665_),
    .A2(\datamem.data_ram[9][2] ),
    .A3(_11675_),
    .B1(_11682_),
    .X(_03271_));
 sky130_fd_sc_hd__buf_2 _26665_ (.A(_11104_),
    .X(_11683_));
 sky130_fd_sc_hd__buf_2 _26666_ (.A(_10063_),
    .X(_11684_));
 sky130_fd_sc_hd__and2_1 _26667_ (.A(_11684_),
    .B(_11677_),
    .X(_11685_));
 sky130_fd_sc_hd__a31o_1 _26668_ (.A1(_11683_),
    .A2(\datamem.data_ram[9][3] ),
    .A3(_11675_),
    .B1(_11685_),
    .X(_03272_));
 sky130_fd_sc_hd__and2_1 _26669_ (.A(_11645_),
    .B(_11677_),
    .X(_11686_));
 sky130_fd_sc_hd__a31o_1 _26670_ (.A1(_11683_),
    .A2(\datamem.data_ram[9][4] ),
    .A3(_11675_),
    .B1(_11686_),
    .X(_03273_));
 sky130_fd_sc_hd__buf_2 _26671_ (.A(_10069_),
    .X(_11687_));
 sky130_fd_sc_hd__and2_1 _26672_ (.A(_11687_),
    .B(_11677_),
    .X(_11688_));
 sky130_fd_sc_hd__a31o_1 _26673_ (.A1(_11683_),
    .A2(\datamem.data_ram[9][5] ),
    .A3(_11675_),
    .B1(_11688_),
    .X(_03274_));
 sky130_fd_sc_hd__buf_2 _26674_ (.A(_10072_),
    .X(_11689_));
 sky130_fd_sc_hd__and2_1 _26675_ (.A(_11689_),
    .B(_11677_),
    .X(_11690_));
 sky130_fd_sc_hd__a31o_1 _26676_ (.A1(_11683_),
    .A2(\datamem.data_ram[9][6] ),
    .A3(_11675_),
    .B1(_11690_),
    .X(_03275_));
 sky130_fd_sc_hd__and2_1 _26677_ (.A(_11672_),
    .B(_11677_),
    .X(_11691_));
 sky130_fd_sc_hd__a31o_1 _26678_ (.A1(_11683_),
    .A2(\datamem.data_ram[9][7] ),
    .A3(_11675_),
    .B1(_11691_),
    .X(_03276_));
 sky130_fd_sc_hd__or3_1 _26679_ (.A(_07191_),
    .B(_10946_),
    .C(_11494_),
    .X(_11692_));
 sky130_fd_sc_hd__clkbuf_2 _26680_ (.A(_11692_),
    .X(_11693_));
 sky130_fd_sc_hd__and3_1 _26681_ (.A(_10297_),
    .B(_11054_),
    .C(_11609_),
    .X(_11694_));
 sky130_fd_sc_hd__and2_1 _26682_ (.A(_11676_),
    .B(_11694_),
    .X(_11695_));
 sky130_fd_sc_hd__a31o_1 _26683_ (.A1(_11683_),
    .A2(\datamem.data_ram[16][0] ),
    .A3(_11693_),
    .B1(_11695_),
    .X(_03277_));
 sky130_fd_sc_hd__and2_1 _26684_ (.A(_11679_),
    .B(_11694_),
    .X(_11696_));
 sky130_fd_sc_hd__a31o_1 _26685_ (.A1(_11683_),
    .A2(\datamem.data_ram[16][1] ),
    .A3(_11693_),
    .B1(_11696_),
    .X(_03278_));
 sky130_fd_sc_hd__and2_1 _26686_ (.A(_11681_),
    .B(_11694_),
    .X(_11697_));
 sky130_fd_sc_hd__a31o_1 _26687_ (.A1(_11683_),
    .A2(\datamem.data_ram[16][2] ),
    .A3(_11693_),
    .B1(_11697_),
    .X(_03279_));
 sky130_fd_sc_hd__and2_1 _26688_ (.A(_11684_),
    .B(_11694_),
    .X(_11698_));
 sky130_fd_sc_hd__a31o_1 _26689_ (.A1(_11683_),
    .A2(\datamem.data_ram[16][3] ),
    .A3(_11693_),
    .B1(_11698_),
    .X(_03280_));
 sky130_fd_sc_hd__and2_1 _26690_ (.A(_11645_),
    .B(_11694_),
    .X(_11699_));
 sky130_fd_sc_hd__a31o_1 _26691_ (.A1(_11683_),
    .A2(\datamem.data_ram[16][4] ),
    .A3(_11693_),
    .B1(_11699_),
    .X(_03281_));
 sky130_fd_sc_hd__clkbuf_4 _26692_ (.A(_11104_),
    .X(_11700_));
 sky130_fd_sc_hd__and2_1 _26693_ (.A(_11687_),
    .B(_11694_),
    .X(_11701_));
 sky130_fd_sc_hd__a31o_1 _26694_ (.A1(_11700_),
    .A2(\datamem.data_ram[16][5] ),
    .A3(_11693_),
    .B1(_11701_),
    .X(_03282_));
 sky130_fd_sc_hd__and2_1 _26695_ (.A(_11689_),
    .B(_11694_),
    .X(_11702_));
 sky130_fd_sc_hd__a31o_1 _26696_ (.A1(_11700_),
    .A2(\datamem.data_ram[16][6] ),
    .A3(_11693_),
    .B1(_11702_),
    .X(_03283_));
 sky130_fd_sc_hd__and2_1 _26697_ (.A(_11672_),
    .B(_11694_),
    .X(_11703_));
 sky130_fd_sc_hd__a31o_1 _26698_ (.A1(_11700_),
    .A2(\datamem.data_ram[16][7] ),
    .A3(_11693_),
    .B1(_11703_),
    .X(_03284_));
 sky130_fd_sc_hd__a21oi_4 _26699_ (.A1(_10741_),
    .A2(_11123_),
    .B1(_10998_),
    .Y(_11704_));
 sky130_fd_sc_hd__mux2_1 _26700_ (.A0(_10811_),
    .A1(\datamem.data_ram[3][24] ),
    .S(_11704_),
    .X(_11705_));
 sky130_fd_sc_hd__clkbuf_1 _26701_ (.A(_11705_),
    .X(_03285_));
 sky130_fd_sc_hd__mux2_1 _26702_ (.A0(_10814_),
    .A1(\datamem.data_ram[3][25] ),
    .S(_11704_),
    .X(_11706_));
 sky130_fd_sc_hd__clkbuf_1 _26703_ (.A(_11706_),
    .X(_03286_));
 sky130_fd_sc_hd__mux2_1 _26704_ (.A0(_10816_),
    .A1(\datamem.data_ram[3][26] ),
    .S(_11704_),
    .X(_11707_));
 sky130_fd_sc_hd__clkbuf_1 _26705_ (.A(_11707_),
    .X(_03287_));
 sky130_fd_sc_hd__mux2_1 _26706_ (.A0(_10818_),
    .A1(\datamem.data_ram[3][27] ),
    .S(_11704_),
    .X(_11708_));
 sky130_fd_sc_hd__clkbuf_1 _26707_ (.A(_11708_),
    .X(_03288_));
 sky130_fd_sc_hd__mux2_1 _26708_ (.A0(_10820_),
    .A1(\datamem.data_ram[3][28] ),
    .S(_11704_),
    .X(_11709_));
 sky130_fd_sc_hd__clkbuf_1 _26709_ (.A(_11709_),
    .X(_03289_));
 sky130_fd_sc_hd__mux2_1 _26710_ (.A0(_10822_),
    .A1(\datamem.data_ram[3][29] ),
    .S(_11704_),
    .X(_11710_));
 sky130_fd_sc_hd__clkbuf_1 _26711_ (.A(_11710_),
    .X(_03290_));
 sky130_fd_sc_hd__mux2_1 _26712_ (.A0(_10824_),
    .A1(\datamem.data_ram[3][30] ),
    .S(_11704_),
    .X(_11711_));
 sky130_fd_sc_hd__clkbuf_1 _26713_ (.A(_11711_),
    .X(_03291_));
 sky130_fd_sc_hd__mux2_1 _26714_ (.A0(_10826_),
    .A1(\datamem.data_ram[3][31] ),
    .S(_11704_),
    .X(_11712_));
 sky130_fd_sc_hd__clkbuf_1 _26715_ (.A(_11712_),
    .X(_03292_));
 sky130_fd_sc_hd__buf_8 _26716_ (.A(_10500_),
    .X(_11713_));
 sky130_fd_sc_hd__a21oi_4 _26717_ (.A1(_10838_),
    .A2(_10960_),
    .B1(_11713_),
    .Y(_11714_));
 sky130_fd_sc_hd__mux2_1 _26718_ (.A0(_10751_),
    .A1(\datamem.data_ram[8][16] ),
    .S(_11714_),
    .X(_11715_));
 sky130_fd_sc_hd__clkbuf_1 _26719_ (.A(_11715_),
    .X(_03293_));
 sky130_fd_sc_hd__mux2_1 _26720_ (.A0(_10754_),
    .A1(\datamem.data_ram[8][17] ),
    .S(_11714_),
    .X(_11716_));
 sky130_fd_sc_hd__clkbuf_1 _26721_ (.A(_11716_),
    .X(_03294_));
 sky130_fd_sc_hd__mux2_1 _26722_ (.A0(_10756_),
    .A1(\datamem.data_ram[8][18] ),
    .S(_11714_),
    .X(_11717_));
 sky130_fd_sc_hd__clkbuf_1 _26723_ (.A(_11717_),
    .X(_03295_));
 sky130_fd_sc_hd__mux2_1 _26724_ (.A0(_10758_),
    .A1(\datamem.data_ram[8][19] ),
    .S(_11714_),
    .X(_11718_));
 sky130_fd_sc_hd__clkbuf_1 _26725_ (.A(_11718_),
    .X(_03296_));
 sky130_fd_sc_hd__mux2_1 _26726_ (.A0(_10760_),
    .A1(\datamem.data_ram[8][20] ),
    .S(_11714_),
    .X(_11719_));
 sky130_fd_sc_hd__clkbuf_1 _26727_ (.A(_11719_),
    .X(_03297_));
 sky130_fd_sc_hd__mux2_1 _26728_ (.A0(_10762_),
    .A1(\datamem.data_ram[8][21] ),
    .S(_11714_),
    .X(_11720_));
 sky130_fd_sc_hd__clkbuf_1 _26729_ (.A(_11720_),
    .X(_03298_));
 sky130_fd_sc_hd__mux2_1 _26730_ (.A0(_10764_),
    .A1(\datamem.data_ram[8][22] ),
    .S(_11714_),
    .X(_11721_));
 sky130_fd_sc_hd__clkbuf_1 _26731_ (.A(_11721_),
    .X(_03299_));
 sky130_fd_sc_hd__mux2_1 _26732_ (.A0(_10766_),
    .A1(\datamem.data_ram[8][23] ),
    .S(_11714_),
    .X(_11722_));
 sky130_fd_sc_hd__clkbuf_1 _26733_ (.A(_11722_),
    .X(_03300_));
 sky130_fd_sc_hd__or2_1 _26734_ (.A(_09227_),
    .B(_11603_),
    .X(_11723_));
 sky130_fd_sc_hd__clkbuf_4 _26735_ (.A(_11723_),
    .X(_11724_));
 sky130_fd_sc_hd__buf_2 _26736_ (.A(_09227_),
    .X(_11725_));
 sky130_fd_sc_hd__nor2_1 _26737_ (.A(_11725_),
    .B(_11603_),
    .Y(_11726_));
 sky130_fd_sc_hd__and2_1 _26738_ (.A(_11676_),
    .B(_11726_),
    .X(_11727_));
 sky130_fd_sc_hd__a31o_1 _26739_ (.A1(_11700_),
    .A2(\datamem.data_ram[61][0] ),
    .A3(_11724_),
    .B1(_11727_),
    .X(_03301_));
 sky130_fd_sc_hd__and2_1 _26740_ (.A(_11679_),
    .B(_11726_),
    .X(_11728_));
 sky130_fd_sc_hd__a31o_1 _26741_ (.A1(_11700_),
    .A2(\datamem.data_ram[61][1] ),
    .A3(_11724_),
    .B1(_11728_),
    .X(_03302_));
 sky130_fd_sc_hd__and2_1 _26742_ (.A(_11681_),
    .B(_11726_),
    .X(_11729_));
 sky130_fd_sc_hd__a31o_1 _26743_ (.A1(_11700_),
    .A2(\datamem.data_ram[61][2] ),
    .A3(_11724_),
    .B1(_11729_),
    .X(_03303_));
 sky130_fd_sc_hd__and2_1 _26744_ (.A(_11684_),
    .B(_11726_),
    .X(_11730_));
 sky130_fd_sc_hd__a31o_1 _26745_ (.A1(_11700_),
    .A2(\datamem.data_ram[61][3] ),
    .A3(_11724_),
    .B1(_11730_),
    .X(_03304_));
 sky130_fd_sc_hd__and2_1 _26746_ (.A(_11645_),
    .B(_11726_),
    .X(_11731_));
 sky130_fd_sc_hd__a31o_1 _26747_ (.A1(_11700_),
    .A2(\datamem.data_ram[61][4] ),
    .A3(_11724_),
    .B1(_11731_),
    .X(_03305_));
 sky130_fd_sc_hd__and2_1 _26748_ (.A(_11687_),
    .B(_11726_),
    .X(_11732_));
 sky130_fd_sc_hd__a31o_1 _26749_ (.A1(_11700_),
    .A2(\datamem.data_ram[61][5] ),
    .A3(_11724_),
    .B1(_11732_),
    .X(_03306_));
 sky130_fd_sc_hd__and2_1 _26750_ (.A(_11689_),
    .B(_11726_),
    .X(_11733_));
 sky130_fd_sc_hd__a31o_1 _26751_ (.A1(_11700_),
    .A2(\datamem.data_ram[61][6] ),
    .A3(_11724_),
    .B1(_11733_),
    .X(_03307_));
 sky130_fd_sc_hd__mux2_1 _26752_ (.A0(_10783_),
    .A1(_08356_),
    .S(_11724_),
    .X(_11734_));
 sky130_fd_sc_hd__clkbuf_1 _26753_ (.A(_11734_),
    .X(_03308_));
 sky130_fd_sc_hd__buf_2 _26754_ (.A(_11104_),
    .X(_11735_));
 sky130_fd_sc_hd__or2_1 _26755_ (.A(_11725_),
    .B(_10947_),
    .X(_11736_));
 sky130_fd_sc_hd__buf_2 _26756_ (.A(_11736_),
    .X(_11737_));
 sky130_fd_sc_hd__nor2_2 _26757_ (.A(_11725_),
    .B(_10947_),
    .Y(_11738_));
 sky130_fd_sc_hd__and2_1 _26758_ (.A(_11676_),
    .B(_11738_),
    .X(_11739_));
 sky130_fd_sc_hd__a31o_1 _26759_ (.A1(_11735_),
    .A2(\datamem.data_ram[62][0] ),
    .A3(_11737_),
    .B1(_11739_),
    .X(_03309_));
 sky130_fd_sc_hd__and2_1 _26760_ (.A(_11679_),
    .B(_11738_),
    .X(_11740_));
 sky130_fd_sc_hd__a31o_1 _26761_ (.A1(_11735_),
    .A2(\datamem.data_ram[62][1] ),
    .A3(_11737_),
    .B1(_11740_),
    .X(_03310_));
 sky130_fd_sc_hd__and2_1 _26762_ (.A(_11681_),
    .B(_11738_),
    .X(_11741_));
 sky130_fd_sc_hd__a31o_1 _26763_ (.A1(_11735_),
    .A2(\datamem.data_ram[62][2] ),
    .A3(_11737_),
    .B1(_11741_),
    .X(_03311_));
 sky130_fd_sc_hd__and2_1 _26764_ (.A(_11684_),
    .B(_11738_),
    .X(_11742_));
 sky130_fd_sc_hd__a31o_1 _26765_ (.A1(_11735_),
    .A2(\datamem.data_ram[62][3] ),
    .A3(_11737_),
    .B1(_11742_),
    .X(_03312_));
 sky130_fd_sc_hd__and2_1 _26766_ (.A(_11645_),
    .B(_11738_),
    .X(_11743_));
 sky130_fd_sc_hd__a31o_1 _26767_ (.A1(_11735_),
    .A2(\datamem.data_ram[62][4] ),
    .A3(_11737_),
    .B1(_11743_),
    .X(_03313_));
 sky130_fd_sc_hd__and2_1 _26768_ (.A(_11687_),
    .B(_11738_),
    .X(_11744_));
 sky130_fd_sc_hd__a31o_1 _26769_ (.A1(_11735_),
    .A2(\datamem.data_ram[62][5] ),
    .A3(_11737_),
    .B1(_11744_),
    .X(_03314_));
 sky130_fd_sc_hd__and2_1 _26770_ (.A(_11689_),
    .B(_11738_),
    .X(_11745_));
 sky130_fd_sc_hd__a31o_1 _26771_ (.A1(_11735_),
    .A2(\datamem.data_ram[62][6] ),
    .A3(_11737_),
    .B1(_11745_),
    .X(_03315_));
 sky130_fd_sc_hd__and2_1 _26772_ (.A(_11672_),
    .B(_11738_),
    .X(_11746_));
 sky130_fd_sc_hd__a31o_1 _26773_ (.A1(_11735_),
    .A2(\datamem.data_ram[62][7] ),
    .A3(_11737_),
    .B1(_11746_),
    .X(_03316_));
 sky130_fd_sc_hd__or3_1 _26774_ (.A(_07791_),
    .B(_11725_),
    .C(_11494_),
    .X(_11747_));
 sky130_fd_sc_hd__buf_2 _26775_ (.A(_11747_),
    .X(_11748_));
 sky130_fd_sc_hd__and3_2 _26776_ (.A(_10325_),
    .B(_08066_),
    .C(_11609_),
    .X(_11749_));
 sky130_fd_sc_hd__and2_1 _26777_ (.A(_11676_),
    .B(_11749_),
    .X(_11750_));
 sky130_fd_sc_hd__a31o_1 _26778_ (.A1(_11735_),
    .A2(\datamem.data_ram[63][0] ),
    .A3(_11748_),
    .B1(_11750_),
    .X(_03317_));
 sky130_fd_sc_hd__and2_1 _26779_ (.A(_11679_),
    .B(_11749_),
    .X(_11751_));
 sky130_fd_sc_hd__a31o_1 _26780_ (.A1(_11735_),
    .A2(\datamem.data_ram[63][1] ),
    .A3(_11748_),
    .B1(_11751_),
    .X(_03318_));
 sky130_fd_sc_hd__buf_2 _26781_ (.A(_06587_),
    .X(_11752_));
 sky130_fd_sc_hd__clkbuf_4 _26782_ (.A(_11752_),
    .X(_11753_));
 sky130_fd_sc_hd__and2_1 _26783_ (.A(_11681_),
    .B(_11749_),
    .X(_11754_));
 sky130_fd_sc_hd__a31o_1 _26784_ (.A1(_11753_),
    .A2(\datamem.data_ram[63][2] ),
    .A3(_11748_),
    .B1(_11754_),
    .X(_03319_));
 sky130_fd_sc_hd__and2_1 _26785_ (.A(_11684_),
    .B(_11749_),
    .X(_11755_));
 sky130_fd_sc_hd__a31o_1 _26786_ (.A1(_11753_),
    .A2(\datamem.data_ram[63][3] ),
    .A3(_11748_),
    .B1(_11755_),
    .X(_03320_));
 sky130_fd_sc_hd__and2_1 _26787_ (.A(_11645_),
    .B(_11749_),
    .X(_11756_));
 sky130_fd_sc_hd__a31o_1 _26788_ (.A1(_11753_),
    .A2(\datamem.data_ram[63][4] ),
    .A3(_11748_),
    .B1(_11756_),
    .X(_03321_));
 sky130_fd_sc_hd__and2_1 _26789_ (.A(_11687_),
    .B(_11749_),
    .X(_11757_));
 sky130_fd_sc_hd__a31o_1 _26790_ (.A1(_11753_),
    .A2(\datamem.data_ram[63][5] ),
    .A3(_11748_),
    .B1(_11757_),
    .X(_03322_));
 sky130_fd_sc_hd__and2_1 _26791_ (.A(_11689_),
    .B(_11749_),
    .X(_11758_));
 sky130_fd_sc_hd__a31o_1 _26792_ (.A1(_11753_),
    .A2(\datamem.data_ram[63][6] ),
    .A3(_11748_),
    .B1(_11758_),
    .X(_03323_));
 sky130_fd_sc_hd__and2_1 _26793_ (.A(_11672_),
    .B(_11749_),
    .X(_11759_));
 sky130_fd_sc_hd__a31o_1 _26794_ (.A1(_11753_),
    .A2(\datamem.data_ram[63][7] ),
    .A3(_11748_),
    .B1(_11759_),
    .X(_03324_));
 sky130_fd_sc_hd__or3_1 _26795_ (.A(_07191_),
    .B(_11725_),
    .C(_11494_),
    .X(_11760_));
 sky130_fd_sc_hd__buf_2 _26796_ (.A(_11760_),
    .X(_11761_));
 sky130_fd_sc_hd__and3_2 _26797_ (.A(_10297_),
    .B(_08066_),
    .C(_11609_),
    .X(_11762_));
 sky130_fd_sc_hd__and2_1 _26798_ (.A(_11676_),
    .B(_11762_),
    .X(_11763_));
 sky130_fd_sc_hd__a31o_1 _26799_ (.A1(_11753_),
    .A2(\datamem.data_ram[56][0] ),
    .A3(_11761_),
    .B1(_11763_),
    .X(_03325_));
 sky130_fd_sc_hd__and2_1 _26800_ (.A(_11679_),
    .B(_11762_),
    .X(_11764_));
 sky130_fd_sc_hd__a31o_1 _26801_ (.A1(_11753_),
    .A2(\datamem.data_ram[56][1] ),
    .A3(_11761_),
    .B1(_11764_),
    .X(_03326_));
 sky130_fd_sc_hd__and2_1 _26802_ (.A(_11681_),
    .B(_11762_),
    .X(_11765_));
 sky130_fd_sc_hd__a31o_1 _26803_ (.A1(_11753_),
    .A2(\datamem.data_ram[56][2] ),
    .A3(_11761_),
    .B1(_11765_),
    .X(_03327_));
 sky130_fd_sc_hd__and2_1 _26804_ (.A(_11684_),
    .B(_11762_),
    .X(_11766_));
 sky130_fd_sc_hd__a31o_1 _26805_ (.A1(_11753_),
    .A2(\datamem.data_ram[56][3] ),
    .A3(_11761_),
    .B1(_11766_),
    .X(_03328_));
 sky130_fd_sc_hd__buf_2 _26806_ (.A(_11752_),
    .X(_11767_));
 sky130_fd_sc_hd__and2_1 _26807_ (.A(_11645_),
    .B(_11762_),
    .X(_11768_));
 sky130_fd_sc_hd__a31o_1 _26808_ (.A1(_11767_),
    .A2(\datamem.data_ram[56][4] ),
    .A3(_11761_),
    .B1(_11768_),
    .X(_03329_));
 sky130_fd_sc_hd__and2_1 _26809_ (.A(_11687_),
    .B(_11762_),
    .X(_11769_));
 sky130_fd_sc_hd__a31o_1 _26810_ (.A1(_11767_),
    .A2(\datamem.data_ram[56][5] ),
    .A3(_11761_),
    .B1(_11769_),
    .X(_03330_));
 sky130_fd_sc_hd__and2_1 _26811_ (.A(_11689_),
    .B(_11762_),
    .X(_11770_));
 sky130_fd_sc_hd__a31o_1 _26812_ (.A1(_11767_),
    .A2(\datamem.data_ram[56][6] ),
    .A3(_11761_),
    .B1(_11770_),
    .X(_03331_));
 sky130_fd_sc_hd__and2_1 _26813_ (.A(_11672_),
    .B(_11762_),
    .X(_11771_));
 sky130_fd_sc_hd__a31o_1 _26814_ (.A1(_11767_),
    .A2(\datamem.data_ram[56][7] ),
    .A3(_11761_),
    .B1(_11771_),
    .X(_03332_));
 sky130_fd_sc_hd__or3_1 _26815_ (.A(_07808_),
    .B(_11725_),
    .C(_11494_),
    .X(_11772_));
 sky130_fd_sc_hd__buf_2 _26816_ (.A(_11772_),
    .X(_11773_));
 sky130_fd_sc_hd__and3_2 _26817_ (.A(_10268_),
    .B(_08066_),
    .C(_11609_),
    .X(_11774_));
 sky130_fd_sc_hd__and2_1 _26818_ (.A(_11676_),
    .B(_11774_),
    .X(_11775_));
 sky130_fd_sc_hd__a31o_1 _26819_ (.A1(_11767_),
    .A2(\datamem.data_ram[57][0] ),
    .A3(_11773_),
    .B1(_11775_),
    .X(_03333_));
 sky130_fd_sc_hd__and2_1 _26820_ (.A(_11679_),
    .B(_11774_),
    .X(_11776_));
 sky130_fd_sc_hd__a31o_1 _26821_ (.A1(_11767_),
    .A2(\datamem.data_ram[57][1] ),
    .A3(_11773_),
    .B1(_11776_),
    .X(_03334_));
 sky130_fd_sc_hd__and2_1 _26822_ (.A(_11681_),
    .B(_11774_),
    .X(_11777_));
 sky130_fd_sc_hd__a31o_1 _26823_ (.A1(_11767_),
    .A2(\datamem.data_ram[57][2] ),
    .A3(_11773_),
    .B1(_11777_),
    .X(_03335_));
 sky130_fd_sc_hd__and2_1 _26824_ (.A(_11684_),
    .B(_11774_),
    .X(_11778_));
 sky130_fd_sc_hd__a31o_1 _26825_ (.A1(_11767_),
    .A2(\datamem.data_ram[57][3] ),
    .A3(_11773_),
    .B1(_11778_),
    .X(_03336_));
 sky130_fd_sc_hd__and2_1 _26826_ (.A(_11645_),
    .B(_11774_),
    .X(_11779_));
 sky130_fd_sc_hd__a31o_1 _26827_ (.A1(_11767_),
    .A2(\datamem.data_ram[57][4] ),
    .A3(_11773_),
    .B1(_11779_),
    .X(_03337_));
 sky130_fd_sc_hd__and2_1 _26828_ (.A(_11687_),
    .B(_11774_),
    .X(_11780_));
 sky130_fd_sc_hd__a31o_1 _26829_ (.A1(_11767_),
    .A2(\datamem.data_ram[57][5] ),
    .A3(_11773_),
    .B1(_11780_),
    .X(_03338_));
 sky130_fd_sc_hd__buf_2 _26830_ (.A(_11752_),
    .X(_11781_));
 sky130_fd_sc_hd__and2_1 _26831_ (.A(_11689_),
    .B(_11774_),
    .X(_11782_));
 sky130_fd_sc_hd__a31o_1 _26832_ (.A1(_11781_),
    .A2(\datamem.data_ram[57][6] ),
    .A3(_11773_),
    .B1(_11782_),
    .X(_03339_));
 sky130_fd_sc_hd__and2_1 _26833_ (.A(_11672_),
    .B(_11774_),
    .X(_11783_));
 sky130_fd_sc_hd__a31o_1 _26834_ (.A1(_11781_),
    .A2(\datamem.data_ram[57][7] ),
    .A3(_11773_),
    .B1(_11783_),
    .X(_03340_));
 sky130_fd_sc_hd__or3_1 _26835_ (.A(_07182_),
    .B(_10918_),
    .C(_10897_),
    .X(_11784_));
 sky130_fd_sc_hd__clkbuf_2 _26836_ (.A(_11784_),
    .X(_11785_));
 sky130_fd_sc_hd__and3_1 _26837_ (.A(_09351_),
    .B(_10921_),
    .C(_10922_),
    .X(_11786_));
 sky130_fd_sc_hd__and2_1 _26838_ (.A(_11676_),
    .B(_11786_),
    .X(_11787_));
 sky130_fd_sc_hd__a31o_1 _26839_ (.A1(_11781_),
    .A2(\datamem.data_ram[36][0] ),
    .A3(_11785_),
    .B1(_11787_),
    .X(_03341_));
 sky130_fd_sc_hd__and2_1 _26840_ (.A(_11679_),
    .B(_11786_),
    .X(_11788_));
 sky130_fd_sc_hd__a31o_1 _26841_ (.A1(_11781_),
    .A2(\datamem.data_ram[36][1] ),
    .A3(_11785_),
    .B1(_11788_),
    .X(_03342_));
 sky130_fd_sc_hd__and2_1 _26842_ (.A(_11681_),
    .B(_11786_),
    .X(_11789_));
 sky130_fd_sc_hd__a31o_1 _26843_ (.A1(_11781_),
    .A2(\datamem.data_ram[36][2] ),
    .A3(_11785_),
    .B1(_11789_),
    .X(_03343_));
 sky130_fd_sc_hd__and2_1 _26844_ (.A(_11684_),
    .B(_11786_),
    .X(_11790_));
 sky130_fd_sc_hd__a31o_1 _26845_ (.A1(_11781_),
    .A2(\datamem.data_ram[36][3] ),
    .A3(_11785_),
    .B1(_11790_),
    .X(_03344_));
 sky130_fd_sc_hd__and2_1 _26846_ (.A(_11645_),
    .B(_11786_),
    .X(_11791_));
 sky130_fd_sc_hd__a31o_1 _26847_ (.A1(_11781_),
    .A2(\datamem.data_ram[36][4] ),
    .A3(_11785_),
    .B1(_11791_),
    .X(_03345_));
 sky130_fd_sc_hd__and2_1 _26848_ (.A(_11687_),
    .B(_11786_),
    .X(_11792_));
 sky130_fd_sc_hd__a31o_1 _26849_ (.A1(_11781_),
    .A2(\datamem.data_ram[36][5] ),
    .A3(_11785_),
    .B1(_11792_),
    .X(_03346_));
 sky130_fd_sc_hd__and2_1 _26850_ (.A(_11689_),
    .B(_11786_),
    .X(_11793_));
 sky130_fd_sc_hd__a31o_1 _26851_ (.A1(_11781_),
    .A2(\datamem.data_ram[36][6] ),
    .A3(_11785_),
    .B1(_11793_),
    .X(_03347_));
 sky130_fd_sc_hd__and2_1 _26852_ (.A(_11672_),
    .B(_11786_),
    .X(_11794_));
 sky130_fd_sc_hd__a31o_1 _26853_ (.A1(_11781_),
    .A2(\datamem.data_ram[36][7] ),
    .A3(_11785_),
    .B1(_11794_),
    .X(_03348_));
 sky130_fd_sc_hd__clkbuf_4 _26854_ (.A(_11752_),
    .X(_11795_));
 sky130_fd_sc_hd__or2_1 _26855_ (.A(_11725_),
    .B(_11039_),
    .X(_11796_));
 sky130_fd_sc_hd__buf_2 _26856_ (.A(_11796_),
    .X(_11797_));
 sky130_fd_sc_hd__nor2_2 _26857_ (.A(_11725_),
    .B(_11039_),
    .Y(_11798_));
 sky130_fd_sc_hd__and2_1 _26858_ (.A(_11676_),
    .B(_11798_),
    .X(_11799_));
 sky130_fd_sc_hd__a31o_1 _26859_ (.A1(_11795_),
    .A2(\datamem.data_ram[60][0] ),
    .A3(_11797_),
    .B1(_11799_),
    .X(_03349_));
 sky130_fd_sc_hd__and2_1 _26860_ (.A(_11679_),
    .B(_11798_),
    .X(_11800_));
 sky130_fd_sc_hd__a31o_1 _26861_ (.A1(_11795_),
    .A2(\datamem.data_ram[60][1] ),
    .A3(_11797_),
    .B1(_11800_),
    .X(_03350_));
 sky130_fd_sc_hd__and2_1 _26862_ (.A(_11681_),
    .B(_11798_),
    .X(_11801_));
 sky130_fd_sc_hd__a31o_1 _26863_ (.A1(_11795_),
    .A2(\datamem.data_ram[60][2] ),
    .A3(_11797_),
    .B1(_11801_),
    .X(_03351_));
 sky130_fd_sc_hd__and2_1 _26864_ (.A(_11684_),
    .B(_11798_),
    .X(_11802_));
 sky130_fd_sc_hd__a31o_1 _26865_ (.A1(_11795_),
    .A2(\datamem.data_ram[60][3] ),
    .A3(_11797_),
    .B1(_11802_),
    .X(_03352_));
 sky130_fd_sc_hd__clkbuf_4 _26866_ (.A(_10066_),
    .X(_11803_));
 sky130_fd_sc_hd__and2_1 _26867_ (.A(_11803_),
    .B(_11798_),
    .X(_11804_));
 sky130_fd_sc_hd__a31o_1 _26868_ (.A1(_11795_),
    .A2(\datamem.data_ram[60][4] ),
    .A3(_11797_),
    .B1(_11804_),
    .X(_03353_));
 sky130_fd_sc_hd__and2_1 _26869_ (.A(_11687_),
    .B(_11798_),
    .X(_11805_));
 sky130_fd_sc_hd__a31o_1 _26870_ (.A1(_11795_),
    .A2(\datamem.data_ram[60][5] ),
    .A3(_11797_),
    .B1(_11805_),
    .X(_03354_));
 sky130_fd_sc_hd__and2_1 _26871_ (.A(_11689_),
    .B(_11798_),
    .X(_11806_));
 sky130_fd_sc_hd__a31o_1 _26872_ (.A1(_11795_),
    .A2(\datamem.data_ram[60][6] ),
    .A3(_11797_),
    .B1(_11806_),
    .X(_03355_));
 sky130_fd_sc_hd__and2_1 _26873_ (.A(_11672_),
    .B(_11798_),
    .X(_11807_));
 sky130_fd_sc_hd__a31o_1 _26874_ (.A1(_11795_),
    .A2(\datamem.data_ram[60][7] ),
    .A3(_11797_),
    .B1(_11807_),
    .X(_03356_));
 sky130_fd_sc_hd__or2_1 _26875_ (.A(_11725_),
    .B(_11075_),
    .X(_11808_));
 sky130_fd_sc_hd__buf_2 _26876_ (.A(_11808_),
    .X(_11809_));
 sky130_fd_sc_hd__nor2_2 _26877_ (.A(_11725_),
    .B(_11075_),
    .Y(_11810_));
 sky130_fd_sc_hd__and2_1 _26878_ (.A(_11676_),
    .B(_11810_),
    .X(_11811_));
 sky130_fd_sc_hd__a31o_1 _26879_ (.A1(_11795_),
    .A2(\datamem.data_ram[59][0] ),
    .A3(_11809_),
    .B1(_11811_),
    .X(_03357_));
 sky130_fd_sc_hd__and2_1 _26880_ (.A(_11679_),
    .B(_11810_),
    .X(_11812_));
 sky130_fd_sc_hd__a31o_1 _26881_ (.A1(_11795_),
    .A2(\datamem.data_ram[59][1] ),
    .A3(_11809_),
    .B1(_11812_),
    .X(_03358_));
 sky130_fd_sc_hd__clkbuf_4 _26882_ (.A(_11752_),
    .X(_11813_));
 sky130_fd_sc_hd__and2_1 _26883_ (.A(_11681_),
    .B(_11810_),
    .X(_11814_));
 sky130_fd_sc_hd__a31o_1 _26884_ (.A1(_11813_),
    .A2(\datamem.data_ram[59][2] ),
    .A3(_11809_),
    .B1(_11814_),
    .X(_03359_));
 sky130_fd_sc_hd__and2_1 _26885_ (.A(_11684_),
    .B(_11810_),
    .X(_11815_));
 sky130_fd_sc_hd__a31o_1 _26886_ (.A1(_11813_),
    .A2(\datamem.data_ram[59][3] ),
    .A3(_11809_),
    .B1(_11815_),
    .X(_03360_));
 sky130_fd_sc_hd__and2_1 _26887_ (.A(_11803_),
    .B(_11810_),
    .X(_11816_));
 sky130_fd_sc_hd__a31o_1 _26888_ (.A1(_11813_),
    .A2(\datamem.data_ram[59][4] ),
    .A3(_11809_),
    .B1(_11816_),
    .X(_03361_));
 sky130_fd_sc_hd__and2_1 _26889_ (.A(_11687_),
    .B(_11810_),
    .X(_11817_));
 sky130_fd_sc_hd__a31o_1 _26890_ (.A1(_11813_),
    .A2(\datamem.data_ram[59][5] ),
    .A3(_11809_),
    .B1(_11817_),
    .X(_03362_));
 sky130_fd_sc_hd__and2_1 _26891_ (.A(_11689_),
    .B(_11810_),
    .X(_11818_));
 sky130_fd_sc_hd__a31o_1 _26892_ (.A1(_11813_),
    .A2(\datamem.data_ram[59][6] ),
    .A3(_11809_),
    .B1(_11818_),
    .X(_03363_));
 sky130_fd_sc_hd__and2_1 _26893_ (.A(_11672_),
    .B(_11810_),
    .X(_11819_));
 sky130_fd_sc_hd__a31o_1 _26894_ (.A1(_11813_),
    .A2(\datamem.data_ram[59][7] ),
    .A3(_11809_),
    .B1(_11819_),
    .X(_03364_));
 sky130_fd_sc_hd__or3_1 _26895_ (.A(_07191_),
    .B(_10918_),
    .C(_10897_),
    .X(_11820_));
 sky130_fd_sc_hd__buf_2 _26896_ (.A(_11820_),
    .X(_11821_));
 sky130_fd_sc_hd__clkbuf_4 _26897_ (.A(_10047_),
    .X(_11822_));
 sky130_fd_sc_hd__and3_2 _26898_ (.A(_10297_),
    .B(_10921_),
    .C(_10922_),
    .X(_11823_));
 sky130_fd_sc_hd__and2_1 _26899_ (.A(_11822_),
    .B(_11823_),
    .X(_11824_));
 sky130_fd_sc_hd__a31o_1 _26900_ (.A1(_11813_),
    .A2(\datamem.data_ram[32][0] ),
    .A3(_11821_),
    .B1(_11824_),
    .X(_03365_));
 sky130_fd_sc_hd__clkbuf_4 _26901_ (.A(_10057_),
    .X(_11825_));
 sky130_fd_sc_hd__and2_1 _26902_ (.A(_11825_),
    .B(_11823_),
    .X(_11826_));
 sky130_fd_sc_hd__a31o_1 _26903_ (.A1(_11813_),
    .A2(\datamem.data_ram[32][1] ),
    .A3(_11821_),
    .B1(_11826_),
    .X(_03366_));
 sky130_fd_sc_hd__clkbuf_4 _26904_ (.A(_10060_),
    .X(_11827_));
 sky130_fd_sc_hd__and2_1 _26905_ (.A(_11827_),
    .B(_11823_),
    .X(_11828_));
 sky130_fd_sc_hd__a31o_1 _26906_ (.A1(_11813_),
    .A2(\datamem.data_ram[32][2] ),
    .A3(_11821_),
    .B1(_11828_),
    .X(_03367_));
 sky130_fd_sc_hd__clkbuf_4 _26907_ (.A(_10063_),
    .X(_11829_));
 sky130_fd_sc_hd__and2_1 _26908_ (.A(_11829_),
    .B(_11823_),
    .X(_11830_));
 sky130_fd_sc_hd__a31o_1 _26909_ (.A1(_11813_),
    .A2(\datamem.data_ram[32][3] ),
    .A3(_11821_),
    .B1(_11830_),
    .X(_03368_));
 sky130_fd_sc_hd__clkbuf_4 _26910_ (.A(_11752_),
    .X(_11831_));
 sky130_fd_sc_hd__and2_1 _26911_ (.A(_11803_),
    .B(_11823_),
    .X(_11832_));
 sky130_fd_sc_hd__a31o_1 _26912_ (.A1(_11831_),
    .A2(\datamem.data_ram[32][4] ),
    .A3(_11821_),
    .B1(_11832_),
    .X(_03369_));
 sky130_fd_sc_hd__clkbuf_4 _26913_ (.A(_10069_),
    .X(_11833_));
 sky130_fd_sc_hd__and2_1 _26914_ (.A(_11833_),
    .B(_11823_),
    .X(_11834_));
 sky130_fd_sc_hd__a31o_1 _26915_ (.A1(_11831_),
    .A2(\datamem.data_ram[32][5] ),
    .A3(_11821_),
    .B1(_11834_),
    .X(_03370_));
 sky130_fd_sc_hd__buf_2 _26916_ (.A(_10072_),
    .X(_11835_));
 sky130_fd_sc_hd__and2_1 _26917_ (.A(_11835_),
    .B(_11823_),
    .X(_11836_));
 sky130_fd_sc_hd__a31o_1 _26918_ (.A1(_11831_),
    .A2(\datamem.data_ram[32][6] ),
    .A3(_11821_),
    .B1(_11836_),
    .X(_03371_));
 sky130_fd_sc_hd__clkbuf_4 _26919_ (.A(_10075_),
    .X(_11837_));
 sky130_fd_sc_hd__and2_1 _26920_ (.A(_11837_),
    .B(_11823_),
    .X(_11838_));
 sky130_fd_sc_hd__a31o_1 _26921_ (.A1(_11831_),
    .A2(\datamem.data_ram[32][7] ),
    .A3(_11821_),
    .B1(_11838_),
    .X(_03372_));
 sky130_fd_sc_hd__buf_2 _26922_ (.A(_10043_),
    .X(_11839_));
 sky130_fd_sc_hd__or3_1 _26923_ (.A(_07791_),
    .B(_10402_),
    .C(_11839_),
    .X(_11840_));
 sky130_fd_sc_hd__buf_2 _26924_ (.A(_11840_),
    .X(_11841_));
 sky130_fd_sc_hd__and3_2 _26925_ (.A(_10325_),
    .B(_08059_),
    .C(_11609_),
    .X(_11842_));
 sky130_fd_sc_hd__and2_1 _26926_ (.A(_11822_),
    .B(_11842_),
    .X(_11843_));
 sky130_fd_sc_hd__a31o_1 _26927_ (.A1(_11831_),
    .A2(\datamem.data_ram[55][0] ),
    .A3(_11841_),
    .B1(_11843_),
    .X(_03373_));
 sky130_fd_sc_hd__and2_1 _26928_ (.A(_11825_),
    .B(_11842_),
    .X(_11844_));
 sky130_fd_sc_hd__a31o_1 _26929_ (.A1(_11831_),
    .A2(\datamem.data_ram[55][1] ),
    .A3(_11841_),
    .B1(_11844_),
    .X(_03374_));
 sky130_fd_sc_hd__and2_1 _26930_ (.A(_11827_),
    .B(_11842_),
    .X(_11845_));
 sky130_fd_sc_hd__a31o_1 _26931_ (.A1(_11831_),
    .A2(\datamem.data_ram[55][2] ),
    .A3(_11841_),
    .B1(_11845_),
    .X(_03375_));
 sky130_fd_sc_hd__and2_1 _26932_ (.A(_11829_),
    .B(_11842_),
    .X(_11846_));
 sky130_fd_sc_hd__a31o_1 _26933_ (.A1(_11831_),
    .A2(\datamem.data_ram[55][3] ),
    .A3(_11841_),
    .B1(_11846_),
    .X(_03376_));
 sky130_fd_sc_hd__and2_1 _26934_ (.A(_11803_),
    .B(_11842_),
    .X(_11847_));
 sky130_fd_sc_hd__a31o_1 _26935_ (.A1(_11831_),
    .A2(\datamem.data_ram[55][4] ),
    .A3(_11841_),
    .B1(_11847_),
    .X(_03377_));
 sky130_fd_sc_hd__and2_1 _26936_ (.A(_11833_),
    .B(_11842_),
    .X(_11848_));
 sky130_fd_sc_hd__a31o_1 _26937_ (.A1(_11831_),
    .A2(\datamem.data_ram[55][5] ),
    .A3(_11841_),
    .B1(_11848_),
    .X(_03378_));
 sky130_fd_sc_hd__clkbuf_4 _26938_ (.A(_11752_),
    .X(_11849_));
 sky130_fd_sc_hd__and2_1 _26939_ (.A(_11835_),
    .B(_11842_),
    .X(_11850_));
 sky130_fd_sc_hd__a31o_1 _26940_ (.A1(_11849_),
    .A2(\datamem.data_ram[55][6] ),
    .A3(_11841_),
    .B1(_11850_),
    .X(_03379_));
 sky130_fd_sc_hd__and2_1 _26941_ (.A(_11837_),
    .B(_11842_),
    .X(_11851_));
 sky130_fd_sc_hd__a31o_1 _26942_ (.A1(_11849_),
    .A2(\datamem.data_ram[55][7] ),
    .A3(_11841_),
    .B1(_11851_),
    .X(_03380_));
 sky130_fd_sc_hd__or3_1 _26943_ (.A(_07182_),
    .B(_11109_),
    .C(_11839_),
    .X(_11852_));
 sky130_fd_sc_hd__buf_2 _26944_ (.A(_11852_),
    .X(_11853_));
 sky130_fd_sc_hd__and3_1 _26945_ (.A(_09351_),
    .B(_11112_),
    .C(_11609_),
    .X(_11854_));
 sky130_fd_sc_hd__and2_1 _26946_ (.A(_11822_),
    .B(_11854_),
    .X(_11855_));
 sky130_fd_sc_hd__a31o_1 _26947_ (.A1(_11849_),
    .A2(\datamem.data_ram[28][0] ),
    .A3(_11853_),
    .B1(_11855_),
    .X(_03381_));
 sky130_fd_sc_hd__and2_1 _26948_ (.A(_11825_),
    .B(_11854_),
    .X(_11856_));
 sky130_fd_sc_hd__a31o_1 _26949_ (.A1(_11849_),
    .A2(\datamem.data_ram[28][1] ),
    .A3(_11853_),
    .B1(_11856_),
    .X(_03382_));
 sky130_fd_sc_hd__and2_1 _26950_ (.A(_11827_),
    .B(_11854_),
    .X(_11857_));
 sky130_fd_sc_hd__a31o_1 _26951_ (.A1(_11849_),
    .A2(\datamem.data_ram[28][2] ),
    .A3(_11853_),
    .B1(_11857_),
    .X(_03383_));
 sky130_fd_sc_hd__and2_1 _26952_ (.A(_11829_),
    .B(_11854_),
    .X(_11858_));
 sky130_fd_sc_hd__a31o_1 _26953_ (.A1(_11849_),
    .A2(\datamem.data_ram[28][3] ),
    .A3(_11853_),
    .B1(_11858_),
    .X(_03384_));
 sky130_fd_sc_hd__and2_1 _26954_ (.A(_11803_),
    .B(_11854_),
    .X(_11859_));
 sky130_fd_sc_hd__a31o_1 _26955_ (.A1(_11849_),
    .A2(\datamem.data_ram[28][4] ),
    .A3(_11853_),
    .B1(_11859_),
    .X(_03385_));
 sky130_fd_sc_hd__and2_1 _26956_ (.A(_11833_),
    .B(_11854_),
    .X(_11860_));
 sky130_fd_sc_hd__a31o_1 _26957_ (.A1(_11849_),
    .A2(\datamem.data_ram[28][5] ),
    .A3(_11853_),
    .B1(_11860_),
    .X(_03386_));
 sky130_fd_sc_hd__and2_1 _26958_ (.A(_11835_),
    .B(_11854_),
    .X(_11861_));
 sky130_fd_sc_hd__a31o_1 _26959_ (.A1(_11849_),
    .A2(\datamem.data_ram[28][6] ),
    .A3(_11853_),
    .B1(_11861_),
    .X(_03387_));
 sky130_fd_sc_hd__and2_1 _26960_ (.A(_11837_),
    .B(_11854_),
    .X(_11862_));
 sky130_fd_sc_hd__a31o_1 _26961_ (.A1(_11849_),
    .A2(\datamem.data_ram[28][7] ),
    .A3(_11853_),
    .B1(_11862_),
    .X(_03388_));
 sky130_fd_sc_hd__clkbuf_4 _26962_ (.A(_11752_),
    .X(_11863_));
 sky130_fd_sc_hd__or2_1 _26963_ (.A(_10402_),
    .B(_10947_),
    .X(_11864_));
 sky130_fd_sc_hd__clkbuf_2 _26964_ (.A(_11864_),
    .X(_11865_));
 sky130_fd_sc_hd__nor2_1 _26965_ (.A(_10402_),
    .B(_10947_),
    .Y(_11866_));
 sky130_fd_sc_hd__and2_1 _26966_ (.A(_11822_),
    .B(_11866_),
    .X(_11867_));
 sky130_fd_sc_hd__a31o_1 _26967_ (.A1(_11863_),
    .A2(\datamem.data_ram[54][0] ),
    .A3(_11865_),
    .B1(_11867_),
    .X(_03389_));
 sky130_fd_sc_hd__and2_1 _26968_ (.A(_11825_),
    .B(_11866_),
    .X(_11868_));
 sky130_fd_sc_hd__a31o_1 _26969_ (.A1(_11863_),
    .A2(\datamem.data_ram[54][1] ),
    .A3(_11865_),
    .B1(_11868_),
    .X(_03390_));
 sky130_fd_sc_hd__and2_1 _26970_ (.A(_11827_),
    .B(_11866_),
    .X(_11869_));
 sky130_fd_sc_hd__a31o_1 _26971_ (.A1(_11863_),
    .A2(\datamem.data_ram[54][2] ),
    .A3(_11865_),
    .B1(_11869_),
    .X(_03391_));
 sky130_fd_sc_hd__and2_1 _26972_ (.A(_11829_),
    .B(_11866_),
    .X(_11870_));
 sky130_fd_sc_hd__a31o_1 _26973_ (.A1(_11863_),
    .A2(\datamem.data_ram[54][3] ),
    .A3(_11865_),
    .B1(_11870_),
    .X(_03392_));
 sky130_fd_sc_hd__and2_1 _26974_ (.A(_11803_),
    .B(_11866_),
    .X(_11871_));
 sky130_fd_sc_hd__a31o_1 _26975_ (.A1(_11863_),
    .A2(\datamem.data_ram[54][4] ),
    .A3(_11865_),
    .B1(_11871_),
    .X(_03393_));
 sky130_fd_sc_hd__and2_1 _26976_ (.A(_11833_),
    .B(_11866_),
    .X(_11872_));
 sky130_fd_sc_hd__a31o_1 _26977_ (.A1(_11863_),
    .A2(\datamem.data_ram[54][5] ),
    .A3(_11865_),
    .B1(_11872_),
    .X(_03394_));
 sky130_fd_sc_hd__and2_1 _26978_ (.A(_11835_),
    .B(_11866_),
    .X(_11873_));
 sky130_fd_sc_hd__a31o_1 _26979_ (.A1(_11863_),
    .A2(\datamem.data_ram[54][6] ),
    .A3(_11865_),
    .B1(_11873_),
    .X(_03395_));
 sky130_fd_sc_hd__and2_1 _26980_ (.A(_11837_),
    .B(_11866_),
    .X(_11874_));
 sky130_fd_sc_hd__a31o_1 _26981_ (.A1(_11863_),
    .A2(\datamem.data_ram[54][7] ),
    .A3(_11865_),
    .B1(_11874_),
    .X(_03396_));
 sky130_fd_sc_hd__a21oi_4 _26982_ (.A1(_10113_),
    .A2(_10337_),
    .B1(_11713_),
    .Y(_11875_));
 sky130_fd_sc_hd__mux2_1 _26983_ (.A0(_10751_),
    .A1(\datamem.data_ram[53][16] ),
    .S(_11875_),
    .X(_11876_));
 sky130_fd_sc_hd__clkbuf_1 _26984_ (.A(_11876_),
    .X(_03397_));
 sky130_fd_sc_hd__mux2_1 _26985_ (.A0(_10754_),
    .A1(\datamem.data_ram[53][17] ),
    .S(_11875_),
    .X(_11877_));
 sky130_fd_sc_hd__clkbuf_1 _26986_ (.A(_11877_),
    .X(_03398_));
 sky130_fd_sc_hd__mux2_1 _26987_ (.A0(_10756_),
    .A1(\datamem.data_ram[53][18] ),
    .S(_11875_),
    .X(_11878_));
 sky130_fd_sc_hd__clkbuf_1 _26988_ (.A(_11878_),
    .X(_03399_));
 sky130_fd_sc_hd__mux2_1 _26989_ (.A0(_10758_),
    .A1(\datamem.data_ram[53][19] ),
    .S(_11875_),
    .X(_11879_));
 sky130_fd_sc_hd__clkbuf_1 _26990_ (.A(_11879_),
    .X(_03400_));
 sky130_fd_sc_hd__mux2_1 _26991_ (.A0(_10760_),
    .A1(\datamem.data_ram[53][20] ),
    .S(_11875_),
    .X(_11880_));
 sky130_fd_sc_hd__clkbuf_1 _26992_ (.A(_11880_),
    .X(_03401_));
 sky130_fd_sc_hd__mux2_1 _26993_ (.A0(_10762_),
    .A1(\datamem.data_ram[53][21] ),
    .S(_11875_),
    .X(_11881_));
 sky130_fd_sc_hd__clkbuf_1 _26994_ (.A(_11881_),
    .X(_03402_));
 sky130_fd_sc_hd__mux2_1 _26995_ (.A0(_10764_),
    .A1(\datamem.data_ram[53][22] ),
    .S(_11875_),
    .X(_11882_));
 sky130_fd_sc_hd__clkbuf_1 _26996_ (.A(_11882_),
    .X(_03403_));
 sky130_fd_sc_hd__mux2_1 _26997_ (.A0(_10766_),
    .A1(\datamem.data_ram[53][23] ),
    .S(_11875_),
    .X(_11883_));
 sky130_fd_sc_hd__clkbuf_1 _26998_ (.A(_11883_),
    .X(_03404_));
 sky130_fd_sc_hd__or3_1 _26999_ (.A(_07019_),
    .B(_10918_),
    .C(_10897_),
    .X(_11884_));
 sky130_fd_sc_hd__clkbuf_2 _27000_ (.A(_11884_),
    .X(_11885_));
 sky130_fd_sc_hd__and3_1 _27001_ (.A(_09299_),
    .B(_10921_),
    .C(_10922_),
    .X(_11886_));
 sky130_fd_sc_hd__and2_1 _27002_ (.A(_11822_),
    .B(_11886_),
    .X(_11887_));
 sky130_fd_sc_hd__a31o_1 _27003_ (.A1(_11863_),
    .A2(\datamem.data_ram[37][0] ),
    .A3(_11885_),
    .B1(_11887_),
    .X(_03405_));
 sky130_fd_sc_hd__and2_1 _27004_ (.A(_11825_),
    .B(_11886_),
    .X(_11888_));
 sky130_fd_sc_hd__a31o_1 _27005_ (.A1(_11863_),
    .A2(\datamem.data_ram[37][1] ),
    .A3(_11885_),
    .B1(_11888_),
    .X(_03406_));
 sky130_fd_sc_hd__clkbuf_4 _27006_ (.A(_11752_),
    .X(_11889_));
 sky130_fd_sc_hd__and2_1 _27007_ (.A(_11827_),
    .B(_11886_),
    .X(_11890_));
 sky130_fd_sc_hd__a31o_1 _27008_ (.A1(_11889_),
    .A2(\datamem.data_ram[37][2] ),
    .A3(_11885_),
    .B1(_11890_),
    .X(_03407_));
 sky130_fd_sc_hd__and2_1 _27009_ (.A(_11829_),
    .B(_11886_),
    .X(_11891_));
 sky130_fd_sc_hd__a31o_1 _27010_ (.A1(_11889_),
    .A2(\datamem.data_ram[37][3] ),
    .A3(_11885_),
    .B1(_11891_),
    .X(_03408_));
 sky130_fd_sc_hd__and2_1 _27011_ (.A(_11803_),
    .B(_11886_),
    .X(_11892_));
 sky130_fd_sc_hd__a31o_1 _27012_ (.A1(_11889_),
    .A2(\datamem.data_ram[37][4] ),
    .A3(_11885_),
    .B1(_11892_),
    .X(_03409_));
 sky130_fd_sc_hd__and2_1 _27013_ (.A(_11833_),
    .B(_11886_),
    .X(_11893_));
 sky130_fd_sc_hd__a31o_1 _27014_ (.A1(_11889_),
    .A2(\datamem.data_ram[37][5] ),
    .A3(_11885_),
    .B1(_11893_),
    .X(_03410_));
 sky130_fd_sc_hd__and2_1 _27015_ (.A(_11835_),
    .B(_11886_),
    .X(_11894_));
 sky130_fd_sc_hd__a31o_1 _27016_ (.A1(_11889_),
    .A2(\datamem.data_ram[37][6] ),
    .A3(_11885_),
    .B1(_11894_),
    .X(_03411_));
 sky130_fd_sc_hd__and2_1 _27017_ (.A(_11837_),
    .B(_11886_),
    .X(_11895_));
 sky130_fd_sc_hd__a31o_1 _27018_ (.A1(_11889_),
    .A2(\datamem.data_ram[37][7] ),
    .A3(_11885_),
    .B1(_11895_),
    .X(_03412_));
 sky130_fd_sc_hd__or3_1 _27019_ (.A(_07791_),
    .B(_11109_),
    .C(_11839_),
    .X(_11896_));
 sky130_fd_sc_hd__clkbuf_2 _27020_ (.A(_11896_),
    .X(_11897_));
 sky130_fd_sc_hd__buf_2 _27021_ (.A(_10051_),
    .X(_11898_));
 sky130_fd_sc_hd__and3_1 _27022_ (.A(_10325_),
    .B(_11112_),
    .C(_11898_),
    .X(_11899_));
 sky130_fd_sc_hd__and2_1 _27023_ (.A(_11822_),
    .B(_11899_),
    .X(_11900_));
 sky130_fd_sc_hd__a31o_1 _27024_ (.A1(_11889_),
    .A2(\datamem.data_ram[31][0] ),
    .A3(_11897_),
    .B1(_11900_),
    .X(_03413_));
 sky130_fd_sc_hd__and2_1 _27025_ (.A(_11825_),
    .B(_11899_),
    .X(_11901_));
 sky130_fd_sc_hd__a31o_1 _27026_ (.A1(_11889_),
    .A2(\datamem.data_ram[31][1] ),
    .A3(_11897_),
    .B1(_11901_),
    .X(_03414_));
 sky130_fd_sc_hd__and2_1 _27027_ (.A(_11827_),
    .B(_11899_),
    .X(_11902_));
 sky130_fd_sc_hd__a31o_1 _27028_ (.A1(_11889_),
    .A2(\datamem.data_ram[31][2] ),
    .A3(_11897_),
    .B1(_11902_),
    .X(_03415_));
 sky130_fd_sc_hd__and2_1 _27029_ (.A(_11829_),
    .B(_11899_),
    .X(_11903_));
 sky130_fd_sc_hd__a31o_1 _27030_ (.A1(_11889_),
    .A2(\datamem.data_ram[31][3] ),
    .A3(_11897_),
    .B1(_11903_),
    .X(_03416_));
 sky130_fd_sc_hd__clkbuf_4 _27031_ (.A(_11752_),
    .X(_11904_));
 sky130_fd_sc_hd__and2_1 _27032_ (.A(_11803_),
    .B(_11899_),
    .X(_11905_));
 sky130_fd_sc_hd__a31o_1 _27033_ (.A1(_11904_),
    .A2(\datamem.data_ram[31][4] ),
    .A3(_11897_),
    .B1(_11905_),
    .X(_03417_));
 sky130_fd_sc_hd__and2_1 _27034_ (.A(_11833_),
    .B(_11899_),
    .X(_11906_));
 sky130_fd_sc_hd__a31o_1 _27035_ (.A1(_11904_),
    .A2(\datamem.data_ram[31][5] ),
    .A3(_11897_),
    .B1(_11906_),
    .X(_03418_));
 sky130_fd_sc_hd__and2_1 _27036_ (.A(_11835_),
    .B(_11899_),
    .X(_11907_));
 sky130_fd_sc_hd__a31o_1 _27037_ (.A1(_11904_),
    .A2(\datamem.data_ram[31][6] ),
    .A3(_11897_),
    .B1(_11907_),
    .X(_03419_));
 sky130_fd_sc_hd__and2_1 _27038_ (.A(_11837_),
    .B(_11899_),
    .X(_11908_));
 sky130_fd_sc_hd__a31o_1 _27039_ (.A1(_11904_),
    .A2(\datamem.data_ram[31][7] ),
    .A3(_11897_),
    .B1(_11908_),
    .X(_03420_));
 sky130_fd_sc_hd__or2_1 _27040_ (.A(_10402_),
    .B(_11039_),
    .X(_11909_));
 sky130_fd_sc_hd__clkbuf_2 _27041_ (.A(_11909_),
    .X(_11910_));
 sky130_fd_sc_hd__nor2_1 _27042_ (.A(_10402_),
    .B(_11039_),
    .Y(_11911_));
 sky130_fd_sc_hd__and2_1 _27043_ (.A(_11822_),
    .B(_11911_),
    .X(_11912_));
 sky130_fd_sc_hd__a31o_1 _27044_ (.A1(_11904_),
    .A2(\datamem.data_ram[52][0] ),
    .A3(_11910_),
    .B1(_11912_),
    .X(_03421_));
 sky130_fd_sc_hd__and2_1 _27045_ (.A(_11825_),
    .B(_11911_),
    .X(_11913_));
 sky130_fd_sc_hd__a31o_1 _27046_ (.A1(_11904_),
    .A2(\datamem.data_ram[52][1] ),
    .A3(_11910_),
    .B1(_11913_),
    .X(_03422_));
 sky130_fd_sc_hd__and2_1 _27047_ (.A(_11827_),
    .B(_11911_),
    .X(_11914_));
 sky130_fd_sc_hd__a31o_1 _27048_ (.A1(_11904_),
    .A2(\datamem.data_ram[52][2] ),
    .A3(_11910_),
    .B1(_11914_),
    .X(_03423_));
 sky130_fd_sc_hd__and2_1 _27049_ (.A(_11829_),
    .B(_11911_),
    .X(_11915_));
 sky130_fd_sc_hd__a31o_1 _27050_ (.A1(_11904_),
    .A2(\datamem.data_ram[52][3] ),
    .A3(_11910_),
    .B1(_11915_),
    .X(_03424_));
 sky130_fd_sc_hd__and2_1 _27051_ (.A(_11803_),
    .B(_11911_),
    .X(_11916_));
 sky130_fd_sc_hd__a31o_1 _27052_ (.A1(_11904_),
    .A2(\datamem.data_ram[52][4] ),
    .A3(_11910_),
    .B1(_11916_),
    .X(_03425_));
 sky130_fd_sc_hd__and2_1 _27053_ (.A(_11833_),
    .B(_11911_),
    .X(_11917_));
 sky130_fd_sc_hd__a31o_1 _27054_ (.A1(_11904_),
    .A2(\datamem.data_ram[52][5] ),
    .A3(_11910_),
    .B1(_11917_),
    .X(_03426_));
 sky130_fd_sc_hd__buf_2 _27055_ (.A(_06587_),
    .X(_11918_));
 sky130_fd_sc_hd__clkbuf_4 _27056_ (.A(_11918_),
    .X(_11919_));
 sky130_fd_sc_hd__and2_1 _27057_ (.A(_11835_),
    .B(_11911_),
    .X(_11920_));
 sky130_fd_sc_hd__a31o_1 _27058_ (.A1(_11919_),
    .A2(\datamem.data_ram[52][6] ),
    .A3(_11910_),
    .B1(_11920_),
    .X(_03427_));
 sky130_fd_sc_hd__and2_1 _27059_ (.A(_11837_),
    .B(_11911_),
    .X(_11921_));
 sky130_fd_sc_hd__a31o_1 _27060_ (.A1(_11919_),
    .A2(\datamem.data_ram[52][7] ),
    .A3(_11910_),
    .B1(_11921_),
    .X(_03428_));
 sky130_fd_sc_hd__or3_1 _27061_ (.A(_07077_),
    .B(_11109_),
    .C(_11839_),
    .X(_11922_));
 sky130_fd_sc_hd__clkbuf_2 _27062_ (.A(_11922_),
    .X(_11923_));
 sky130_fd_sc_hd__and3_1 _27063_ (.A(_10142_),
    .B(_11112_),
    .C(_11898_),
    .X(_11924_));
 sky130_fd_sc_hd__and2_1 _27064_ (.A(_11822_),
    .B(_11924_),
    .X(_11925_));
 sky130_fd_sc_hd__a31o_1 _27065_ (.A1(_11919_),
    .A2(\datamem.data_ram[27][0] ),
    .A3(_11923_),
    .B1(_11925_),
    .X(_03429_));
 sky130_fd_sc_hd__and2_1 _27066_ (.A(_11825_),
    .B(_11924_),
    .X(_11926_));
 sky130_fd_sc_hd__a31o_1 _27067_ (.A1(_11919_),
    .A2(\datamem.data_ram[27][1] ),
    .A3(_11923_),
    .B1(_11926_),
    .X(_03430_));
 sky130_fd_sc_hd__and2_1 _27068_ (.A(_11827_),
    .B(_11924_),
    .X(_11927_));
 sky130_fd_sc_hd__a31o_1 _27069_ (.A1(_11919_),
    .A2(\datamem.data_ram[27][2] ),
    .A3(_11923_),
    .B1(_11927_),
    .X(_03431_));
 sky130_fd_sc_hd__and2_1 _27070_ (.A(_11829_),
    .B(_11924_),
    .X(_11928_));
 sky130_fd_sc_hd__a31o_1 _27071_ (.A1(_11919_),
    .A2(\datamem.data_ram[27][3] ),
    .A3(_11923_),
    .B1(_11928_),
    .X(_03432_));
 sky130_fd_sc_hd__and2_1 _27072_ (.A(_11803_),
    .B(_11924_),
    .X(_11929_));
 sky130_fd_sc_hd__a31o_1 _27073_ (.A1(_11919_),
    .A2(\datamem.data_ram[27][4] ),
    .A3(_11923_),
    .B1(_11929_),
    .X(_03433_));
 sky130_fd_sc_hd__and2_1 _27074_ (.A(_11833_),
    .B(_11924_),
    .X(_11930_));
 sky130_fd_sc_hd__a31o_1 _27075_ (.A1(_11919_),
    .A2(\datamem.data_ram[27][5] ),
    .A3(_11923_),
    .B1(_11930_),
    .X(_03434_));
 sky130_fd_sc_hd__and2_1 _27076_ (.A(_11835_),
    .B(_11924_),
    .X(_11931_));
 sky130_fd_sc_hd__a31o_1 _27077_ (.A1(_11919_),
    .A2(\datamem.data_ram[27][6] ),
    .A3(_11923_),
    .B1(_11931_),
    .X(_03435_));
 sky130_fd_sc_hd__and2_1 _27078_ (.A(_11837_),
    .B(_11924_),
    .X(_11932_));
 sky130_fd_sc_hd__a31o_1 _27079_ (.A1(_11919_),
    .A2(\datamem.data_ram[27][7] ),
    .A3(_11923_),
    .B1(_11932_),
    .X(_03436_));
 sky130_fd_sc_hd__nor2_1 _27080_ (.A(_11153_),
    .B(_11146_),
    .Y(_11933_));
 sky130_fd_sc_hd__mux2_1 _27081_ (.A0(\rvcpu.ALUResultE[0] ),
    .A1(_06354_),
    .S(_11598_),
    .X(_11934_));
 sky130_fd_sc_hd__or2_1 _27082_ (.A(_11526_),
    .B(_11934_),
    .X(_11935_));
 sky130_fd_sc_hd__o211a_1 _27083_ (.A1(\rvcpu.dp.pcreg.q[0] ),
    .A2(_11933_),
    .B1(_11935_),
    .C1(_10041_),
    .X(_03437_));
 sky130_fd_sc_hd__mux2_1 _27084_ (.A0(\rvcpu.ALUResultE[1] ),
    .A1(_06358_),
    .S(_11598_),
    .X(_11936_));
 sky130_fd_sc_hd__or2_1 _27085_ (.A(_11526_),
    .B(_11936_),
    .X(_11937_));
 sky130_fd_sc_hd__o211a_1 _27086_ (.A1(\rvcpu.dp.pcreg.q[1] ),
    .A2(_11933_),
    .B1(_11937_),
    .C1(_10041_),
    .X(_03438_));
 sky130_fd_sc_hd__buf_2 _27087_ (.A(_11918_),
    .X(_11938_));
 sky130_fd_sc_hd__or2_1 _27088_ (.A(_10402_),
    .B(_11075_),
    .X(_11939_));
 sky130_fd_sc_hd__clkbuf_2 _27089_ (.A(_11939_),
    .X(_11940_));
 sky130_fd_sc_hd__nor2_1 _27090_ (.A(_10402_),
    .B(_11075_),
    .Y(_11941_));
 sky130_fd_sc_hd__and2_1 _27091_ (.A(_11822_),
    .B(_11941_),
    .X(_11942_));
 sky130_fd_sc_hd__a31o_1 _27092_ (.A1(_11938_),
    .A2(\datamem.data_ram[51][0] ),
    .A3(_11940_),
    .B1(_11942_),
    .X(_03439_));
 sky130_fd_sc_hd__and2_1 _27093_ (.A(_11825_),
    .B(_11941_),
    .X(_11943_));
 sky130_fd_sc_hd__a31o_1 _27094_ (.A1(_11938_),
    .A2(\datamem.data_ram[51][1] ),
    .A3(_11940_),
    .B1(_11943_),
    .X(_03440_));
 sky130_fd_sc_hd__and2_1 _27095_ (.A(_11827_),
    .B(_11941_),
    .X(_11944_));
 sky130_fd_sc_hd__a31o_1 _27096_ (.A1(_11938_),
    .A2(\datamem.data_ram[51][2] ),
    .A3(_11940_),
    .B1(_11944_),
    .X(_03441_));
 sky130_fd_sc_hd__and2_1 _27097_ (.A(_11829_),
    .B(_11941_),
    .X(_11945_));
 sky130_fd_sc_hd__a31o_1 _27098_ (.A1(_11938_),
    .A2(\datamem.data_ram[51][3] ),
    .A3(_11940_),
    .B1(_11945_),
    .X(_03442_));
 sky130_fd_sc_hd__clkbuf_4 _27099_ (.A(_10066_),
    .X(_11946_));
 sky130_fd_sc_hd__and2_1 _27100_ (.A(_11946_),
    .B(_11941_),
    .X(_11947_));
 sky130_fd_sc_hd__a31o_1 _27101_ (.A1(_11938_),
    .A2(\datamem.data_ram[51][4] ),
    .A3(_11940_),
    .B1(_11947_),
    .X(_03443_));
 sky130_fd_sc_hd__and2_1 _27102_ (.A(_11833_),
    .B(_11941_),
    .X(_11948_));
 sky130_fd_sc_hd__a31o_1 _27103_ (.A1(_11938_),
    .A2(\datamem.data_ram[51][5] ),
    .A3(_11940_),
    .B1(_11948_),
    .X(_03444_));
 sky130_fd_sc_hd__and2_1 _27104_ (.A(_11835_),
    .B(_11941_),
    .X(_11949_));
 sky130_fd_sc_hd__a31o_1 _27105_ (.A1(_11938_),
    .A2(\datamem.data_ram[51][6] ),
    .A3(_11940_),
    .B1(_11949_),
    .X(_03445_));
 sky130_fd_sc_hd__and2_1 _27106_ (.A(_11837_),
    .B(_11941_),
    .X(_11950_));
 sky130_fd_sc_hd__a31o_1 _27107_ (.A1(_11938_),
    .A2(\datamem.data_ram[51][7] ),
    .A3(_11940_),
    .B1(_11950_),
    .X(_03446_));
 sky130_fd_sc_hd__or2_1 _27108_ (.A(_11109_),
    .B(_10778_),
    .X(_11951_));
 sky130_fd_sc_hd__clkbuf_2 _27109_ (.A(_11951_),
    .X(_11952_));
 sky130_fd_sc_hd__nor2_1 _27110_ (.A(_11109_),
    .B(_10778_),
    .Y(_11953_));
 sky130_fd_sc_hd__and2_1 _27111_ (.A(_11822_),
    .B(_11953_),
    .X(_11954_));
 sky130_fd_sc_hd__a31o_1 _27112_ (.A1(_11938_),
    .A2(\datamem.data_ram[26][0] ),
    .A3(_11952_),
    .B1(_11954_),
    .X(_03447_));
 sky130_fd_sc_hd__and2_1 _27113_ (.A(_11825_),
    .B(_11953_),
    .X(_11955_));
 sky130_fd_sc_hd__a31o_1 _27114_ (.A1(_11938_),
    .A2(\datamem.data_ram[26][1] ),
    .A3(_11952_),
    .B1(_11955_),
    .X(_03448_));
 sky130_fd_sc_hd__buf_2 _27115_ (.A(_11918_),
    .X(_11956_));
 sky130_fd_sc_hd__and2_1 _27116_ (.A(_11827_),
    .B(_11953_),
    .X(_11957_));
 sky130_fd_sc_hd__a31o_1 _27117_ (.A1(_11956_),
    .A2(\datamem.data_ram[26][2] ),
    .A3(_11952_),
    .B1(_11957_),
    .X(_03449_));
 sky130_fd_sc_hd__and2_1 _27118_ (.A(_11829_),
    .B(_11953_),
    .X(_11958_));
 sky130_fd_sc_hd__a31o_1 _27119_ (.A1(_11956_),
    .A2(\datamem.data_ram[26][3] ),
    .A3(_11952_),
    .B1(_11958_),
    .X(_03450_));
 sky130_fd_sc_hd__and2_1 _27120_ (.A(_11946_),
    .B(_11953_),
    .X(_11959_));
 sky130_fd_sc_hd__a31o_1 _27121_ (.A1(_11956_),
    .A2(\datamem.data_ram[26][4] ),
    .A3(_11952_),
    .B1(_11959_),
    .X(_03451_));
 sky130_fd_sc_hd__and2_1 _27122_ (.A(_11833_),
    .B(_11953_),
    .X(_11960_));
 sky130_fd_sc_hd__a31o_1 _27123_ (.A1(_11956_),
    .A2(\datamem.data_ram[26][5] ),
    .A3(_11952_),
    .B1(_11960_),
    .X(_03452_));
 sky130_fd_sc_hd__and2_1 _27124_ (.A(_11835_),
    .B(_11953_),
    .X(_11961_));
 sky130_fd_sc_hd__a31o_1 _27125_ (.A1(_11956_),
    .A2(\datamem.data_ram[26][6] ),
    .A3(_11952_),
    .B1(_11961_),
    .X(_03453_));
 sky130_fd_sc_hd__and2_1 _27126_ (.A(_11837_),
    .B(_11953_),
    .X(_11962_));
 sky130_fd_sc_hd__a31o_1 _27127_ (.A1(_11956_),
    .A2(\datamem.data_ram[26][7] ),
    .A3(_11952_),
    .B1(_11962_),
    .X(_03454_));
 sky130_fd_sc_hd__or3_1 _27128_ (.A(_07203_),
    .B(_10326_),
    .C(_11839_),
    .X(_11963_));
 sky130_fd_sc_hd__buf_2 _27129_ (.A(_11963_),
    .X(_11964_));
 sky130_fd_sc_hd__buf_2 _27130_ (.A(_10047_),
    .X(_11965_));
 sky130_fd_sc_hd__and3_1 _27131_ (.A(_10209_),
    .B(_08059_),
    .C(_11898_),
    .X(_11966_));
 sky130_fd_sc_hd__and2_1 _27132_ (.A(_11965_),
    .B(_11966_),
    .X(_11967_));
 sky130_fd_sc_hd__a31o_1 _27133_ (.A1(_11956_),
    .A2(\datamem.data_ram[50][0] ),
    .A3(_11964_),
    .B1(_11967_),
    .X(_03455_));
 sky130_fd_sc_hd__clkbuf_4 _27134_ (.A(_10057_),
    .X(_11968_));
 sky130_fd_sc_hd__and2_1 _27135_ (.A(_11968_),
    .B(_11966_),
    .X(_11969_));
 sky130_fd_sc_hd__a31o_1 _27136_ (.A1(_11956_),
    .A2(\datamem.data_ram[50][1] ),
    .A3(_11964_),
    .B1(_11969_),
    .X(_03456_));
 sky130_fd_sc_hd__clkbuf_4 _27137_ (.A(_10060_),
    .X(_11970_));
 sky130_fd_sc_hd__and2_1 _27138_ (.A(_11970_),
    .B(_11966_),
    .X(_11971_));
 sky130_fd_sc_hd__a31o_1 _27139_ (.A1(_11956_),
    .A2(\datamem.data_ram[50][2] ),
    .A3(_11964_),
    .B1(_11971_),
    .X(_03457_));
 sky130_fd_sc_hd__clkbuf_4 _27140_ (.A(_10063_),
    .X(_11972_));
 sky130_fd_sc_hd__and2_1 _27141_ (.A(_11972_),
    .B(_11966_),
    .X(_11973_));
 sky130_fd_sc_hd__a31o_1 _27142_ (.A1(_11956_),
    .A2(\datamem.data_ram[50][3] ),
    .A3(_11964_),
    .B1(_11973_),
    .X(_03458_));
 sky130_fd_sc_hd__buf_2 _27143_ (.A(_11918_),
    .X(_11974_));
 sky130_fd_sc_hd__and2_1 _27144_ (.A(_11946_),
    .B(_11966_),
    .X(_11975_));
 sky130_fd_sc_hd__a31o_1 _27145_ (.A1(_11974_),
    .A2(\datamem.data_ram[50][4] ),
    .A3(_11964_),
    .B1(_11975_),
    .X(_03459_));
 sky130_fd_sc_hd__buf_2 _27146_ (.A(_10069_),
    .X(_11976_));
 sky130_fd_sc_hd__and2_1 _27147_ (.A(_11976_),
    .B(_11966_),
    .X(_11977_));
 sky130_fd_sc_hd__a31o_1 _27148_ (.A1(_11974_),
    .A2(\datamem.data_ram[50][5] ),
    .A3(_11964_),
    .B1(_11977_),
    .X(_03460_));
 sky130_fd_sc_hd__clkbuf_4 _27149_ (.A(_10072_),
    .X(_11978_));
 sky130_fd_sc_hd__and2_1 _27150_ (.A(_11978_),
    .B(_11966_),
    .X(_11979_));
 sky130_fd_sc_hd__a31o_1 _27151_ (.A1(_11974_),
    .A2(\datamem.data_ram[50][6] ),
    .A3(_11964_),
    .B1(_11979_),
    .X(_03461_));
 sky130_fd_sc_hd__clkbuf_4 _27152_ (.A(_10075_),
    .X(_11980_));
 sky130_fd_sc_hd__and2_1 _27153_ (.A(_11980_),
    .B(_11966_),
    .X(_11981_));
 sky130_fd_sc_hd__a31o_1 _27154_ (.A1(_11974_),
    .A2(\datamem.data_ram[50][7] ),
    .A3(_11964_),
    .B1(_11981_),
    .X(_03462_));
 sky130_fd_sc_hd__or3_1 _27155_ (.A(_07808_),
    .B(_10326_),
    .C(_11839_),
    .X(_11982_));
 sky130_fd_sc_hd__buf_2 _27156_ (.A(_11982_),
    .X(_11983_));
 sky130_fd_sc_hd__and3_1 _27157_ (.A(_10268_),
    .B(_08059_),
    .C(_11898_),
    .X(_11984_));
 sky130_fd_sc_hd__and2_1 _27158_ (.A(_11965_),
    .B(_11984_),
    .X(_11985_));
 sky130_fd_sc_hd__a31o_1 _27159_ (.A1(_11974_),
    .A2(\datamem.data_ram[49][0] ),
    .A3(_11983_),
    .B1(_11985_),
    .X(_03463_));
 sky130_fd_sc_hd__and2_1 _27160_ (.A(_11968_),
    .B(_11984_),
    .X(_11986_));
 sky130_fd_sc_hd__a31o_1 _27161_ (.A1(_11974_),
    .A2(\datamem.data_ram[49][1] ),
    .A3(_11983_),
    .B1(_11986_),
    .X(_03464_));
 sky130_fd_sc_hd__and2_1 _27162_ (.A(_11970_),
    .B(_11984_),
    .X(_11987_));
 sky130_fd_sc_hd__a31o_1 _27163_ (.A1(_11974_),
    .A2(\datamem.data_ram[49][2] ),
    .A3(_11983_),
    .B1(_11987_),
    .X(_03465_));
 sky130_fd_sc_hd__and2_1 _27164_ (.A(_11972_),
    .B(_11984_),
    .X(_11988_));
 sky130_fd_sc_hd__a31o_1 _27165_ (.A1(_11974_),
    .A2(\datamem.data_ram[49][3] ),
    .A3(_11983_),
    .B1(_11988_),
    .X(_03466_));
 sky130_fd_sc_hd__and2_1 _27166_ (.A(_11946_),
    .B(_11984_),
    .X(_11989_));
 sky130_fd_sc_hd__a31o_1 _27167_ (.A1(_11974_),
    .A2(\datamem.data_ram[49][4] ),
    .A3(_11983_),
    .B1(_11989_),
    .X(_03467_));
 sky130_fd_sc_hd__and2_1 _27168_ (.A(_11976_),
    .B(_11984_),
    .X(_11990_));
 sky130_fd_sc_hd__a31o_1 _27169_ (.A1(_11974_),
    .A2(\datamem.data_ram[49][5] ),
    .A3(_11983_),
    .B1(_11990_),
    .X(_03468_));
 sky130_fd_sc_hd__buf_2 _27170_ (.A(_11918_),
    .X(_11991_));
 sky130_fd_sc_hd__and2_1 _27171_ (.A(_11978_),
    .B(_11984_),
    .X(_11992_));
 sky130_fd_sc_hd__a31o_1 _27172_ (.A1(_11991_),
    .A2(\datamem.data_ram[49][6] ),
    .A3(_11983_),
    .B1(_11992_),
    .X(_03469_));
 sky130_fd_sc_hd__and2_1 _27173_ (.A(_11980_),
    .B(_11984_),
    .X(_11993_));
 sky130_fd_sc_hd__a31o_1 _27174_ (.A1(_11991_),
    .A2(\datamem.data_ram[49][7] ),
    .A3(_11983_),
    .B1(_11993_),
    .X(_03470_));
 sky130_fd_sc_hd__or3_1 _27175_ (.A(_07028_),
    .B(_11109_),
    .C(_11839_),
    .X(_11994_));
 sky130_fd_sc_hd__buf_2 _27176_ (.A(_11994_),
    .X(_11995_));
 sky130_fd_sc_hd__and3_1 _27177_ (.A(_09226_),
    .B(_11112_),
    .C(_11898_),
    .X(_11996_));
 sky130_fd_sc_hd__and2_1 _27178_ (.A(_11965_),
    .B(_11996_),
    .X(_11997_));
 sky130_fd_sc_hd__a31o_1 _27179_ (.A1(_11991_),
    .A2(\datamem.data_ram[30][0] ),
    .A3(_11995_),
    .B1(_11997_),
    .X(_03471_));
 sky130_fd_sc_hd__and2_1 _27180_ (.A(_11968_),
    .B(_11996_),
    .X(_11998_));
 sky130_fd_sc_hd__a31o_1 _27181_ (.A1(_11991_),
    .A2(\datamem.data_ram[30][1] ),
    .A3(_11995_),
    .B1(_11998_),
    .X(_03472_));
 sky130_fd_sc_hd__and2_1 _27182_ (.A(_11970_),
    .B(_11996_),
    .X(_11999_));
 sky130_fd_sc_hd__a31o_1 _27183_ (.A1(_11991_),
    .A2(\datamem.data_ram[30][2] ),
    .A3(_11995_),
    .B1(_11999_),
    .X(_03473_));
 sky130_fd_sc_hd__and2_1 _27184_ (.A(_11972_),
    .B(_11996_),
    .X(_12000_));
 sky130_fd_sc_hd__a31o_1 _27185_ (.A1(_11991_),
    .A2(\datamem.data_ram[30][3] ),
    .A3(_11995_),
    .B1(_12000_),
    .X(_03474_));
 sky130_fd_sc_hd__and2_1 _27186_ (.A(_11946_),
    .B(_11996_),
    .X(_12001_));
 sky130_fd_sc_hd__a31o_1 _27187_ (.A1(_11991_),
    .A2(\datamem.data_ram[30][4] ),
    .A3(_11995_),
    .B1(_12001_),
    .X(_03475_));
 sky130_fd_sc_hd__and2_1 _27188_ (.A(_11976_),
    .B(_11996_),
    .X(_12002_));
 sky130_fd_sc_hd__a31o_1 _27189_ (.A1(_11991_),
    .A2(\datamem.data_ram[30][5] ),
    .A3(_11995_),
    .B1(_12002_),
    .X(_03476_));
 sky130_fd_sc_hd__and2_1 _27190_ (.A(_11978_),
    .B(_11996_),
    .X(_12003_));
 sky130_fd_sc_hd__a31o_1 _27191_ (.A1(_11991_),
    .A2(\datamem.data_ram[30][6] ),
    .A3(_11995_),
    .B1(_12003_),
    .X(_03477_));
 sky130_fd_sc_hd__and2_1 _27192_ (.A(_11980_),
    .B(_11996_),
    .X(_12004_));
 sky130_fd_sc_hd__a31o_1 _27193_ (.A1(_11991_),
    .A2(\datamem.data_ram[30][7] ),
    .A3(_11995_),
    .B1(_12004_),
    .X(_03478_));
 sky130_fd_sc_hd__buf_2 _27194_ (.A(_11918_),
    .X(_12005_));
 sky130_fd_sc_hd__or2_1 _27195_ (.A(_10402_),
    .B(_10980_),
    .X(_12006_));
 sky130_fd_sc_hd__clkbuf_2 _27196_ (.A(_12006_),
    .X(_12007_));
 sky130_fd_sc_hd__nor2_2 _27197_ (.A(_10402_),
    .B(_10980_),
    .Y(_12008_));
 sky130_fd_sc_hd__and2_1 _27198_ (.A(_11965_),
    .B(_12008_),
    .X(_12009_));
 sky130_fd_sc_hd__a31o_1 _27199_ (.A1(_12005_),
    .A2(\datamem.data_ram[48][0] ),
    .A3(_12007_),
    .B1(_12009_),
    .X(_03479_));
 sky130_fd_sc_hd__and2_1 _27200_ (.A(_11968_),
    .B(_12008_),
    .X(_12010_));
 sky130_fd_sc_hd__a31o_1 _27201_ (.A1(_12005_),
    .A2(\datamem.data_ram[48][1] ),
    .A3(_12007_),
    .B1(_12010_),
    .X(_03480_));
 sky130_fd_sc_hd__and2_1 _27202_ (.A(_11970_),
    .B(_12008_),
    .X(_12011_));
 sky130_fd_sc_hd__a31o_1 _27203_ (.A1(_12005_),
    .A2(\datamem.data_ram[48][2] ),
    .A3(_12007_),
    .B1(_12011_),
    .X(_03481_));
 sky130_fd_sc_hd__and2_1 _27204_ (.A(_11972_),
    .B(_12008_),
    .X(_12012_));
 sky130_fd_sc_hd__a31o_1 _27205_ (.A1(_12005_),
    .A2(\datamem.data_ram[48][3] ),
    .A3(_12007_),
    .B1(_12012_),
    .X(_03482_));
 sky130_fd_sc_hd__and2_1 _27206_ (.A(_11946_),
    .B(_12008_),
    .X(_12013_));
 sky130_fd_sc_hd__a31o_1 _27207_ (.A1(_12005_),
    .A2(\datamem.data_ram[48][4] ),
    .A3(_12007_),
    .B1(_12013_),
    .X(_03483_));
 sky130_fd_sc_hd__and2_1 _27208_ (.A(_11976_),
    .B(_12008_),
    .X(_12014_));
 sky130_fd_sc_hd__a31o_1 _27209_ (.A1(_12005_),
    .A2(\datamem.data_ram[48][5] ),
    .A3(_12007_),
    .B1(_12014_),
    .X(_03484_));
 sky130_fd_sc_hd__and2_1 _27210_ (.A(_11978_),
    .B(_12008_),
    .X(_12015_));
 sky130_fd_sc_hd__a31o_1 _27211_ (.A1(_12005_),
    .A2(\datamem.data_ram[48][6] ),
    .A3(_12007_),
    .B1(_12015_),
    .X(_03485_));
 sky130_fd_sc_hd__and2_1 _27212_ (.A(_11980_),
    .B(_12008_),
    .X(_12016_));
 sky130_fd_sc_hd__a31o_1 _27213_ (.A1(_12005_),
    .A2(\datamem.data_ram[48][7] ),
    .A3(_12007_),
    .B1(_12016_),
    .X(_03486_));
 sky130_fd_sc_hd__or3_1 _27214_ (.A(_07019_),
    .B(_11109_),
    .C(_11839_),
    .X(_12017_));
 sky130_fd_sc_hd__clkbuf_2 _27215_ (.A(_12017_),
    .X(_12018_));
 sky130_fd_sc_hd__and3_1 _27216_ (.A(_09299_),
    .B(_11112_),
    .C(_11898_),
    .X(_12019_));
 sky130_fd_sc_hd__and2_1 _27217_ (.A(_11965_),
    .B(_12019_),
    .X(_12020_));
 sky130_fd_sc_hd__a31o_1 _27218_ (.A1(_12005_),
    .A2(\datamem.data_ram[29][0] ),
    .A3(_12018_),
    .B1(_12020_),
    .X(_03487_));
 sky130_fd_sc_hd__and2_1 _27219_ (.A(_11968_),
    .B(_12019_),
    .X(_12021_));
 sky130_fd_sc_hd__a31o_1 _27220_ (.A1(_12005_),
    .A2(\datamem.data_ram[29][1] ),
    .A3(_12018_),
    .B1(_12021_),
    .X(_03488_));
 sky130_fd_sc_hd__clkbuf_4 _27221_ (.A(_11918_),
    .X(_12022_));
 sky130_fd_sc_hd__and2_1 _27222_ (.A(_11970_),
    .B(_12019_),
    .X(_12023_));
 sky130_fd_sc_hd__a31o_1 _27223_ (.A1(_12022_),
    .A2(\datamem.data_ram[29][2] ),
    .A3(_12018_),
    .B1(_12023_),
    .X(_03489_));
 sky130_fd_sc_hd__and2_1 _27224_ (.A(_11972_),
    .B(_12019_),
    .X(_12024_));
 sky130_fd_sc_hd__a31o_1 _27225_ (.A1(_12022_),
    .A2(\datamem.data_ram[29][3] ),
    .A3(_12018_),
    .B1(_12024_),
    .X(_03490_));
 sky130_fd_sc_hd__and2_1 _27226_ (.A(_11946_),
    .B(_12019_),
    .X(_12025_));
 sky130_fd_sc_hd__a31o_1 _27227_ (.A1(_12022_),
    .A2(\datamem.data_ram[29][4] ),
    .A3(_12018_),
    .B1(_12025_),
    .X(_03491_));
 sky130_fd_sc_hd__and2_1 _27228_ (.A(_11976_),
    .B(_12019_),
    .X(_12026_));
 sky130_fd_sc_hd__a31o_1 _27229_ (.A1(_12022_),
    .A2(\datamem.data_ram[29][5] ),
    .A3(_12018_),
    .B1(_12026_),
    .X(_03492_));
 sky130_fd_sc_hd__and2_1 _27230_ (.A(_11978_),
    .B(_12019_),
    .X(_12027_));
 sky130_fd_sc_hd__a31o_1 _27231_ (.A1(_12022_),
    .A2(\datamem.data_ram[29][6] ),
    .A3(_12018_),
    .B1(_12027_),
    .X(_03493_));
 sky130_fd_sc_hd__and2_1 _27232_ (.A(_11980_),
    .B(_12019_),
    .X(_12028_));
 sky130_fd_sc_hd__a31o_1 _27233_ (.A1(_12022_),
    .A2(\datamem.data_ram[29][7] ),
    .A3(_12018_),
    .B1(_12028_),
    .X(_03494_));
 sky130_fd_sc_hd__or3_1 _27234_ (.A(_07808_),
    .B(_10043_),
    .C(_10897_),
    .X(_12029_));
 sky130_fd_sc_hd__clkbuf_2 _27235_ (.A(_12029_),
    .X(_12030_));
 sky130_fd_sc_hd__and3_1 _27236_ (.A(_10268_),
    .B(_10921_),
    .C(_10922_),
    .X(_12031_));
 sky130_fd_sc_hd__and2_1 _27237_ (.A(_11965_),
    .B(_12031_),
    .X(_12032_));
 sky130_fd_sc_hd__a31o_1 _27238_ (.A1(_12022_),
    .A2(\datamem.data_ram[33][0] ),
    .A3(_12030_),
    .B1(_12032_),
    .X(_03495_));
 sky130_fd_sc_hd__and2_1 _27239_ (.A(_11968_),
    .B(_12031_),
    .X(_12033_));
 sky130_fd_sc_hd__a31o_1 _27240_ (.A1(_12022_),
    .A2(\datamem.data_ram[33][1] ),
    .A3(_12030_),
    .B1(_12033_),
    .X(_03496_));
 sky130_fd_sc_hd__and2_1 _27241_ (.A(_11970_),
    .B(_12031_),
    .X(_12034_));
 sky130_fd_sc_hd__a31o_1 _27242_ (.A1(_12022_),
    .A2(\datamem.data_ram[33][2] ),
    .A3(_12030_),
    .B1(_12034_),
    .X(_03497_));
 sky130_fd_sc_hd__and2_1 _27243_ (.A(_11972_),
    .B(_12031_),
    .X(_12035_));
 sky130_fd_sc_hd__a31o_1 _27244_ (.A1(_12022_),
    .A2(\datamem.data_ram[33][3] ),
    .A3(_12030_),
    .B1(_12035_),
    .X(_03498_));
 sky130_fd_sc_hd__buf_2 _27245_ (.A(_11918_),
    .X(_12036_));
 sky130_fd_sc_hd__and2_1 _27246_ (.A(_11946_),
    .B(_12031_),
    .X(_12037_));
 sky130_fd_sc_hd__a31o_1 _27247_ (.A1(_12036_),
    .A2(\datamem.data_ram[33][4] ),
    .A3(_12030_),
    .B1(_12037_),
    .X(_03499_));
 sky130_fd_sc_hd__and2_1 _27248_ (.A(_11976_),
    .B(_12031_),
    .X(_12038_));
 sky130_fd_sc_hd__a31o_1 _27249_ (.A1(_12036_),
    .A2(\datamem.data_ram[33][5] ),
    .A3(_12030_),
    .B1(_12038_),
    .X(_03500_));
 sky130_fd_sc_hd__and2_1 _27250_ (.A(_11978_),
    .B(_12031_),
    .X(_12039_));
 sky130_fd_sc_hd__a31o_1 _27251_ (.A1(_12036_),
    .A2(\datamem.data_ram[33][6] ),
    .A3(_12030_),
    .B1(_12039_),
    .X(_03501_));
 sky130_fd_sc_hd__and2_1 _27252_ (.A(_11980_),
    .B(_12031_),
    .X(_12040_));
 sky130_fd_sc_hd__a31o_1 _27253_ (.A1(_12036_),
    .A2(\datamem.data_ram[33][7] ),
    .A3(_12030_),
    .B1(_12040_),
    .X(_03502_));
 sky130_fd_sc_hd__nor3_1 _27254_ (.A(_07791_),
    .B(_10043_),
    .C(_10600_),
    .Y(_12041_));
 sky130_fd_sc_hd__nor2_2 _27255_ (.A(_09231_),
    .B(net52),
    .Y(_12042_));
 sky130_fd_sc_hd__a22o_1 _27256_ (.A1(_10048_),
    .A2(net52),
    .B1(_12042_),
    .B2(\datamem.data_ram[47][0] ),
    .X(_03503_));
 sky130_fd_sc_hd__a22o_1 _27257_ (.A1(_10058_),
    .A2(net52),
    .B1(_12042_),
    .B2(\datamem.data_ram[47][1] ),
    .X(_03504_));
 sky130_fd_sc_hd__a22o_1 _27258_ (.A1(_10061_),
    .A2(net52),
    .B1(_12042_),
    .B2(\datamem.data_ram[47][2] ),
    .X(_03505_));
 sky130_fd_sc_hd__a22o_1 _27259_ (.A1(_10064_),
    .A2(net52),
    .B1(_12042_),
    .B2(\datamem.data_ram[47][3] ),
    .X(_03506_));
 sky130_fd_sc_hd__a22o_1 _27260_ (.A1(_10782_),
    .A2(net52),
    .B1(_12042_),
    .B2(\datamem.data_ram[47][4] ),
    .X(_03507_));
 sky130_fd_sc_hd__a22o_1 _27261_ (.A1(_10070_),
    .A2(net52),
    .B1(_12042_),
    .B2(\datamem.data_ram[47][5] ),
    .X(_03508_));
 sky130_fd_sc_hd__a22o_1 _27262_ (.A1(_10073_),
    .A2(_12041_),
    .B1(_12042_),
    .B2(\datamem.data_ram[47][6] ),
    .X(_03509_));
 sky130_fd_sc_hd__a22o_1 _27263_ (.A1(_10783_),
    .A2(_12041_),
    .B1(_12042_),
    .B2(\datamem.data_ram[47][7] ),
    .X(_03510_));
 sky130_fd_sc_hd__a21oi_4 _27264_ (.A1(_10838_),
    .A2(_10997_),
    .B1(_11713_),
    .Y(_12043_));
 sky130_fd_sc_hd__mux2_1 _27265_ (.A0(_10811_),
    .A1(\datamem.data_ram[8][24] ),
    .S(_12043_),
    .X(_12044_));
 sky130_fd_sc_hd__clkbuf_1 _27266_ (.A(_12044_),
    .X(_03511_));
 sky130_fd_sc_hd__mux2_1 _27267_ (.A0(_10814_),
    .A1(\datamem.data_ram[8][25] ),
    .S(_12043_),
    .X(_12045_));
 sky130_fd_sc_hd__clkbuf_1 _27268_ (.A(_12045_),
    .X(_03512_));
 sky130_fd_sc_hd__mux2_1 _27269_ (.A0(_10816_),
    .A1(\datamem.data_ram[8][26] ),
    .S(_12043_),
    .X(_12046_));
 sky130_fd_sc_hd__clkbuf_1 _27270_ (.A(_12046_),
    .X(_03513_));
 sky130_fd_sc_hd__mux2_1 _27271_ (.A0(_10818_),
    .A1(\datamem.data_ram[8][27] ),
    .S(_12043_),
    .X(_12047_));
 sky130_fd_sc_hd__clkbuf_1 _27272_ (.A(_12047_),
    .X(_03514_));
 sky130_fd_sc_hd__mux2_1 _27273_ (.A0(_10820_),
    .A1(\datamem.data_ram[8][28] ),
    .S(_12043_),
    .X(_12048_));
 sky130_fd_sc_hd__clkbuf_1 _27274_ (.A(_12048_),
    .X(_03515_));
 sky130_fd_sc_hd__mux2_1 _27275_ (.A0(_10822_),
    .A1(\datamem.data_ram[8][29] ),
    .S(_12043_),
    .X(_12049_));
 sky130_fd_sc_hd__clkbuf_1 _27276_ (.A(_12049_),
    .X(_03516_));
 sky130_fd_sc_hd__mux2_1 _27277_ (.A0(_10824_),
    .A1(\datamem.data_ram[8][30] ),
    .S(_12043_),
    .X(_12050_));
 sky130_fd_sc_hd__clkbuf_1 _27278_ (.A(_12050_),
    .X(_03517_));
 sky130_fd_sc_hd__mux2_1 _27279_ (.A0(_10826_),
    .A1(\datamem.data_ram[8][31] ),
    .S(_12043_),
    .X(_12051_));
 sky130_fd_sc_hd__clkbuf_1 _27280_ (.A(_12051_),
    .X(_03518_));
 sky130_fd_sc_hd__or3_1 _27281_ (.A(_07791_),
    .B(_08133_),
    .C(_11839_),
    .X(_12052_));
 sky130_fd_sc_hd__clkbuf_2 _27282_ (.A(_12052_),
    .X(_12053_));
 sky130_fd_sc_hd__and3_1 _27283_ (.A(_10325_),
    .B(_11054_),
    .C(_11898_),
    .X(_12054_));
 sky130_fd_sc_hd__and2_1 _27284_ (.A(_11965_),
    .B(_12054_),
    .X(_12055_));
 sky130_fd_sc_hd__a31o_1 _27285_ (.A1(_12036_),
    .A2(\datamem.data_ram[23][0] ),
    .A3(_12053_),
    .B1(_12055_),
    .X(_03519_));
 sky130_fd_sc_hd__and2_1 _27286_ (.A(_11968_),
    .B(_12054_),
    .X(_12056_));
 sky130_fd_sc_hd__a31o_1 _27287_ (.A1(_12036_),
    .A2(\datamem.data_ram[23][1] ),
    .A3(_12053_),
    .B1(_12056_),
    .X(_03520_));
 sky130_fd_sc_hd__and2_1 _27288_ (.A(_11970_),
    .B(_12054_),
    .X(_12057_));
 sky130_fd_sc_hd__a31o_1 _27289_ (.A1(_12036_),
    .A2(\datamem.data_ram[23][2] ),
    .A3(_12053_),
    .B1(_12057_),
    .X(_03521_));
 sky130_fd_sc_hd__and2_1 _27290_ (.A(_11972_),
    .B(_12054_),
    .X(_12058_));
 sky130_fd_sc_hd__a31o_1 _27291_ (.A1(_12036_),
    .A2(\datamem.data_ram[23][3] ),
    .A3(_12053_),
    .B1(_12058_),
    .X(_03522_));
 sky130_fd_sc_hd__and2_1 _27292_ (.A(_11946_),
    .B(_12054_),
    .X(_12059_));
 sky130_fd_sc_hd__a31o_1 _27293_ (.A1(_12036_),
    .A2(\datamem.data_ram[23][4] ),
    .A3(_12053_),
    .B1(_12059_),
    .X(_03523_));
 sky130_fd_sc_hd__and2_1 _27294_ (.A(_11976_),
    .B(_12054_),
    .X(_12060_));
 sky130_fd_sc_hd__a31o_1 _27295_ (.A1(_12036_),
    .A2(\datamem.data_ram[23][5] ),
    .A3(_12053_),
    .B1(_12060_),
    .X(_03524_));
 sky130_fd_sc_hd__buf_2 _27296_ (.A(_11918_),
    .X(_12061_));
 sky130_fd_sc_hd__and2_1 _27297_ (.A(_11978_),
    .B(_12054_),
    .X(_12062_));
 sky130_fd_sc_hd__a31o_1 _27298_ (.A1(_12061_),
    .A2(\datamem.data_ram[23][6] ),
    .A3(_12053_),
    .B1(_12062_),
    .X(_03525_));
 sky130_fd_sc_hd__and2_1 _27299_ (.A(_11980_),
    .B(_12054_),
    .X(_12063_));
 sky130_fd_sc_hd__a31o_1 _27300_ (.A1(_12061_),
    .A2(\datamem.data_ram[23][7] ),
    .A3(_12053_),
    .B1(_12063_),
    .X(_03526_));
 sky130_fd_sc_hd__or3_1 _27301_ (.A(_07203_),
    .B(_09227_),
    .C(_11839_),
    .X(_12064_));
 sky130_fd_sc_hd__clkbuf_2 _27302_ (.A(_12064_),
    .X(_12065_));
 sky130_fd_sc_hd__and3_1 _27303_ (.A(_10209_),
    .B(_08066_),
    .C(_11898_),
    .X(_12066_));
 sky130_fd_sc_hd__and2_1 _27304_ (.A(_11965_),
    .B(_12066_),
    .X(_12067_));
 sky130_fd_sc_hd__a31o_1 _27305_ (.A1(_12061_),
    .A2(\datamem.data_ram[58][0] ),
    .A3(_12065_),
    .B1(_12067_),
    .X(_03527_));
 sky130_fd_sc_hd__and2_1 _27306_ (.A(_11968_),
    .B(_12066_),
    .X(_12068_));
 sky130_fd_sc_hd__a31o_1 _27307_ (.A1(_12061_),
    .A2(\datamem.data_ram[58][1] ),
    .A3(_12065_),
    .B1(_12068_),
    .X(_03528_));
 sky130_fd_sc_hd__and2_1 _27308_ (.A(_11970_),
    .B(_12066_),
    .X(_12069_));
 sky130_fd_sc_hd__a31o_1 _27309_ (.A1(_12061_),
    .A2(\datamem.data_ram[58][2] ),
    .A3(_12065_),
    .B1(_12069_),
    .X(_03529_));
 sky130_fd_sc_hd__and2_1 _27310_ (.A(_11972_),
    .B(_12066_),
    .X(_12070_));
 sky130_fd_sc_hd__a31o_1 _27311_ (.A1(_12061_),
    .A2(\datamem.data_ram[58][3] ),
    .A3(_12065_),
    .B1(_12070_),
    .X(_03530_));
 sky130_fd_sc_hd__and2_1 _27312_ (.A(_11946_),
    .B(_12066_),
    .X(_12071_));
 sky130_fd_sc_hd__a31o_1 _27313_ (.A1(_12061_),
    .A2(\datamem.data_ram[58][4] ),
    .A3(_12065_),
    .B1(_12071_),
    .X(_03531_));
 sky130_fd_sc_hd__and2_1 _27314_ (.A(_11976_),
    .B(_12066_),
    .X(_12072_));
 sky130_fd_sc_hd__a31o_1 _27315_ (.A1(_12061_),
    .A2(\datamem.data_ram[58][5] ),
    .A3(_12065_),
    .B1(_12072_),
    .X(_03532_));
 sky130_fd_sc_hd__and2_1 _27316_ (.A(_11978_),
    .B(_12066_),
    .X(_12073_));
 sky130_fd_sc_hd__a31o_1 _27317_ (.A1(_12061_),
    .A2(\datamem.data_ram[58][6] ),
    .A3(_12065_),
    .B1(_12073_),
    .X(_03533_));
 sky130_fd_sc_hd__and2_1 _27318_ (.A(_11980_),
    .B(_12066_),
    .X(_12074_));
 sky130_fd_sc_hd__a31o_1 _27319_ (.A1(_12061_),
    .A2(\datamem.data_ram[58][7] ),
    .A3(_12065_),
    .B1(_12074_),
    .X(_03534_));
 sky130_fd_sc_hd__and3_1 _27320_ (.A(_10979_),
    .B(_10049_),
    .C(_10051_),
    .X(_12075_));
 sky130_fd_sc_hd__clkbuf_2 _27321_ (.A(_12075_),
    .X(_12076_));
 sky130_fd_sc_hd__nor2_2 _27322_ (.A(_10780_),
    .B(_12076_),
    .Y(_12077_));
 sky130_fd_sc_hd__a22o_1 _27323_ (.A1(_10048_),
    .A2(_12076_),
    .B1(_12077_),
    .B2(\datamem.data_ram[0][0] ),
    .X(_03535_));
 sky130_fd_sc_hd__a22o_1 _27324_ (.A1(_10058_),
    .A2(_12076_),
    .B1(_12077_),
    .B2(\datamem.data_ram[0][1] ),
    .X(_03536_));
 sky130_fd_sc_hd__or3_2 _27325_ (.A(_07191_),
    .B(_10042_),
    .C(_10044_),
    .X(_12078_));
 sky130_fd_sc_hd__nand2_1 _27326_ (.A(_11533_),
    .B(_12078_),
    .Y(_12079_));
 sky130_fd_sc_hd__o22a_1 _27327_ (.A1(_10061_),
    .A2(_12078_),
    .B1(_12079_),
    .B2(\datamem.data_ram[0][2] ),
    .X(_03537_));
 sky130_fd_sc_hd__o22a_1 _27328_ (.A1(_10064_),
    .A2(_12078_),
    .B1(_12079_),
    .B2(\datamem.data_ram[0][3] ),
    .X(_03538_));
 sky130_fd_sc_hd__o22a_1 _27329_ (.A1(_10782_),
    .A2(_12078_),
    .B1(_12079_),
    .B2(\datamem.data_ram[0][4] ),
    .X(_03539_));
 sky130_fd_sc_hd__a22o_1 _27330_ (.A1(_10070_),
    .A2(_12076_),
    .B1(_12077_),
    .B2(\datamem.data_ram[0][5] ),
    .X(_03540_));
 sky130_fd_sc_hd__a22o_1 _27331_ (.A1(_10073_),
    .A2(_12076_),
    .B1(_12077_),
    .B2(\datamem.data_ram[0][6] ),
    .X(_03541_));
 sky130_fd_sc_hd__a22o_1 _27332_ (.A1(_10783_),
    .A2(_12076_),
    .B1(_12077_),
    .B2(\datamem.data_ram[0][7] ),
    .X(_03542_));
 sky130_fd_sc_hd__clkbuf_2 _27333_ (.A(_09297_),
    .X(_12080_));
 sky130_fd_sc_hd__a21oi_4 _27334_ (.A1(_10598_),
    .A2(_11123_),
    .B1(_11713_),
    .Y(_12081_));
 sky130_fd_sc_hd__mux2_1 _27335_ (.A0(_12080_),
    .A1(\datamem.data_ram[7][24] ),
    .S(_12081_),
    .X(_12082_));
 sky130_fd_sc_hd__clkbuf_1 _27336_ (.A(_12082_),
    .X(_03543_));
 sky130_fd_sc_hd__buf_2 _27337_ (.A(_09305_),
    .X(_12083_));
 sky130_fd_sc_hd__mux2_1 _27338_ (.A0(_12083_),
    .A1(\datamem.data_ram[7][25] ),
    .S(_12081_),
    .X(_12084_));
 sky130_fd_sc_hd__clkbuf_1 _27339_ (.A(_12084_),
    .X(_03544_));
 sky130_fd_sc_hd__buf_2 _27340_ (.A(_09309_),
    .X(_12085_));
 sky130_fd_sc_hd__mux2_1 _27341_ (.A0(_12085_),
    .A1(\datamem.data_ram[7][26] ),
    .S(_12081_),
    .X(_12086_));
 sky130_fd_sc_hd__clkbuf_1 _27342_ (.A(_12086_),
    .X(_03545_));
 sky130_fd_sc_hd__buf_2 _27343_ (.A(_09313_),
    .X(_12087_));
 sky130_fd_sc_hd__mux2_1 _27344_ (.A0(_12087_),
    .A1(\datamem.data_ram[7][27] ),
    .S(_12081_),
    .X(_12088_));
 sky130_fd_sc_hd__clkbuf_1 _27345_ (.A(_12088_),
    .X(_03546_));
 sky130_fd_sc_hd__buf_2 _27346_ (.A(_09317_),
    .X(_12089_));
 sky130_fd_sc_hd__mux2_1 _27347_ (.A0(_12089_),
    .A1(\datamem.data_ram[7][28] ),
    .S(_12081_),
    .X(_12090_));
 sky130_fd_sc_hd__clkbuf_1 _27348_ (.A(_12090_),
    .X(_03547_));
 sky130_fd_sc_hd__buf_2 _27349_ (.A(_09321_),
    .X(_12091_));
 sky130_fd_sc_hd__mux2_1 _27350_ (.A0(_12091_),
    .A1(\datamem.data_ram[7][29] ),
    .S(_12081_),
    .X(_12092_));
 sky130_fd_sc_hd__clkbuf_1 _27351_ (.A(_12092_),
    .X(_03548_));
 sky130_fd_sc_hd__clkbuf_2 _27352_ (.A(_09325_),
    .X(_12093_));
 sky130_fd_sc_hd__mux2_1 _27353_ (.A0(_12093_),
    .A1(\datamem.data_ram[7][30] ),
    .S(_12081_),
    .X(_12094_));
 sky130_fd_sc_hd__clkbuf_1 _27354_ (.A(_12094_),
    .X(_03549_));
 sky130_fd_sc_hd__buf_2 _27355_ (.A(_09329_),
    .X(_12095_));
 sky130_fd_sc_hd__mux2_1 _27356_ (.A0(_12095_),
    .A1(\datamem.data_ram[7][31] ),
    .S(_12081_),
    .X(_12096_));
 sky130_fd_sc_hd__clkbuf_1 _27357_ (.A(_12096_),
    .X(_03550_));
 sky130_fd_sc_hd__a21oi_4 _27358_ (.A1(_10520_),
    .A2(_10997_),
    .B1(_11713_),
    .Y(_12097_));
 sky130_fd_sc_hd__mux2_1 _27359_ (.A0(_12080_),
    .A1(\datamem.data_ram[10][24] ),
    .S(_12097_),
    .X(_12098_));
 sky130_fd_sc_hd__clkbuf_1 _27360_ (.A(_12098_),
    .X(_03551_));
 sky130_fd_sc_hd__mux2_1 _27361_ (.A0(_12083_),
    .A1(\datamem.data_ram[10][25] ),
    .S(_12097_),
    .X(_12099_));
 sky130_fd_sc_hd__clkbuf_1 _27362_ (.A(_12099_),
    .X(_03552_));
 sky130_fd_sc_hd__mux2_1 _27363_ (.A0(_12085_),
    .A1(\datamem.data_ram[10][26] ),
    .S(_12097_),
    .X(_12100_));
 sky130_fd_sc_hd__clkbuf_1 _27364_ (.A(_12100_),
    .X(_03553_));
 sky130_fd_sc_hd__mux2_1 _27365_ (.A0(_12087_),
    .A1(\datamem.data_ram[10][27] ),
    .S(_12097_),
    .X(_12101_));
 sky130_fd_sc_hd__clkbuf_1 _27366_ (.A(_12101_),
    .X(_03554_));
 sky130_fd_sc_hd__mux2_1 _27367_ (.A0(_12089_),
    .A1(\datamem.data_ram[10][28] ),
    .S(_12097_),
    .X(_12102_));
 sky130_fd_sc_hd__clkbuf_1 _27368_ (.A(_12102_),
    .X(_03555_));
 sky130_fd_sc_hd__mux2_1 _27369_ (.A0(_12091_),
    .A1(\datamem.data_ram[10][29] ),
    .S(_12097_),
    .X(_12103_));
 sky130_fd_sc_hd__clkbuf_1 _27370_ (.A(_12103_),
    .X(_03556_));
 sky130_fd_sc_hd__mux2_1 _27371_ (.A0(_12093_),
    .A1(\datamem.data_ram[10][30] ),
    .S(_12097_),
    .X(_12104_));
 sky130_fd_sc_hd__clkbuf_1 _27372_ (.A(_12104_),
    .X(_03557_));
 sky130_fd_sc_hd__mux2_1 _27373_ (.A0(_12095_),
    .A1(\datamem.data_ram[10][31] ),
    .S(_12097_),
    .X(_12105_));
 sky130_fd_sc_hd__clkbuf_1 _27374_ (.A(_12105_),
    .X(_03558_));
 sky130_fd_sc_hd__nor2_8 _27375_ (.A(net112),
    .B(_10896_),
    .Y(_12106_));
 sky130_fd_sc_hd__a21oi_1 _27376_ (.A1(_10598_),
    .A2(_12106_),
    .B1(_11713_),
    .Y(_12107_));
 sky130_fd_sc_hd__mux2_1 _27377_ (.A0(_10724_),
    .A1(\datamem.data_ram[39][8] ),
    .S(net86),
    .X(_12108_));
 sky130_fd_sc_hd__clkbuf_1 _27378_ (.A(_12108_),
    .X(_03559_));
 sky130_fd_sc_hd__mux2_1 _27379_ (.A0(_10727_),
    .A1(\datamem.data_ram[39][9] ),
    .S(net86),
    .X(_12109_));
 sky130_fd_sc_hd__clkbuf_1 _27380_ (.A(_12109_),
    .X(_03560_));
 sky130_fd_sc_hd__mux2_1 _27381_ (.A0(_10729_),
    .A1(\datamem.data_ram[39][10] ),
    .S(net86),
    .X(_12110_));
 sky130_fd_sc_hd__clkbuf_1 _27382_ (.A(_12110_),
    .X(_03561_));
 sky130_fd_sc_hd__mux2_1 _27383_ (.A0(_10731_),
    .A1(\datamem.data_ram[39][11] ),
    .S(net86),
    .X(_12111_));
 sky130_fd_sc_hd__clkbuf_1 _27384_ (.A(_12111_),
    .X(_03562_));
 sky130_fd_sc_hd__mux2_1 _27385_ (.A0(_10733_),
    .A1(\datamem.data_ram[39][12] ),
    .S(net86),
    .X(_12112_));
 sky130_fd_sc_hd__clkbuf_1 _27386_ (.A(_12112_),
    .X(_03563_));
 sky130_fd_sc_hd__mux2_1 _27387_ (.A0(_10735_),
    .A1(\datamem.data_ram[39][13] ),
    .S(_12107_),
    .X(_12113_));
 sky130_fd_sc_hd__clkbuf_1 _27388_ (.A(_12113_),
    .X(_03564_));
 sky130_fd_sc_hd__mux2_1 _27389_ (.A0(_10737_),
    .A1(\datamem.data_ram[39][14] ),
    .S(net86),
    .X(_12114_));
 sky130_fd_sc_hd__clkbuf_1 _27390_ (.A(_12114_),
    .X(_03565_));
 sky130_fd_sc_hd__mux2_1 _27391_ (.A0(_10739_),
    .A1(\datamem.data_ram[39][15] ),
    .S(net86),
    .X(_12115_));
 sky130_fd_sc_hd__clkbuf_1 _27392_ (.A(_12115_),
    .X(_03566_));
 sky130_fd_sc_hd__a21oi_2 _27393_ (.A1(_10668_),
    .A2(_10898_),
    .B1(_11713_),
    .Y(_12116_));
 sky130_fd_sc_hd__mux2_1 _27394_ (.A0(_12080_),
    .A1(\datamem.data_ram[38][24] ),
    .S(net85),
    .X(_12117_));
 sky130_fd_sc_hd__clkbuf_1 _27395_ (.A(_12117_),
    .X(_03567_));
 sky130_fd_sc_hd__mux2_1 _27396_ (.A0(_12083_),
    .A1(\datamem.data_ram[38][25] ),
    .S(net85),
    .X(_12118_));
 sky130_fd_sc_hd__clkbuf_1 _27397_ (.A(_12118_),
    .X(_03568_));
 sky130_fd_sc_hd__mux2_1 _27398_ (.A0(_12085_),
    .A1(\datamem.data_ram[38][26] ),
    .S(net85),
    .X(_12119_));
 sky130_fd_sc_hd__clkbuf_1 _27399_ (.A(_12119_),
    .X(_03569_));
 sky130_fd_sc_hd__mux2_1 _27400_ (.A0(_12087_),
    .A1(\datamem.data_ram[38][27] ),
    .S(net85),
    .X(_12120_));
 sky130_fd_sc_hd__clkbuf_1 _27401_ (.A(_12120_),
    .X(_03570_));
 sky130_fd_sc_hd__mux2_1 _27402_ (.A0(_12089_),
    .A1(\datamem.data_ram[38][28] ),
    .S(net85),
    .X(_12121_));
 sky130_fd_sc_hd__clkbuf_1 _27403_ (.A(_12121_),
    .X(_03571_));
 sky130_fd_sc_hd__mux2_1 _27404_ (.A0(_12091_),
    .A1(\datamem.data_ram[38][29] ),
    .S(net85),
    .X(_12122_));
 sky130_fd_sc_hd__clkbuf_1 _27405_ (.A(_12122_),
    .X(_03572_));
 sky130_fd_sc_hd__mux2_1 _27406_ (.A0(_12093_),
    .A1(\datamem.data_ram[38][30] ),
    .S(_12116_),
    .X(_12123_));
 sky130_fd_sc_hd__clkbuf_1 _27407_ (.A(_12123_),
    .X(_03573_));
 sky130_fd_sc_hd__mux2_1 _27408_ (.A0(_12095_),
    .A1(\datamem.data_ram[38][31] ),
    .S(_12116_),
    .X(_12124_));
 sky130_fd_sc_hd__clkbuf_1 _27409_ (.A(_12124_),
    .X(_03574_));
 sky130_fd_sc_hd__buf_2 _27410_ (.A(_09223_),
    .X(_12125_));
 sky130_fd_sc_hd__a21oi_4 _27411_ (.A1(_10668_),
    .A2(_10908_),
    .B1(_11713_),
    .Y(_12126_));
 sky130_fd_sc_hd__mux2_1 _27412_ (.A0(_12125_),
    .A1(\datamem.data_ram[38][16] ),
    .S(_12126_),
    .X(_12127_));
 sky130_fd_sc_hd__clkbuf_1 _27413_ (.A(_12127_),
    .X(_03575_));
 sky130_fd_sc_hd__clkbuf_2 _27414_ (.A(_09235_),
    .X(_12128_));
 sky130_fd_sc_hd__mux2_1 _27415_ (.A0(_12128_),
    .A1(\datamem.data_ram[38][17] ),
    .S(_12126_),
    .X(_12129_));
 sky130_fd_sc_hd__clkbuf_1 _27416_ (.A(_12129_),
    .X(_03576_));
 sky130_fd_sc_hd__clkbuf_2 _27417_ (.A(_09239_),
    .X(_12130_));
 sky130_fd_sc_hd__mux2_1 _27418_ (.A0(_12130_),
    .A1(\datamem.data_ram[38][18] ),
    .S(_12126_),
    .X(_12131_));
 sky130_fd_sc_hd__clkbuf_1 _27419_ (.A(_12131_),
    .X(_03577_));
 sky130_fd_sc_hd__clkbuf_2 _27420_ (.A(_09243_),
    .X(_12132_));
 sky130_fd_sc_hd__mux2_1 _27421_ (.A0(_12132_),
    .A1(\datamem.data_ram[38][19] ),
    .S(_12126_),
    .X(_12133_));
 sky130_fd_sc_hd__clkbuf_1 _27422_ (.A(_12133_),
    .X(_03578_));
 sky130_fd_sc_hd__clkbuf_2 _27423_ (.A(_09247_),
    .X(_12134_));
 sky130_fd_sc_hd__mux2_1 _27424_ (.A0(_12134_),
    .A1(\datamem.data_ram[38][20] ),
    .S(_12126_),
    .X(_12135_));
 sky130_fd_sc_hd__clkbuf_1 _27425_ (.A(_12135_),
    .X(_03579_));
 sky130_fd_sc_hd__buf_2 _27426_ (.A(_09251_),
    .X(_12136_));
 sky130_fd_sc_hd__mux2_1 _27427_ (.A0(_12136_),
    .A1(\datamem.data_ram[38][21] ),
    .S(_12126_),
    .X(_12137_));
 sky130_fd_sc_hd__clkbuf_1 _27428_ (.A(_12137_),
    .X(_03580_));
 sky130_fd_sc_hd__clkbuf_2 _27429_ (.A(_09255_),
    .X(_12138_));
 sky130_fd_sc_hd__mux2_1 _27430_ (.A0(_12138_),
    .A1(\datamem.data_ram[38][22] ),
    .S(_12126_),
    .X(_12139_));
 sky130_fd_sc_hd__clkbuf_1 _27431_ (.A(_12139_),
    .X(_03581_));
 sky130_fd_sc_hd__clkbuf_2 _27432_ (.A(_09259_),
    .X(_12140_));
 sky130_fd_sc_hd__mux2_1 _27433_ (.A0(_12140_),
    .A1(\datamem.data_ram[38][23] ),
    .S(_12126_),
    .X(_12141_));
 sky130_fd_sc_hd__clkbuf_1 _27434_ (.A(_12141_),
    .X(_03582_));
 sky130_fd_sc_hd__buf_2 _27435_ (.A(_09266_),
    .X(_12142_));
 sky130_fd_sc_hd__a21oi_4 _27436_ (.A1(_10668_),
    .A2(_12106_),
    .B1(_11713_),
    .Y(_12143_));
 sky130_fd_sc_hd__mux2_1 _27437_ (.A0(_12142_),
    .A1(\datamem.data_ram[38][8] ),
    .S(net84),
    .X(_12144_));
 sky130_fd_sc_hd__clkbuf_1 _27438_ (.A(_12144_),
    .X(_03583_));
 sky130_fd_sc_hd__clkbuf_2 _27439_ (.A(_09272_),
    .X(_12145_));
 sky130_fd_sc_hd__mux2_1 _27440_ (.A0(_12145_),
    .A1(\datamem.data_ram[38][9] ),
    .S(_12143_),
    .X(_12146_));
 sky130_fd_sc_hd__clkbuf_1 _27441_ (.A(_12146_),
    .X(_03584_));
 sky130_fd_sc_hd__clkbuf_2 _27442_ (.A(_09275_),
    .X(_12147_));
 sky130_fd_sc_hd__mux2_1 _27443_ (.A0(_12147_),
    .A1(\datamem.data_ram[38][10] ),
    .S(net84),
    .X(_12148_));
 sky130_fd_sc_hd__clkbuf_1 _27444_ (.A(_12148_),
    .X(_03585_));
 sky130_fd_sc_hd__clkbuf_2 _27445_ (.A(_09278_),
    .X(_12149_));
 sky130_fd_sc_hd__mux2_1 _27446_ (.A0(_12149_),
    .A1(\datamem.data_ram[38][11] ),
    .S(net84),
    .X(_12150_));
 sky130_fd_sc_hd__clkbuf_1 _27447_ (.A(_12150_),
    .X(_03586_));
 sky130_fd_sc_hd__clkbuf_2 _27448_ (.A(_09281_),
    .X(_12151_));
 sky130_fd_sc_hd__mux2_1 _27449_ (.A0(_12151_),
    .A1(\datamem.data_ram[38][12] ),
    .S(net84),
    .X(_12152_));
 sky130_fd_sc_hd__clkbuf_1 _27450_ (.A(_12152_),
    .X(_03587_));
 sky130_fd_sc_hd__buf_2 _27451_ (.A(_09284_),
    .X(_12153_));
 sky130_fd_sc_hd__mux2_1 _27452_ (.A0(_12153_),
    .A1(\datamem.data_ram[38][13] ),
    .S(_12143_),
    .X(_12154_));
 sky130_fd_sc_hd__clkbuf_1 _27453_ (.A(_12154_),
    .X(_03588_));
 sky130_fd_sc_hd__clkbuf_2 _27454_ (.A(_09287_),
    .X(_12155_));
 sky130_fd_sc_hd__mux2_1 _27455_ (.A0(_12155_),
    .A1(\datamem.data_ram[38][14] ),
    .S(_12143_),
    .X(_12156_));
 sky130_fd_sc_hd__clkbuf_1 _27456_ (.A(_12156_),
    .X(_03589_));
 sky130_fd_sc_hd__clkbuf_2 _27457_ (.A(_09290_),
    .X(_12157_));
 sky130_fd_sc_hd__mux2_1 _27458_ (.A0(_12157_),
    .A1(\datamem.data_ram[38][15] ),
    .S(_12143_),
    .X(_12158_));
 sky130_fd_sc_hd__clkbuf_1 _27459_ (.A(_12158_),
    .X(_03590_));
 sky130_fd_sc_hd__a21oi_2 _27460_ (.A1(_10113_),
    .A2(_10898_),
    .B1(_11713_),
    .Y(_12159_));
 sky130_fd_sc_hd__mux2_1 _27461_ (.A0(_12080_),
    .A1(\datamem.data_ram[37][24] ),
    .S(net83),
    .X(_12160_));
 sky130_fd_sc_hd__clkbuf_1 _27462_ (.A(_12160_),
    .X(_03591_));
 sky130_fd_sc_hd__mux2_1 _27463_ (.A0(_12083_),
    .A1(\datamem.data_ram[37][25] ),
    .S(net83),
    .X(_12161_));
 sky130_fd_sc_hd__clkbuf_1 _27464_ (.A(_12161_),
    .X(_03592_));
 sky130_fd_sc_hd__mux2_1 _27465_ (.A0(_12085_),
    .A1(\datamem.data_ram[37][26] ),
    .S(net83),
    .X(_12162_));
 sky130_fd_sc_hd__clkbuf_1 _27466_ (.A(_12162_),
    .X(_03593_));
 sky130_fd_sc_hd__mux2_1 _27467_ (.A0(_12087_),
    .A1(\datamem.data_ram[37][27] ),
    .S(net83),
    .X(_12163_));
 sky130_fd_sc_hd__clkbuf_1 _27468_ (.A(_12163_),
    .X(_03594_));
 sky130_fd_sc_hd__mux2_1 _27469_ (.A0(_12089_),
    .A1(\datamem.data_ram[37][28] ),
    .S(net83),
    .X(_12164_));
 sky130_fd_sc_hd__clkbuf_1 _27470_ (.A(_12164_),
    .X(_03595_));
 sky130_fd_sc_hd__mux2_1 _27471_ (.A0(_12091_),
    .A1(\datamem.data_ram[37][29] ),
    .S(net83),
    .X(_12165_));
 sky130_fd_sc_hd__clkbuf_1 _27472_ (.A(_12165_),
    .X(_03596_));
 sky130_fd_sc_hd__mux2_1 _27473_ (.A0(_12093_),
    .A1(\datamem.data_ram[37][30] ),
    .S(_12159_),
    .X(_12166_));
 sky130_fd_sc_hd__clkbuf_1 _27474_ (.A(_12166_),
    .X(_03597_));
 sky130_fd_sc_hd__mux2_1 _27475_ (.A0(_12095_),
    .A1(\datamem.data_ram[37][31] ),
    .S(_12159_),
    .X(_12167_));
 sky130_fd_sc_hd__clkbuf_1 _27476_ (.A(_12167_),
    .X(_03598_));
 sky130_fd_sc_hd__buf_6 _27477_ (.A(_10500_),
    .X(_12168_));
 sky130_fd_sc_hd__a21oi_4 _27478_ (.A1(_10113_),
    .A2(_10908_),
    .B1(_12168_),
    .Y(_12169_));
 sky130_fd_sc_hd__mux2_1 _27479_ (.A0(_12125_),
    .A1(\datamem.data_ram[37][16] ),
    .S(_12169_),
    .X(_12170_));
 sky130_fd_sc_hd__clkbuf_1 _27480_ (.A(_12170_),
    .X(_03599_));
 sky130_fd_sc_hd__mux2_1 _27481_ (.A0(_12128_),
    .A1(\datamem.data_ram[37][17] ),
    .S(_12169_),
    .X(_12171_));
 sky130_fd_sc_hd__clkbuf_1 _27482_ (.A(_12171_),
    .X(_03600_));
 sky130_fd_sc_hd__mux2_1 _27483_ (.A0(_12130_),
    .A1(\datamem.data_ram[37][18] ),
    .S(_12169_),
    .X(_12172_));
 sky130_fd_sc_hd__clkbuf_1 _27484_ (.A(_12172_),
    .X(_03601_));
 sky130_fd_sc_hd__mux2_1 _27485_ (.A0(_12132_),
    .A1(\datamem.data_ram[37][19] ),
    .S(_12169_),
    .X(_12173_));
 sky130_fd_sc_hd__clkbuf_1 _27486_ (.A(_12173_),
    .X(_03602_));
 sky130_fd_sc_hd__mux2_1 _27487_ (.A0(_12134_),
    .A1(\datamem.data_ram[37][20] ),
    .S(_12169_),
    .X(_12174_));
 sky130_fd_sc_hd__clkbuf_1 _27488_ (.A(_12174_),
    .X(_03603_));
 sky130_fd_sc_hd__mux2_1 _27489_ (.A0(_12136_),
    .A1(\datamem.data_ram[37][21] ),
    .S(_12169_),
    .X(_12175_));
 sky130_fd_sc_hd__clkbuf_1 _27490_ (.A(_12175_),
    .X(_03604_));
 sky130_fd_sc_hd__mux2_1 _27491_ (.A0(_12138_),
    .A1(\datamem.data_ram[37][22] ),
    .S(_12169_),
    .X(_12176_));
 sky130_fd_sc_hd__clkbuf_1 _27492_ (.A(_12176_),
    .X(_03605_));
 sky130_fd_sc_hd__mux2_1 _27493_ (.A0(_12140_),
    .A1(\datamem.data_ram[37][23] ),
    .S(_12169_),
    .X(_12177_));
 sky130_fd_sc_hd__clkbuf_1 _27494_ (.A(_12177_),
    .X(_03606_));
 sky130_fd_sc_hd__buf_8 _27495_ (.A(_07132_),
    .X(_12178_));
 sky130_fd_sc_hd__a21oi_4 _27496_ (.A1(_12178_),
    .A2(_12106_),
    .B1(_12168_),
    .Y(_12179_));
 sky130_fd_sc_hd__mux2_1 _27497_ (.A0(_12142_),
    .A1(\datamem.data_ram[37][8] ),
    .S(_12179_),
    .X(_12180_));
 sky130_fd_sc_hd__clkbuf_1 _27498_ (.A(_12180_),
    .X(_03607_));
 sky130_fd_sc_hd__mux2_1 _27499_ (.A0(_12145_),
    .A1(\datamem.data_ram[37][9] ),
    .S(_12179_),
    .X(_12181_));
 sky130_fd_sc_hd__clkbuf_1 _27500_ (.A(_12181_),
    .X(_03608_));
 sky130_fd_sc_hd__mux2_1 _27501_ (.A0(_12147_),
    .A1(\datamem.data_ram[37][10] ),
    .S(_12179_),
    .X(_12182_));
 sky130_fd_sc_hd__clkbuf_1 _27502_ (.A(_12182_),
    .X(_03609_));
 sky130_fd_sc_hd__mux2_1 _27503_ (.A0(_12149_),
    .A1(\datamem.data_ram[37][11] ),
    .S(_12179_),
    .X(_12183_));
 sky130_fd_sc_hd__clkbuf_1 _27504_ (.A(_12183_),
    .X(_03610_));
 sky130_fd_sc_hd__mux2_1 _27505_ (.A0(_12151_),
    .A1(\datamem.data_ram[37][12] ),
    .S(_12179_),
    .X(_12184_));
 sky130_fd_sc_hd__clkbuf_1 _27506_ (.A(_12184_),
    .X(_03611_));
 sky130_fd_sc_hd__mux2_1 _27507_ (.A0(_12153_),
    .A1(\datamem.data_ram[37][13] ),
    .S(_12179_),
    .X(_12185_));
 sky130_fd_sc_hd__clkbuf_1 _27508_ (.A(_12185_),
    .X(_03612_));
 sky130_fd_sc_hd__mux2_1 _27509_ (.A0(_12155_),
    .A1(\datamem.data_ram[37][14] ),
    .S(_12179_),
    .X(_12186_));
 sky130_fd_sc_hd__clkbuf_1 _27510_ (.A(_12186_),
    .X(_03613_));
 sky130_fd_sc_hd__mux2_1 _27511_ (.A0(_12157_),
    .A1(\datamem.data_ram[37][15] ),
    .S(_12179_),
    .X(_12187_));
 sky130_fd_sc_hd__clkbuf_1 _27512_ (.A(_12187_),
    .X(_03614_));
 sky130_fd_sc_hd__a21oi_2 _27513_ (.A1(_10542_),
    .A2(_10898_),
    .B1(_12168_),
    .Y(_12188_));
 sky130_fd_sc_hd__mux2_1 _27514_ (.A0(_12080_),
    .A1(\datamem.data_ram[36][24] ),
    .S(net99),
    .X(_12189_));
 sky130_fd_sc_hd__clkbuf_1 _27515_ (.A(_12189_),
    .X(_03615_));
 sky130_fd_sc_hd__mux2_1 _27516_ (.A0(_12083_),
    .A1(\datamem.data_ram[36][25] ),
    .S(net99),
    .X(_12190_));
 sky130_fd_sc_hd__clkbuf_1 _27517_ (.A(_12190_),
    .X(_03616_));
 sky130_fd_sc_hd__mux2_1 _27518_ (.A0(_12085_),
    .A1(\datamem.data_ram[36][26] ),
    .S(net99),
    .X(_12191_));
 sky130_fd_sc_hd__clkbuf_1 _27519_ (.A(_12191_),
    .X(_03617_));
 sky130_fd_sc_hd__mux2_1 _27520_ (.A0(_12087_),
    .A1(\datamem.data_ram[36][27] ),
    .S(net99),
    .X(_12192_));
 sky130_fd_sc_hd__clkbuf_1 _27521_ (.A(_12192_),
    .X(_03618_));
 sky130_fd_sc_hd__mux2_1 _27522_ (.A0(_12089_),
    .A1(\datamem.data_ram[36][28] ),
    .S(net99),
    .X(_12193_));
 sky130_fd_sc_hd__clkbuf_1 _27523_ (.A(_12193_),
    .X(_03619_));
 sky130_fd_sc_hd__mux2_1 _27524_ (.A0(_12091_),
    .A1(\datamem.data_ram[36][29] ),
    .S(net99),
    .X(_12194_));
 sky130_fd_sc_hd__clkbuf_1 _27525_ (.A(_12194_),
    .X(_03620_));
 sky130_fd_sc_hd__mux2_1 _27526_ (.A0(_12093_),
    .A1(\datamem.data_ram[36][30] ),
    .S(_12188_),
    .X(_12195_));
 sky130_fd_sc_hd__clkbuf_1 _27527_ (.A(_12195_),
    .X(_03621_));
 sky130_fd_sc_hd__mux2_1 _27528_ (.A0(_12095_),
    .A1(\datamem.data_ram[36][31] ),
    .S(_12188_),
    .X(_12196_));
 sky130_fd_sc_hd__clkbuf_1 _27529_ (.A(_12196_),
    .X(_03622_));
 sky130_fd_sc_hd__a21oi_4 _27530_ (.A1(_10542_),
    .A2(_10908_),
    .B1(_12168_),
    .Y(_12197_));
 sky130_fd_sc_hd__mux2_1 _27531_ (.A0(_12125_),
    .A1(\datamem.data_ram[36][16] ),
    .S(_12197_),
    .X(_12198_));
 sky130_fd_sc_hd__clkbuf_1 _27532_ (.A(_12198_),
    .X(_03623_));
 sky130_fd_sc_hd__mux2_1 _27533_ (.A0(_12128_),
    .A1(\datamem.data_ram[36][17] ),
    .S(_12197_),
    .X(_12199_));
 sky130_fd_sc_hd__clkbuf_1 _27534_ (.A(_12199_),
    .X(_03624_));
 sky130_fd_sc_hd__mux2_1 _27535_ (.A0(_12130_),
    .A1(\datamem.data_ram[36][18] ),
    .S(_12197_),
    .X(_12200_));
 sky130_fd_sc_hd__clkbuf_1 _27536_ (.A(_12200_),
    .X(_03625_));
 sky130_fd_sc_hd__mux2_1 _27537_ (.A0(_12132_),
    .A1(\datamem.data_ram[36][19] ),
    .S(_12197_),
    .X(_12201_));
 sky130_fd_sc_hd__clkbuf_1 _27538_ (.A(_12201_),
    .X(_03626_));
 sky130_fd_sc_hd__mux2_1 _27539_ (.A0(_12134_),
    .A1(\datamem.data_ram[36][20] ),
    .S(_12197_),
    .X(_12202_));
 sky130_fd_sc_hd__clkbuf_1 _27540_ (.A(_12202_),
    .X(_03627_));
 sky130_fd_sc_hd__mux2_1 _27541_ (.A0(_12136_),
    .A1(\datamem.data_ram[36][21] ),
    .S(_12197_),
    .X(_12203_));
 sky130_fd_sc_hd__clkbuf_1 _27542_ (.A(_12203_),
    .X(_03628_));
 sky130_fd_sc_hd__mux2_1 _27543_ (.A0(_12138_),
    .A1(\datamem.data_ram[36][22] ),
    .S(_12197_),
    .X(_12204_));
 sky130_fd_sc_hd__clkbuf_1 _27544_ (.A(_12204_),
    .X(_03629_));
 sky130_fd_sc_hd__mux2_1 _27545_ (.A0(_12140_),
    .A1(\datamem.data_ram[36][23] ),
    .S(_12197_),
    .X(_12205_));
 sky130_fd_sc_hd__clkbuf_1 _27546_ (.A(_12205_),
    .X(_03630_));
 sky130_fd_sc_hd__a21oi_4 _27547_ (.A1(_10542_),
    .A2(_12106_),
    .B1(_12168_),
    .Y(_12206_));
 sky130_fd_sc_hd__mux2_1 _27548_ (.A0(_12142_),
    .A1(\datamem.data_ram[36][8] ),
    .S(net98),
    .X(_12207_));
 sky130_fd_sc_hd__clkbuf_1 _27549_ (.A(_12207_),
    .X(_03631_));
 sky130_fd_sc_hd__mux2_1 _27550_ (.A0(_12145_),
    .A1(\datamem.data_ram[36][9] ),
    .S(_12206_),
    .X(_12208_));
 sky130_fd_sc_hd__clkbuf_1 _27551_ (.A(_12208_),
    .X(_03632_));
 sky130_fd_sc_hd__mux2_1 _27552_ (.A0(_12147_),
    .A1(\datamem.data_ram[36][10] ),
    .S(net98),
    .X(_12209_));
 sky130_fd_sc_hd__clkbuf_1 _27553_ (.A(_12209_),
    .X(_03633_));
 sky130_fd_sc_hd__mux2_1 _27554_ (.A0(_12149_),
    .A1(\datamem.data_ram[36][11] ),
    .S(net98),
    .X(_12210_));
 sky130_fd_sc_hd__clkbuf_1 _27555_ (.A(_12210_),
    .X(_03634_));
 sky130_fd_sc_hd__mux2_1 _27556_ (.A0(_12151_),
    .A1(\datamem.data_ram[36][12] ),
    .S(net98),
    .X(_12211_));
 sky130_fd_sc_hd__clkbuf_1 _27557_ (.A(_12211_),
    .X(_03635_));
 sky130_fd_sc_hd__mux2_1 _27558_ (.A0(_12153_),
    .A1(\datamem.data_ram[36][13] ),
    .S(_12206_),
    .X(_12212_));
 sky130_fd_sc_hd__clkbuf_1 _27559_ (.A(_12212_),
    .X(_03636_));
 sky130_fd_sc_hd__mux2_1 _27560_ (.A0(_12155_),
    .A1(\datamem.data_ram[36][14] ),
    .S(_12206_),
    .X(_12213_));
 sky130_fd_sc_hd__clkbuf_1 _27561_ (.A(_12213_),
    .X(_03637_));
 sky130_fd_sc_hd__mux2_1 _27562_ (.A0(_12157_),
    .A1(\datamem.data_ram[36][15] ),
    .S(_12206_),
    .X(_12214_));
 sky130_fd_sc_hd__clkbuf_1 _27563_ (.A(_12214_),
    .X(_03638_));
 sky130_fd_sc_hd__a21oi_1 _27564_ (.A1(_10741_),
    .A2(_10898_),
    .B1(_12168_),
    .Y(_12215_));
 sky130_fd_sc_hd__mux2_1 _27565_ (.A0(_12080_),
    .A1(\datamem.data_ram[35][24] ),
    .S(net82),
    .X(_12216_));
 sky130_fd_sc_hd__clkbuf_1 _27566_ (.A(_12216_),
    .X(_03639_));
 sky130_fd_sc_hd__mux2_1 _27567_ (.A0(_12083_),
    .A1(\datamem.data_ram[35][25] ),
    .S(net82),
    .X(_12217_));
 sky130_fd_sc_hd__clkbuf_1 _27568_ (.A(_12217_),
    .X(_03640_));
 sky130_fd_sc_hd__mux2_1 _27569_ (.A0(_12085_),
    .A1(\datamem.data_ram[35][26] ),
    .S(net82),
    .X(_12218_));
 sky130_fd_sc_hd__clkbuf_1 _27570_ (.A(_12218_),
    .X(_03641_));
 sky130_fd_sc_hd__mux2_1 _27571_ (.A0(_12087_),
    .A1(\datamem.data_ram[35][27] ),
    .S(net82),
    .X(_12219_));
 sky130_fd_sc_hd__clkbuf_1 _27572_ (.A(_12219_),
    .X(_03642_));
 sky130_fd_sc_hd__mux2_1 _27573_ (.A0(_12089_),
    .A1(\datamem.data_ram[35][28] ),
    .S(net82),
    .X(_12220_));
 sky130_fd_sc_hd__clkbuf_1 _27574_ (.A(_12220_),
    .X(_03643_));
 sky130_fd_sc_hd__mux2_1 _27575_ (.A0(_12091_),
    .A1(\datamem.data_ram[35][29] ),
    .S(net82),
    .X(_12221_));
 sky130_fd_sc_hd__clkbuf_1 _27576_ (.A(_12221_),
    .X(_03644_));
 sky130_fd_sc_hd__mux2_1 _27577_ (.A0(_12093_),
    .A1(\datamem.data_ram[35][30] ),
    .S(_12215_),
    .X(_12222_));
 sky130_fd_sc_hd__clkbuf_1 _27578_ (.A(_12222_),
    .X(_03645_));
 sky130_fd_sc_hd__mux2_1 _27579_ (.A0(_12095_),
    .A1(\datamem.data_ram[35][31] ),
    .S(net82),
    .X(_12223_));
 sky130_fd_sc_hd__clkbuf_1 _27580_ (.A(_12223_),
    .X(_03646_));
 sky130_fd_sc_hd__a21oi_4 _27581_ (.A1(_10741_),
    .A2(_10908_),
    .B1(_12168_),
    .Y(_12224_));
 sky130_fd_sc_hd__mux2_1 _27582_ (.A0(_12125_),
    .A1(\datamem.data_ram[35][16] ),
    .S(_12224_),
    .X(_12225_));
 sky130_fd_sc_hd__clkbuf_1 _27583_ (.A(_12225_),
    .X(_03647_));
 sky130_fd_sc_hd__mux2_1 _27584_ (.A0(_12128_),
    .A1(\datamem.data_ram[35][17] ),
    .S(_12224_),
    .X(_12226_));
 sky130_fd_sc_hd__clkbuf_1 _27585_ (.A(_12226_),
    .X(_03648_));
 sky130_fd_sc_hd__mux2_1 _27586_ (.A0(_12130_),
    .A1(\datamem.data_ram[35][18] ),
    .S(_12224_),
    .X(_12227_));
 sky130_fd_sc_hd__clkbuf_1 _27587_ (.A(_12227_),
    .X(_03649_));
 sky130_fd_sc_hd__mux2_1 _27588_ (.A0(_12132_),
    .A1(\datamem.data_ram[35][19] ),
    .S(_12224_),
    .X(_12228_));
 sky130_fd_sc_hd__clkbuf_1 _27589_ (.A(_12228_),
    .X(_03650_));
 sky130_fd_sc_hd__mux2_1 _27590_ (.A0(_12134_),
    .A1(\datamem.data_ram[35][20] ),
    .S(_12224_),
    .X(_12229_));
 sky130_fd_sc_hd__clkbuf_1 _27591_ (.A(_12229_),
    .X(_03651_));
 sky130_fd_sc_hd__mux2_1 _27592_ (.A0(_12136_),
    .A1(\datamem.data_ram[35][21] ),
    .S(_12224_),
    .X(_12230_));
 sky130_fd_sc_hd__clkbuf_1 _27593_ (.A(_12230_),
    .X(_03652_));
 sky130_fd_sc_hd__mux2_1 _27594_ (.A0(_12138_),
    .A1(\datamem.data_ram[35][22] ),
    .S(_12224_),
    .X(_12231_));
 sky130_fd_sc_hd__clkbuf_1 _27595_ (.A(_12231_),
    .X(_03653_));
 sky130_fd_sc_hd__mux2_1 _27596_ (.A0(_12140_),
    .A1(\datamem.data_ram[35][23] ),
    .S(_12224_),
    .X(_12232_));
 sky130_fd_sc_hd__clkbuf_1 _27597_ (.A(_12232_),
    .X(_03654_));
 sky130_fd_sc_hd__a21oi_1 _27598_ (.A1(_10741_),
    .A2(_12106_),
    .B1(_12168_),
    .Y(_12233_));
 sky130_fd_sc_hd__mux2_1 _27599_ (.A0(_12142_),
    .A1(\datamem.data_ram[35][8] ),
    .S(net81),
    .X(_12234_));
 sky130_fd_sc_hd__clkbuf_1 _27600_ (.A(_12234_),
    .X(_03655_));
 sky130_fd_sc_hd__mux2_1 _27601_ (.A0(_12145_),
    .A1(\datamem.data_ram[35][9] ),
    .S(net81),
    .X(_12235_));
 sky130_fd_sc_hd__clkbuf_1 _27602_ (.A(_12235_),
    .X(_03656_));
 sky130_fd_sc_hd__mux2_1 _27603_ (.A0(_12147_),
    .A1(\datamem.data_ram[35][10] ),
    .S(net81),
    .X(_12236_));
 sky130_fd_sc_hd__clkbuf_1 _27604_ (.A(_12236_),
    .X(_03657_));
 sky130_fd_sc_hd__mux2_1 _27605_ (.A0(_12149_),
    .A1(\datamem.data_ram[35][11] ),
    .S(net81),
    .X(_12237_));
 sky130_fd_sc_hd__clkbuf_1 _27606_ (.A(_12237_),
    .X(_03658_));
 sky130_fd_sc_hd__mux2_1 _27607_ (.A0(_12151_),
    .A1(\datamem.data_ram[35][12] ),
    .S(net81),
    .X(_12238_));
 sky130_fd_sc_hd__clkbuf_1 _27608_ (.A(_12238_),
    .X(_03659_));
 sky130_fd_sc_hd__mux2_1 _27609_ (.A0(_12153_),
    .A1(\datamem.data_ram[35][13] ),
    .S(net81),
    .X(_12239_));
 sky130_fd_sc_hd__clkbuf_1 _27610_ (.A(_12239_),
    .X(_03660_));
 sky130_fd_sc_hd__mux2_1 _27611_ (.A0(_12155_),
    .A1(\datamem.data_ram[35][14] ),
    .S(_12233_),
    .X(_12240_));
 sky130_fd_sc_hd__clkbuf_1 _27612_ (.A(_12240_),
    .X(_03661_));
 sky130_fd_sc_hd__mux2_1 _27613_ (.A0(_12157_),
    .A1(\datamem.data_ram[35][15] ),
    .S(net81),
    .X(_12241_));
 sky130_fd_sc_hd__clkbuf_1 _27614_ (.A(_12241_),
    .X(_03662_));
 sky130_fd_sc_hd__a21oi_1 _27615_ (.A1(_10520_),
    .A2(_10898_),
    .B1(_12168_),
    .Y(_12242_));
 sky130_fd_sc_hd__mux2_1 _27616_ (.A0(_12080_),
    .A1(\datamem.data_ram[34][24] ),
    .S(net80),
    .X(_12243_));
 sky130_fd_sc_hd__clkbuf_1 _27617_ (.A(_12243_),
    .X(_03663_));
 sky130_fd_sc_hd__mux2_1 _27618_ (.A0(_12083_),
    .A1(\datamem.data_ram[34][25] ),
    .S(net80),
    .X(_12244_));
 sky130_fd_sc_hd__clkbuf_1 _27619_ (.A(_12244_),
    .X(_03664_));
 sky130_fd_sc_hd__mux2_1 _27620_ (.A0(_12085_),
    .A1(\datamem.data_ram[34][26] ),
    .S(net80),
    .X(_12245_));
 sky130_fd_sc_hd__clkbuf_1 _27621_ (.A(_12245_),
    .X(_03665_));
 sky130_fd_sc_hd__mux2_1 _27622_ (.A0(_12087_),
    .A1(\datamem.data_ram[34][27] ),
    .S(net80),
    .X(_12246_));
 sky130_fd_sc_hd__clkbuf_1 _27623_ (.A(_12246_),
    .X(_03666_));
 sky130_fd_sc_hd__mux2_1 _27624_ (.A0(_12089_),
    .A1(\datamem.data_ram[34][28] ),
    .S(net80),
    .X(_12247_));
 sky130_fd_sc_hd__clkbuf_1 _27625_ (.A(_12247_),
    .X(_03667_));
 sky130_fd_sc_hd__mux2_1 _27626_ (.A0(_12091_),
    .A1(\datamem.data_ram[34][29] ),
    .S(net80),
    .X(_12248_));
 sky130_fd_sc_hd__clkbuf_1 _27627_ (.A(_12248_),
    .X(_03668_));
 sky130_fd_sc_hd__mux2_1 _27628_ (.A0(_12093_),
    .A1(\datamem.data_ram[34][30] ),
    .S(_12242_),
    .X(_12249_));
 sky130_fd_sc_hd__clkbuf_1 _27629_ (.A(_12249_),
    .X(_03669_));
 sky130_fd_sc_hd__mux2_1 _27630_ (.A0(_12095_),
    .A1(\datamem.data_ram[34][31] ),
    .S(net80),
    .X(_12250_));
 sky130_fd_sc_hd__clkbuf_1 _27631_ (.A(_12250_),
    .X(_03670_));
 sky130_fd_sc_hd__a21oi_4 _27632_ (.A1(_10520_),
    .A2(_10908_),
    .B1(_12168_),
    .Y(_12251_));
 sky130_fd_sc_hd__mux2_1 _27633_ (.A0(_12125_),
    .A1(\datamem.data_ram[34][16] ),
    .S(_12251_),
    .X(_12252_));
 sky130_fd_sc_hd__clkbuf_1 _27634_ (.A(_12252_),
    .X(_03671_));
 sky130_fd_sc_hd__mux2_1 _27635_ (.A0(_12128_),
    .A1(\datamem.data_ram[34][17] ),
    .S(_12251_),
    .X(_12253_));
 sky130_fd_sc_hd__clkbuf_1 _27636_ (.A(_12253_),
    .X(_03672_));
 sky130_fd_sc_hd__mux2_1 _27637_ (.A0(_12130_),
    .A1(\datamem.data_ram[34][18] ),
    .S(_12251_),
    .X(_12254_));
 sky130_fd_sc_hd__clkbuf_1 _27638_ (.A(_12254_),
    .X(_03673_));
 sky130_fd_sc_hd__mux2_1 _27639_ (.A0(_12132_),
    .A1(\datamem.data_ram[34][19] ),
    .S(_12251_),
    .X(_12255_));
 sky130_fd_sc_hd__clkbuf_1 _27640_ (.A(_12255_),
    .X(_03674_));
 sky130_fd_sc_hd__mux2_1 _27641_ (.A0(_12134_),
    .A1(\datamem.data_ram[34][20] ),
    .S(_12251_),
    .X(_12256_));
 sky130_fd_sc_hd__clkbuf_1 _27642_ (.A(_12256_),
    .X(_03675_));
 sky130_fd_sc_hd__mux2_1 _27643_ (.A0(_12136_),
    .A1(\datamem.data_ram[34][21] ),
    .S(_12251_),
    .X(_12257_));
 sky130_fd_sc_hd__clkbuf_1 _27644_ (.A(_12257_),
    .X(_03676_));
 sky130_fd_sc_hd__mux2_1 _27645_ (.A0(_12138_),
    .A1(\datamem.data_ram[34][22] ),
    .S(_12251_),
    .X(_12258_));
 sky130_fd_sc_hd__clkbuf_1 _27646_ (.A(_12258_),
    .X(_03677_));
 sky130_fd_sc_hd__mux2_1 _27647_ (.A0(_12140_),
    .A1(\datamem.data_ram[34][23] ),
    .S(_12251_),
    .X(_12259_));
 sky130_fd_sc_hd__clkbuf_1 _27648_ (.A(_12259_),
    .X(_03678_));
 sky130_fd_sc_hd__buf_6 _27649_ (.A(_10500_),
    .X(_12260_));
 sky130_fd_sc_hd__a21oi_1 _27650_ (.A1(_10520_),
    .A2(_12106_),
    .B1(_12260_),
    .Y(_12261_));
 sky130_fd_sc_hd__mux2_1 _27651_ (.A0(_12142_),
    .A1(\datamem.data_ram[34][8] ),
    .S(net79),
    .X(_12262_));
 sky130_fd_sc_hd__clkbuf_1 _27652_ (.A(_12262_),
    .X(_03679_));
 sky130_fd_sc_hd__mux2_1 _27653_ (.A0(_12145_),
    .A1(\datamem.data_ram[34][9] ),
    .S(net79),
    .X(_12263_));
 sky130_fd_sc_hd__clkbuf_1 _27654_ (.A(_12263_),
    .X(_03680_));
 sky130_fd_sc_hd__mux2_1 _27655_ (.A0(_12147_),
    .A1(\datamem.data_ram[34][10] ),
    .S(net79),
    .X(_12264_));
 sky130_fd_sc_hd__clkbuf_1 _27656_ (.A(_12264_),
    .X(_03681_));
 sky130_fd_sc_hd__mux2_1 _27657_ (.A0(_12149_),
    .A1(\datamem.data_ram[34][11] ),
    .S(net79),
    .X(_12265_));
 sky130_fd_sc_hd__clkbuf_1 _27658_ (.A(_12265_),
    .X(_03682_));
 sky130_fd_sc_hd__mux2_1 _27659_ (.A0(_12151_),
    .A1(\datamem.data_ram[34][12] ),
    .S(net79),
    .X(_12266_));
 sky130_fd_sc_hd__clkbuf_1 _27660_ (.A(_12266_),
    .X(_03683_));
 sky130_fd_sc_hd__mux2_1 _27661_ (.A0(_12153_),
    .A1(\datamem.data_ram[34][13] ),
    .S(net79),
    .X(_12267_));
 sky130_fd_sc_hd__clkbuf_1 _27662_ (.A(_12267_),
    .X(_03684_));
 sky130_fd_sc_hd__mux2_1 _27663_ (.A0(_12155_),
    .A1(\datamem.data_ram[34][14] ),
    .S(_12261_),
    .X(_12268_));
 sky130_fd_sc_hd__clkbuf_1 _27664_ (.A(_12268_),
    .X(_03685_));
 sky130_fd_sc_hd__mux2_1 _27665_ (.A0(_12157_),
    .A1(\datamem.data_ram[34][15] ),
    .S(net79),
    .X(_12269_));
 sky130_fd_sc_hd__clkbuf_1 _27666_ (.A(_12269_),
    .X(_03686_));
 sky130_fd_sc_hd__a21oi_1 _27667_ (.A1(_10570_),
    .A2(_10898_),
    .B1(_12260_),
    .Y(_12270_));
 sky130_fd_sc_hd__mux2_1 _27668_ (.A0(_12080_),
    .A1(\datamem.data_ram[33][24] ),
    .S(net51),
    .X(_12271_));
 sky130_fd_sc_hd__clkbuf_1 _27669_ (.A(_12271_),
    .X(_03687_));
 sky130_fd_sc_hd__mux2_1 _27670_ (.A0(_12083_),
    .A1(\datamem.data_ram[33][25] ),
    .S(net51),
    .X(_12272_));
 sky130_fd_sc_hd__clkbuf_1 _27671_ (.A(_12272_),
    .X(_03688_));
 sky130_fd_sc_hd__mux2_1 _27672_ (.A0(_12085_),
    .A1(\datamem.data_ram[33][26] ),
    .S(net51),
    .X(_12273_));
 sky130_fd_sc_hd__clkbuf_1 _27673_ (.A(_12273_),
    .X(_03689_));
 sky130_fd_sc_hd__mux2_1 _27674_ (.A0(_12087_),
    .A1(\datamem.data_ram[33][27] ),
    .S(net51),
    .X(_12274_));
 sky130_fd_sc_hd__clkbuf_1 _27675_ (.A(_12274_),
    .X(_03690_));
 sky130_fd_sc_hd__mux2_1 _27676_ (.A0(_12089_),
    .A1(\datamem.data_ram[33][28] ),
    .S(net51),
    .X(_12275_));
 sky130_fd_sc_hd__clkbuf_1 _27677_ (.A(_12275_),
    .X(_03691_));
 sky130_fd_sc_hd__mux2_1 _27678_ (.A0(_12091_),
    .A1(\datamem.data_ram[33][29] ),
    .S(net51),
    .X(_12276_));
 sky130_fd_sc_hd__clkbuf_1 _27679_ (.A(_12276_),
    .X(_03692_));
 sky130_fd_sc_hd__mux2_1 _27680_ (.A0(_12093_),
    .A1(\datamem.data_ram[33][30] ),
    .S(_12270_),
    .X(_12277_));
 sky130_fd_sc_hd__clkbuf_1 _27681_ (.A(_12277_),
    .X(_03693_));
 sky130_fd_sc_hd__mux2_1 _27682_ (.A0(_12095_),
    .A1(\datamem.data_ram[33][31] ),
    .S(net51),
    .X(_12278_));
 sky130_fd_sc_hd__clkbuf_1 _27683_ (.A(_12278_),
    .X(_03694_));
 sky130_fd_sc_hd__buf_8 _27684_ (.A(_06997_),
    .X(_12279_));
 sky130_fd_sc_hd__a21oi_4 _27685_ (.A1(_12279_),
    .A2(_10908_),
    .B1(_12260_),
    .Y(_12280_));
 sky130_fd_sc_hd__mux2_1 _27686_ (.A0(_12125_),
    .A1(\datamem.data_ram[33][16] ),
    .S(_12280_),
    .X(_12281_));
 sky130_fd_sc_hd__clkbuf_1 _27687_ (.A(_12281_),
    .X(_03695_));
 sky130_fd_sc_hd__mux2_1 _27688_ (.A0(_12128_),
    .A1(\datamem.data_ram[33][17] ),
    .S(_12280_),
    .X(_12282_));
 sky130_fd_sc_hd__clkbuf_1 _27689_ (.A(_12282_),
    .X(_03696_));
 sky130_fd_sc_hd__mux2_1 _27690_ (.A0(_12130_),
    .A1(\datamem.data_ram[33][18] ),
    .S(_12280_),
    .X(_12283_));
 sky130_fd_sc_hd__clkbuf_1 _27691_ (.A(_12283_),
    .X(_03697_));
 sky130_fd_sc_hd__mux2_1 _27692_ (.A0(_12132_),
    .A1(\datamem.data_ram[33][19] ),
    .S(_12280_),
    .X(_12284_));
 sky130_fd_sc_hd__clkbuf_1 _27693_ (.A(_12284_),
    .X(_03698_));
 sky130_fd_sc_hd__mux2_1 _27694_ (.A0(_12134_),
    .A1(\datamem.data_ram[33][20] ),
    .S(_12280_),
    .X(_12285_));
 sky130_fd_sc_hd__clkbuf_1 _27695_ (.A(_12285_),
    .X(_03699_));
 sky130_fd_sc_hd__mux2_1 _27696_ (.A0(_12136_),
    .A1(\datamem.data_ram[33][21] ),
    .S(_12280_),
    .X(_12286_));
 sky130_fd_sc_hd__clkbuf_1 _27697_ (.A(_12286_),
    .X(_03700_));
 sky130_fd_sc_hd__mux2_1 _27698_ (.A0(_12138_),
    .A1(\datamem.data_ram[33][22] ),
    .S(_12280_),
    .X(_12287_));
 sky130_fd_sc_hd__clkbuf_1 _27699_ (.A(_12287_),
    .X(_03701_));
 sky130_fd_sc_hd__mux2_1 _27700_ (.A0(_12140_),
    .A1(\datamem.data_ram[33][23] ),
    .S(_12280_),
    .X(_12288_));
 sky130_fd_sc_hd__clkbuf_1 _27701_ (.A(_12288_),
    .X(_03702_));
 sky130_fd_sc_hd__a21oi_4 _27702_ (.A1(_12279_),
    .A2(_12106_),
    .B1(_12260_),
    .Y(_12289_));
 sky130_fd_sc_hd__mux2_1 _27703_ (.A0(_12142_),
    .A1(\datamem.data_ram[33][8] ),
    .S(_12289_),
    .X(_12290_));
 sky130_fd_sc_hd__clkbuf_1 _27704_ (.A(_12290_),
    .X(_03703_));
 sky130_fd_sc_hd__mux2_1 _27705_ (.A0(_12145_),
    .A1(\datamem.data_ram[33][9] ),
    .S(net50),
    .X(_12291_));
 sky130_fd_sc_hd__clkbuf_1 _27706_ (.A(_12291_),
    .X(_03704_));
 sky130_fd_sc_hd__mux2_1 _27707_ (.A0(_12147_),
    .A1(\datamem.data_ram[33][10] ),
    .S(_12289_),
    .X(_12292_));
 sky130_fd_sc_hd__clkbuf_1 _27708_ (.A(_12292_),
    .X(_03705_));
 sky130_fd_sc_hd__mux2_1 _27709_ (.A0(_12149_),
    .A1(\datamem.data_ram[33][11] ),
    .S(net50),
    .X(_12293_));
 sky130_fd_sc_hd__clkbuf_1 _27710_ (.A(_12293_),
    .X(_03706_));
 sky130_fd_sc_hd__mux2_1 _27711_ (.A0(_12151_),
    .A1(\datamem.data_ram[33][12] ),
    .S(_12289_),
    .X(_12294_));
 sky130_fd_sc_hd__clkbuf_1 _27712_ (.A(_12294_),
    .X(_03707_));
 sky130_fd_sc_hd__mux2_1 _27713_ (.A0(_12153_),
    .A1(\datamem.data_ram[33][13] ),
    .S(net50),
    .X(_12295_));
 sky130_fd_sc_hd__clkbuf_1 _27714_ (.A(_12295_),
    .X(_03708_));
 sky130_fd_sc_hd__mux2_1 _27715_ (.A0(_12155_),
    .A1(\datamem.data_ram[33][14] ),
    .S(net50),
    .X(_12296_));
 sky130_fd_sc_hd__clkbuf_1 _27716_ (.A(_12296_),
    .X(_03709_));
 sky130_fd_sc_hd__mux2_1 _27717_ (.A0(_12157_),
    .A1(\datamem.data_ram[33][15] ),
    .S(net50),
    .X(_12297_));
 sky130_fd_sc_hd__clkbuf_1 _27718_ (.A(_12297_),
    .X(_03710_));
 sky130_fd_sc_hd__a21oi_1 _27719_ (.A1(_10838_),
    .A2(_10898_),
    .B1(_12260_),
    .Y(_12298_));
 sky130_fd_sc_hd__mux2_1 _27720_ (.A0(_12080_),
    .A1(\datamem.data_ram[32][24] ),
    .S(net49),
    .X(_12299_));
 sky130_fd_sc_hd__clkbuf_1 _27721_ (.A(_12299_),
    .X(_03711_));
 sky130_fd_sc_hd__mux2_1 _27722_ (.A0(_12083_),
    .A1(\datamem.data_ram[32][25] ),
    .S(net49),
    .X(_12300_));
 sky130_fd_sc_hd__clkbuf_1 _27723_ (.A(_12300_),
    .X(_03712_));
 sky130_fd_sc_hd__mux2_1 _27724_ (.A0(_12085_),
    .A1(\datamem.data_ram[32][26] ),
    .S(net49),
    .X(_12301_));
 sky130_fd_sc_hd__clkbuf_1 _27725_ (.A(_12301_),
    .X(_03713_));
 sky130_fd_sc_hd__mux2_1 _27726_ (.A0(_12087_),
    .A1(\datamem.data_ram[32][27] ),
    .S(net49),
    .X(_12302_));
 sky130_fd_sc_hd__clkbuf_1 _27727_ (.A(_12302_),
    .X(_03714_));
 sky130_fd_sc_hd__mux2_1 _27728_ (.A0(_12089_),
    .A1(\datamem.data_ram[32][28] ),
    .S(net49),
    .X(_12303_));
 sky130_fd_sc_hd__clkbuf_1 _27729_ (.A(_12303_),
    .X(_03715_));
 sky130_fd_sc_hd__mux2_1 _27730_ (.A0(_12091_),
    .A1(\datamem.data_ram[32][29] ),
    .S(net49),
    .X(_12304_));
 sky130_fd_sc_hd__clkbuf_1 _27731_ (.A(_12304_),
    .X(_03716_));
 sky130_fd_sc_hd__mux2_1 _27732_ (.A0(_12093_),
    .A1(\datamem.data_ram[32][30] ),
    .S(_12298_),
    .X(_12305_));
 sky130_fd_sc_hd__clkbuf_1 _27733_ (.A(_12305_),
    .X(_03717_));
 sky130_fd_sc_hd__mux2_1 _27734_ (.A0(_12095_),
    .A1(\datamem.data_ram[32][31] ),
    .S(net49),
    .X(_12306_));
 sky130_fd_sc_hd__clkbuf_1 _27735_ (.A(_12306_),
    .X(_03718_));
 sky130_fd_sc_hd__a21oi_4 _27736_ (.A1(_10838_),
    .A2(_10908_),
    .B1(_12260_),
    .Y(_12307_));
 sky130_fd_sc_hd__mux2_1 _27737_ (.A0(_12125_),
    .A1(\datamem.data_ram[32][16] ),
    .S(_12307_),
    .X(_12308_));
 sky130_fd_sc_hd__clkbuf_1 _27738_ (.A(_12308_),
    .X(_03719_));
 sky130_fd_sc_hd__mux2_1 _27739_ (.A0(_12128_),
    .A1(\datamem.data_ram[32][17] ),
    .S(_12307_),
    .X(_12309_));
 sky130_fd_sc_hd__clkbuf_1 _27740_ (.A(_12309_),
    .X(_03720_));
 sky130_fd_sc_hd__mux2_1 _27741_ (.A0(_12130_),
    .A1(\datamem.data_ram[32][18] ),
    .S(_12307_),
    .X(_12310_));
 sky130_fd_sc_hd__clkbuf_1 _27742_ (.A(_12310_),
    .X(_03721_));
 sky130_fd_sc_hd__mux2_1 _27743_ (.A0(_12132_),
    .A1(\datamem.data_ram[32][19] ),
    .S(_12307_),
    .X(_12311_));
 sky130_fd_sc_hd__clkbuf_1 _27744_ (.A(_12311_),
    .X(_03722_));
 sky130_fd_sc_hd__mux2_1 _27745_ (.A0(_12134_),
    .A1(\datamem.data_ram[32][20] ),
    .S(_12307_),
    .X(_12312_));
 sky130_fd_sc_hd__clkbuf_1 _27746_ (.A(_12312_),
    .X(_03723_));
 sky130_fd_sc_hd__mux2_1 _27747_ (.A0(_12136_),
    .A1(\datamem.data_ram[32][21] ),
    .S(_12307_),
    .X(_12313_));
 sky130_fd_sc_hd__clkbuf_1 _27748_ (.A(_12313_),
    .X(_03724_));
 sky130_fd_sc_hd__mux2_1 _27749_ (.A0(_12138_),
    .A1(\datamem.data_ram[32][22] ),
    .S(_12307_),
    .X(_12314_));
 sky130_fd_sc_hd__clkbuf_1 _27750_ (.A(_12314_),
    .X(_03725_));
 sky130_fd_sc_hd__mux2_1 _27751_ (.A0(_12140_),
    .A1(\datamem.data_ram[32][23] ),
    .S(_12307_),
    .X(_12315_));
 sky130_fd_sc_hd__clkbuf_1 _27752_ (.A(_12315_),
    .X(_03726_));
 sky130_fd_sc_hd__a21oi_4 _27753_ (.A1(_10838_),
    .A2(_12106_),
    .B1(_12260_),
    .Y(_12316_));
 sky130_fd_sc_hd__mux2_1 _27754_ (.A0(_12142_),
    .A1(\datamem.data_ram[32][8] ),
    .S(net48),
    .X(_12317_));
 sky130_fd_sc_hd__clkbuf_1 _27755_ (.A(_12317_),
    .X(_03727_));
 sky130_fd_sc_hd__mux2_1 _27756_ (.A0(_12145_),
    .A1(\datamem.data_ram[32][9] ),
    .S(_12316_),
    .X(_12318_));
 sky130_fd_sc_hd__clkbuf_1 _27757_ (.A(_12318_),
    .X(_03728_));
 sky130_fd_sc_hd__mux2_1 _27758_ (.A0(_12147_),
    .A1(\datamem.data_ram[32][10] ),
    .S(net48),
    .X(_12319_));
 sky130_fd_sc_hd__clkbuf_1 _27759_ (.A(_12319_),
    .X(_03729_));
 sky130_fd_sc_hd__mux2_1 _27760_ (.A0(_12149_),
    .A1(\datamem.data_ram[32][11] ),
    .S(net48),
    .X(_12320_));
 sky130_fd_sc_hd__clkbuf_1 _27761_ (.A(_12320_),
    .X(_03730_));
 sky130_fd_sc_hd__mux2_1 _27762_ (.A0(_12151_),
    .A1(\datamem.data_ram[32][12] ),
    .S(net48),
    .X(_12321_));
 sky130_fd_sc_hd__clkbuf_1 _27763_ (.A(_12321_),
    .X(_03731_));
 sky130_fd_sc_hd__mux2_1 _27764_ (.A0(_12153_),
    .A1(\datamem.data_ram[32][13] ),
    .S(_12316_),
    .X(_12322_));
 sky130_fd_sc_hd__clkbuf_1 _27765_ (.A(_12322_),
    .X(_03732_));
 sky130_fd_sc_hd__mux2_1 _27766_ (.A0(_12155_),
    .A1(\datamem.data_ram[32][14] ),
    .S(_12316_),
    .X(_12323_));
 sky130_fd_sc_hd__clkbuf_1 _27767_ (.A(_12323_),
    .X(_03733_));
 sky130_fd_sc_hd__mux2_1 _27768_ (.A0(_12157_),
    .A1(\datamem.data_ram[32][15] ),
    .S(_12316_),
    .X(_12324_));
 sky130_fd_sc_hd__clkbuf_1 _27769_ (.A(_12324_),
    .X(_03734_));
 sky130_fd_sc_hd__nor2_8 _27770_ (.A(_08125_),
    .B(net111),
    .Y(_12325_));
 sky130_fd_sc_hd__a21oi_4 _27771_ (.A1(_10598_),
    .A2(_12325_),
    .B1(_12260_),
    .Y(_12326_));
 sky130_fd_sc_hd__mux2_1 _27772_ (.A0(_12080_),
    .A1(\datamem.data_ram[31][24] ),
    .S(_12326_),
    .X(_12327_));
 sky130_fd_sc_hd__clkbuf_1 _27773_ (.A(_12327_),
    .X(_03735_));
 sky130_fd_sc_hd__mux2_1 _27774_ (.A0(_12083_),
    .A1(\datamem.data_ram[31][25] ),
    .S(_12326_),
    .X(_12328_));
 sky130_fd_sc_hd__clkbuf_1 _27775_ (.A(_12328_),
    .X(_03736_));
 sky130_fd_sc_hd__mux2_1 _27776_ (.A0(_12085_),
    .A1(\datamem.data_ram[31][26] ),
    .S(_12326_),
    .X(_12329_));
 sky130_fd_sc_hd__clkbuf_1 _27777_ (.A(_12329_),
    .X(_03737_));
 sky130_fd_sc_hd__mux2_1 _27778_ (.A0(_12087_),
    .A1(\datamem.data_ram[31][27] ),
    .S(_12326_),
    .X(_12330_));
 sky130_fd_sc_hd__clkbuf_1 _27779_ (.A(_12330_),
    .X(_03738_));
 sky130_fd_sc_hd__mux2_1 _27780_ (.A0(_12089_),
    .A1(\datamem.data_ram[31][28] ),
    .S(_12326_),
    .X(_12331_));
 sky130_fd_sc_hd__clkbuf_1 _27781_ (.A(_12331_),
    .X(_03739_));
 sky130_fd_sc_hd__mux2_1 _27782_ (.A0(_12091_),
    .A1(\datamem.data_ram[31][29] ),
    .S(_12326_),
    .X(_12332_));
 sky130_fd_sc_hd__clkbuf_1 _27783_ (.A(_12332_),
    .X(_03740_));
 sky130_fd_sc_hd__mux2_1 _27784_ (.A0(_12093_),
    .A1(\datamem.data_ram[31][30] ),
    .S(_12326_),
    .X(_12333_));
 sky130_fd_sc_hd__clkbuf_1 _27785_ (.A(_12333_),
    .X(_03741_));
 sky130_fd_sc_hd__mux2_1 _27786_ (.A0(_12095_),
    .A1(\datamem.data_ram[31][31] ),
    .S(_12326_),
    .X(_12334_));
 sky130_fd_sc_hd__clkbuf_1 _27787_ (.A(_12334_),
    .X(_03742_));
 sky130_fd_sc_hd__nor2_8 _27788_ (.A(_08125_),
    .B(_09228_),
    .Y(_12335_));
 sky130_fd_sc_hd__a21oi_4 _27789_ (.A1(_10598_),
    .A2(_12335_),
    .B1(_12260_),
    .Y(_12336_));
 sky130_fd_sc_hd__mux2_1 _27790_ (.A0(_12125_),
    .A1(\datamem.data_ram[31][16] ),
    .S(_12336_),
    .X(_12337_));
 sky130_fd_sc_hd__clkbuf_1 _27791_ (.A(_12337_),
    .X(_03743_));
 sky130_fd_sc_hd__mux2_1 _27792_ (.A0(_12128_),
    .A1(\datamem.data_ram[31][17] ),
    .S(_12336_),
    .X(_12338_));
 sky130_fd_sc_hd__clkbuf_1 _27793_ (.A(_12338_),
    .X(_03744_));
 sky130_fd_sc_hd__mux2_1 _27794_ (.A0(_12130_),
    .A1(\datamem.data_ram[31][18] ),
    .S(_12336_),
    .X(_12339_));
 sky130_fd_sc_hd__clkbuf_1 _27795_ (.A(_12339_),
    .X(_03745_));
 sky130_fd_sc_hd__mux2_1 _27796_ (.A0(_12132_),
    .A1(\datamem.data_ram[31][19] ),
    .S(_12336_),
    .X(_12340_));
 sky130_fd_sc_hd__clkbuf_1 _27797_ (.A(_12340_),
    .X(_03746_));
 sky130_fd_sc_hd__mux2_1 _27798_ (.A0(_12134_),
    .A1(\datamem.data_ram[31][20] ),
    .S(_12336_),
    .X(_12341_));
 sky130_fd_sc_hd__clkbuf_1 _27799_ (.A(_12341_),
    .X(_03747_));
 sky130_fd_sc_hd__mux2_1 _27800_ (.A0(_12136_),
    .A1(\datamem.data_ram[31][21] ),
    .S(_12336_),
    .X(_12342_));
 sky130_fd_sc_hd__clkbuf_1 _27801_ (.A(_12342_),
    .X(_03748_));
 sky130_fd_sc_hd__mux2_1 _27802_ (.A0(_12138_),
    .A1(\datamem.data_ram[31][22] ),
    .S(_12336_),
    .X(_12343_));
 sky130_fd_sc_hd__clkbuf_1 _27803_ (.A(_12343_),
    .X(_03749_));
 sky130_fd_sc_hd__mux2_1 _27804_ (.A0(_12140_),
    .A1(\datamem.data_ram[31][23] ),
    .S(_12336_),
    .X(_12344_));
 sky130_fd_sc_hd__clkbuf_1 _27805_ (.A(_12344_),
    .X(_03750_));
 sky130_fd_sc_hd__nor2_2 _27806_ (.A(_08125_),
    .B(_09268_),
    .Y(_12345_));
 sky130_fd_sc_hd__a21oi_1 _27807_ (.A1(_10598_),
    .A2(_12345_),
    .B1(_12260_),
    .Y(_12346_));
 sky130_fd_sc_hd__mux2_1 _27808_ (.A0(_12142_),
    .A1(\datamem.data_ram[31][8] ),
    .S(net78),
    .X(_12347_));
 sky130_fd_sc_hd__clkbuf_1 _27809_ (.A(_12347_),
    .X(_03751_));
 sky130_fd_sc_hd__mux2_1 _27810_ (.A0(_12145_),
    .A1(\datamem.data_ram[31][9] ),
    .S(net78),
    .X(_12348_));
 sky130_fd_sc_hd__clkbuf_1 _27811_ (.A(_12348_),
    .X(_03752_));
 sky130_fd_sc_hd__mux2_1 _27812_ (.A0(_12147_),
    .A1(\datamem.data_ram[31][10] ),
    .S(net78),
    .X(_12349_));
 sky130_fd_sc_hd__clkbuf_1 _27813_ (.A(_12349_),
    .X(_03753_));
 sky130_fd_sc_hd__mux2_1 _27814_ (.A0(_12149_),
    .A1(\datamem.data_ram[31][11] ),
    .S(net78),
    .X(_12350_));
 sky130_fd_sc_hd__clkbuf_1 _27815_ (.A(_12350_),
    .X(_03754_));
 sky130_fd_sc_hd__mux2_1 _27816_ (.A0(_12151_),
    .A1(\datamem.data_ram[31][12] ),
    .S(net78),
    .X(_12351_));
 sky130_fd_sc_hd__clkbuf_1 _27817_ (.A(_12351_),
    .X(_03755_));
 sky130_fd_sc_hd__mux2_1 _27818_ (.A0(_12153_),
    .A1(\datamem.data_ram[31][13] ),
    .S(net78),
    .X(_12352_));
 sky130_fd_sc_hd__clkbuf_1 _27819_ (.A(_12352_),
    .X(_03756_));
 sky130_fd_sc_hd__mux2_1 _27820_ (.A0(_12155_),
    .A1(\datamem.data_ram[31][14] ),
    .S(net78),
    .X(_12353_));
 sky130_fd_sc_hd__clkbuf_1 _27821_ (.A(_12353_),
    .X(_03757_));
 sky130_fd_sc_hd__mux2_1 _27822_ (.A0(_12157_),
    .A1(\datamem.data_ram[31][15] ),
    .S(net78),
    .X(_12354_));
 sky130_fd_sc_hd__clkbuf_1 _27823_ (.A(_12354_),
    .X(_03758_));
 sky130_fd_sc_hd__clkbuf_2 _27824_ (.A(_09297_),
    .X(_12355_));
 sky130_fd_sc_hd__buf_6 _27825_ (.A(_10500_),
    .X(_12356_));
 sky130_fd_sc_hd__a21oi_4 _27826_ (.A1(_10668_),
    .A2(_12325_),
    .B1(_12356_),
    .Y(_12357_));
 sky130_fd_sc_hd__mux2_1 _27827_ (.A0(_12355_),
    .A1(\datamem.data_ram[30][24] ),
    .S(_12357_),
    .X(_12358_));
 sky130_fd_sc_hd__clkbuf_1 _27828_ (.A(_12358_),
    .X(_03759_));
 sky130_fd_sc_hd__clkbuf_2 _27829_ (.A(_09305_),
    .X(_12359_));
 sky130_fd_sc_hd__mux2_1 _27830_ (.A0(_12359_),
    .A1(\datamem.data_ram[30][25] ),
    .S(_12357_),
    .X(_12360_));
 sky130_fd_sc_hd__clkbuf_1 _27831_ (.A(_12360_),
    .X(_03760_));
 sky130_fd_sc_hd__clkbuf_2 _27832_ (.A(_09309_),
    .X(_12361_));
 sky130_fd_sc_hd__mux2_1 _27833_ (.A0(_12361_),
    .A1(\datamem.data_ram[30][26] ),
    .S(_12357_),
    .X(_12362_));
 sky130_fd_sc_hd__clkbuf_1 _27834_ (.A(_12362_),
    .X(_03761_));
 sky130_fd_sc_hd__clkbuf_2 _27835_ (.A(_09313_),
    .X(_12363_));
 sky130_fd_sc_hd__mux2_1 _27836_ (.A0(_12363_),
    .A1(\datamem.data_ram[30][27] ),
    .S(_12357_),
    .X(_12364_));
 sky130_fd_sc_hd__clkbuf_1 _27837_ (.A(_12364_),
    .X(_03762_));
 sky130_fd_sc_hd__buf_2 _27838_ (.A(_09317_),
    .X(_12365_));
 sky130_fd_sc_hd__mux2_1 _27839_ (.A0(_12365_),
    .A1(\datamem.data_ram[30][28] ),
    .S(_12357_),
    .X(_12366_));
 sky130_fd_sc_hd__clkbuf_1 _27840_ (.A(_12366_),
    .X(_03763_));
 sky130_fd_sc_hd__clkbuf_2 _27841_ (.A(_09321_),
    .X(_12367_));
 sky130_fd_sc_hd__mux2_1 _27842_ (.A0(_12367_),
    .A1(\datamem.data_ram[30][29] ),
    .S(_12357_),
    .X(_12368_));
 sky130_fd_sc_hd__clkbuf_1 _27843_ (.A(_12368_),
    .X(_03764_));
 sky130_fd_sc_hd__clkbuf_2 _27844_ (.A(_09325_),
    .X(_12369_));
 sky130_fd_sc_hd__mux2_1 _27845_ (.A0(_12369_),
    .A1(\datamem.data_ram[30][30] ),
    .S(_12357_),
    .X(_12370_));
 sky130_fd_sc_hd__clkbuf_1 _27846_ (.A(_12370_),
    .X(_03765_));
 sky130_fd_sc_hd__clkbuf_2 _27847_ (.A(_09329_),
    .X(_12371_));
 sky130_fd_sc_hd__mux2_1 _27848_ (.A0(_12371_),
    .A1(\datamem.data_ram[30][31] ),
    .S(_12357_),
    .X(_12372_));
 sky130_fd_sc_hd__clkbuf_1 _27849_ (.A(_12372_),
    .X(_03766_));
 sky130_fd_sc_hd__a21oi_4 _27850_ (.A1(_10668_),
    .A2(_12335_),
    .B1(_12356_),
    .Y(_12373_));
 sky130_fd_sc_hd__mux2_1 _27851_ (.A0(_12125_),
    .A1(\datamem.data_ram[30][16] ),
    .S(_12373_),
    .X(_12374_));
 sky130_fd_sc_hd__clkbuf_1 _27852_ (.A(_12374_),
    .X(_03767_));
 sky130_fd_sc_hd__mux2_1 _27853_ (.A0(_12128_),
    .A1(\datamem.data_ram[30][17] ),
    .S(_12373_),
    .X(_12375_));
 sky130_fd_sc_hd__clkbuf_1 _27854_ (.A(_12375_),
    .X(_03768_));
 sky130_fd_sc_hd__mux2_1 _27855_ (.A0(_12130_),
    .A1(\datamem.data_ram[30][18] ),
    .S(_12373_),
    .X(_12376_));
 sky130_fd_sc_hd__clkbuf_1 _27856_ (.A(_12376_),
    .X(_03769_));
 sky130_fd_sc_hd__mux2_1 _27857_ (.A0(_12132_),
    .A1(\datamem.data_ram[30][19] ),
    .S(_12373_),
    .X(_12377_));
 sky130_fd_sc_hd__clkbuf_1 _27858_ (.A(_12377_),
    .X(_03770_));
 sky130_fd_sc_hd__mux2_1 _27859_ (.A0(_12134_),
    .A1(\datamem.data_ram[30][20] ),
    .S(_12373_),
    .X(_12378_));
 sky130_fd_sc_hd__clkbuf_1 _27860_ (.A(_12378_),
    .X(_03771_));
 sky130_fd_sc_hd__mux2_1 _27861_ (.A0(_12136_),
    .A1(\datamem.data_ram[30][21] ),
    .S(_12373_),
    .X(_12379_));
 sky130_fd_sc_hd__clkbuf_1 _27862_ (.A(_12379_),
    .X(_03772_));
 sky130_fd_sc_hd__mux2_1 _27863_ (.A0(_12138_),
    .A1(\datamem.data_ram[30][22] ),
    .S(_12373_),
    .X(_12380_));
 sky130_fd_sc_hd__clkbuf_1 _27864_ (.A(_12380_),
    .X(_03773_));
 sky130_fd_sc_hd__mux2_1 _27865_ (.A0(_12140_),
    .A1(\datamem.data_ram[30][23] ),
    .S(_12373_),
    .X(_12381_));
 sky130_fd_sc_hd__clkbuf_1 _27866_ (.A(_12381_),
    .X(_03774_));
 sky130_fd_sc_hd__a21oi_2 _27867_ (.A1(_10668_),
    .A2(_12345_),
    .B1(_12356_),
    .Y(_12382_));
 sky130_fd_sc_hd__mux2_1 _27868_ (.A0(_12142_),
    .A1(\datamem.data_ram[30][8] ),
    .S(net77),
    .X(_12383_));
 sky130_fd_sc_hd__clkbuf_1 _27869_ (.A(_12383_),
    .X(_03775_));
 sky130_fd_sc_hd__mux2_1 _27870_ (.A0(_12145_),
    .A1(\datamem.data_ram[30][9] ),
    .S(net77),
    .X(_12384_));
 sky130_fd_sc_hd__clkbuf_1 _27871_ (.A(_12384_),
    .X(_03776_));
 sky130_fd_sc_hd__mux2_1 _27872_ (.A0(_12147_),
    .A1(\datamem.data_ram[30][10] ),
    .S(net77),
    .X(_12385_));
 sky130_fd_sc_hd__clkbuf_1 _27873_ (.A(_12385_),
    .X(_03777_));
 sky130_fd_sc_hd__mux2_1 _27874_ (.A0(_12149_),
    .A1(\datamem.data_ram[30][11] ),
    .S(net77),
    .X(_12386_));
 sky130_fd_sc_hd__clkbuf_1 _27875_ (.A(_12386_),
    .X(_03778_));
 sky130_fd_sc_hd__mux2_1 _27876_ (.A0(_12151_),
    .A1(\datamem.data_ram[30][12] ),
    .S(net77),
    .X(_12387_));
 sky130_fd_sc_hd__clkbuf_1 _27877_ (.A(_12387_),
    .X(_03779_));
 sky130_fd_sc_hd__mux2_1 _27878_ (.A0(_12153_),
    .A1(\datamem.data_ram[30][13] ),
    .S(net77),
    .X(_12388_));
 sky130_fd_sc_hd__clkbuf_1 _27879_ (.A(_12388_),
    .X(_03780_));
 sky130_fd_sc_hd__mux2_1 _27880_ (.A0(_12155_),
    .A1(\datamem.data_ram[30][14] ),
    .S(_12382_),
    .X(_12389_));
 sky130_fd_sc_hd__clkbuf_1 _27881_ (.A(_12389_),
    .X(_03781_));
 sky130_fd_sc_hd__mux2_1 _27882_ (.A0(_12157_),
    .A1(\datamem.data_ram[30][15] ),
    .S(_12382_),
    .X(_12390_));
 sky130_fd_sc_hd__clkbuf_1 _27883_ (.A(_12390_),
    .X(_03782_));
 sky130_fd_sc_hd__buf_2 _27884_ (.A(_11918_),
    .X(_12391_));
 sky130_fd_sc_hd__or3_1 _27885_ (.A(_07203_),
    .B(_10042_),
    .C(_10918_),
    .X(_12392_));
 sky130_fd_sc_hd__buf_2 _27886_ (.A(_12392_),
    .X(_12393_));
 sky130_fd_sc_hd__and3_2 _27887_ (.A(_10209_),
    .B(_10049_),
    .C(_11898_),
    .X(_12394_));
 sky130_fd_sc_hd__and2_1 _27888_ (.A(_11965_),
    .B(_12394_),
    .X(_12395_));
 sky130_fd_sc_hd__a31o_1 _27889_ (.A1(_12391_),
    .A2(\datamem.data_ram[2][0] ),
    .A3(_12393_),
    .B1(_12395_),
    .X(_03783_));
 sky130_fd_sc_hd__and2_1 _27890_ (.A(_11968_),
    .B(_12394_),
    .X(_12396_));
 sky130_fd_sc_hd__a31o_1 _27891_ (.A1(_12391_),
    .A2(\datamem.data_ram[2][1] ),
    .A3(_12393_),
    .B1(_12396_),
    .X(_03784_));
 sky130_fd_sc_hd__and2_1 _27892_ (.A(_11970_),
    .B(_12394_),
    .X(_12397_));
 sky130_fd_sc_hd__a31o_1 _27893_ (.A1(_12391_),
    .A2(\datamem.data_ram[2][2] ),
    .A3(_12393_),
    .B1(_12397_),
    .X(_03785_));
 sky130_fd_sc_hd__and2_1 _27894_ (.A(_11972_),
    .B(_12394_),
    .X(_12398_));
 sky130_fd_sc_hd__a31o_1 _27895_ (.A1(_12391_),
    .A2(\datamem.data_ram[2][3] ),
    .A3(_12393_),
    .B1(_12398_),
    .X(_03786_));
 sky130_fd_sc_hd__and2_1 _27896_ (.A(_10066_),
    .B(_12394_),
    .X(_12399_));
 sky130_fd_sc_hd__a31o_1 _27897_ (.A1(_12391_),
    .A2(\datamem.data_ram[2][4] ),
    .A3(_12393_),
    .B1(_12399_),
    .X(_03787_));
 sky130_fd_sc_hd__and2_1 _27898_ (.A(_11976_),
    .B(_12394_),
    .X(_12400_));
 sky130_fd_sc_hd__a31o_1 _27899_ (.A1(_12391_),
    .A2(\datamem.data_ram[2][5] ),
    .A3(_12393_),
    .B1(_12400_),
    .X(_03788_));
 sky130_fd_sc_hd__and2_1 _27900_ (.A(_11978_),
    .B(_12394_),
    .X(_12401_));
 sky130_fd_sc_hd__a31o_1 _27901_ (.A1(_12391_),
    .A2(\datamem.data_ram[2][6] ),
    .A3(_12393_),
    .B1(_12401_),
    .X(_03789_));
 sky130_fd_sc_hd__and2_1 _27902_ (.A(_11980_),
    .B(_12394_),
    .X(_12402_));
 sky130_fd_sc_hd__a31o_1 _27903_ (.A1(_12391_),
    .A2(\datamem.data_ram[2][7] ),
    .A3(_12393_),
    .B1(_12402_),
    .X(_03790_));
 sky130_fd_sc_hd__a21oi_1 _27904_ (.A1(_10520_),
    .A2(_10092_),
    .B1(_12356_),
    .Y(_12403_));
 sky130_fd_sc_hd__mux2_1 _27905_ (.A0(_12142_),
    .A1(\datamem.data_ram[2][8] ),
    .S(net47),
    .X(_12404_));
 sky130_fd_sc_hd__clkbuf_1 _27906_ (.A(_12404_),
    .X(_03791_));
 sky130_fd_sc_hd__mux2_1 _27907_ (.A0(_12145_),
    .A1(\datamem.data_ram[2][9] ),
    .S(net47),
    .X(_12405_));
 sky130_fd_sc_hd__clkbuf_1 _27908_ (.A(_12405_),
    .X(_03792_));
 sky130_fd_sc_hd__mux2_1 _27909_ (.A0(_12147_),
    .A1(\datamem.data_ram[2][10] ),
    .S(net47),
    .X(_12406_));
 sky130_fd_sc_hd__clkbuf_1 _27910_ (.A(_12406_),
    .X(_03793_));
 sky130_fd_sc_hd__mux2_1 _27911_ (.A0(_12149_),
    .A1(\datamem.data_ram[2][11] ),
    .S(net47),
    .X(_12407_));
 sky130_fd_sc_hd__clkbuf_1 _27912_ (.A(_12407_),
    .X(_03794_));
 sky130_fd_sc_hd__mux2_1 _27913_ (.A0(_12151_),
    .A1(\datamem.data_ram[2][12] ),
    .S(net47),
    .X(_12408_));
 sky130_fd_sc_hd__clkbuf_1 _27914_ (.A(_12408_),
    .X(_03795_));
 sky130_fd_sc_hd__mux2_1 _27915_ (.A0(_12153_),
    .A1(\datamem.data_ram[2][13] ),
    .S(net47),
    .X(_12409_));
 sky130_fd_sc_hd__clkbuf_1 _27916_ (.A(_12409_),
    .X(_03796_));
 sky130_fd_sc_hd__mux2_1 _27917_ (.A0(_12155_),
    .A1(\datamem.data_ram[2][14] ),
    .S(net47),
    .X(_12410_));
 sky130_fd_sc_hd__clkbuf_1 _27918_ (.A(_12410_),
    .X(_03797_));
 sky130_fd_sc_hd__mux2_1 _27919_ (.A0(_12157_),
    .A1(\datamem.data_ram[2][15] ),
    .S(net47),
    .X(_12411_));
 sky130_fd_sc_hd__clkbuf_1 _27920_ (.A(_12411_),
    .X(_03798_));
 sky130_fd_sc_hd__a21oi_4 _27921_ (.A1(_10777_),
    .A2(_10114_),
    .B1(_12356_),
    .Y(_12412_));
 sky130_fd_sc_hd__mux2_1 _27922_ (.A0(_12125_),
    .A1(\datamem.data_ram[2][16] ),
    .S(_12412_),
    .X(_12413_));
 sky130_fd_sc_hd__clkbuf_1 _27923_ (.A(_12413_),
    .X(_03799_));
 sky130_fd_sc_hd__mux2_1 _27924_ (.A0(_12128_),
    .A1(\datamem.data_ram[2][17] ),
    .S(_12412_),
    .X(_12414_));
 sky130_fd_sc_hd__clkbuf_1 _27925_ (.A(_12414_),
    .X(_03800_));
 sky130_fd_sc_hd__mux2_1 _27926_ (.A0(_12130_),
    .A1(\datamem.data_ram[2][18] ),
    .S(_12412_),
    .X(_12415_));
 sky130_fd_sc_hd__clkbuf_1 _27927_ (.A(_12415_),
    .X(_03801_));
 sky130_fd_sc_hd__mux2_1 _27928_ (.A0(_12132_),
    .A1(\datamem.data_ram[2][19] ),
    .S(_12412_),
    .X(_12416_));
 sky130_fd_sc_hd__clkbuf_1 _27929_ (.A(_12416_),
    .X(_03802_));
 sky130_fd_sc_hd__mux2_1 _27930_ (.A0(_12134_),
    .A1(\datamem.data_ram[2][20] ),
    .S(_12412_),
    .X(_12417_));
 sky130_fd_sc_hd__clkbuf_1 _27931_ (.A(_12417_),
    .X(_03803_));
 sky130_fd_sc_hd__mux2_1 _27932_ (.A0(_12136_),
    .A1(\datamem.data_ram[2][21] ),
    .S(_12412_),
    .X(_12418_));
 sky130_fd_sc_hd__clkbuf_1 _27933_ (.A(_12418_),
    .X(_03804_));
 sky130_fd_sc_hd__mux2_1 _27934_ (.A0(_12138_),
    .A1(\datamem.data_ram[2][22] ),
    .S(_12412_),
    .X(_12419_));
 sky130_fd_sc_hd__clkbuf_1 _27935_ (.A(_12419_),
    .X(_03805_));
 sky130_fd_sc_hd__mux2_1 _27936_ (.A0(_12140_),
    .A1(\datamem.data_ram[2][23] ),
    .S(_12412_),
    .X(_12420_));
 sky130_fd_sc_hd__clkbuf_1 _27937_ (.A(_12420_),
    .X(_03806_));
 sky130_fd_sc_hd__a21oi_4 _27938_ (.A1(_12178_),
    .A2(_12325_),
    .B1(_12356_),
    .Y(_12421_));
 sky130_fd_sc_hd__mux2_1 _27939_ (.A0(_12355_),
    .A1(\datamem.data_ram[29][24] ),
    .S(_12421_),
    .X(_12422_));
 sky130_fd_sc_hd__clkbuf_1 _27940_ (.A(_12422_),
    .X(_03807_));
 sky130_fd_sc_hd__mux2_1 _27941_ (.A0(_12359_),
    .A1(\datamem.data_ram[29][25] ),
    .S(_12421_),
    .X(_12423_));
 sky130_fd_sc_hd__clkbuf_1 _27942_ (.A(_12423_),
    .X(_03808_));
 sky130_fd_sc_hd__mux2_1 _27943_ (.A0(_12361_),
    .A1(\datamem.data_ram[29][26] ),
    .S(_12421_),
    .X(_12424_));
 sky130_fd_sc_hd__clkbuf_1 _27944_ (.A(_12424_),
    .X(_03809_));
 sky130_fd_sc_hd__mux2_1 _27945_ (.A0(_12363_),
    .A1(\datamem.data_ram[29][27] ),
    .S(_12421_),
    .X(_12425_));
 sky130_fd_sc_hd__clkbuf_1 _27946_ (.A(_12425_),
    .X(_03810_));
 sky130_fd_sc_hd__mux2_1 _27947_ (.A0(_12365_),
    .A1(\datamem.data_ram[29][28] ),
    .S(_12421_),
    .X(_12426_));
 sky130_fd_sc_hd__clkbuf_1 _27948_ (.A(_12426_),
    .X(_03811_));
 sky130_fd_sc_hd__mux2_1 _27949_ (.A0(_12367_),
    .A1(\datamem.data_ram[29][29] ),
    .S(_12421_),
    .X(_12427_));
 sky130_fd_sc_hd__clkbuf_1 _27950_ (.A(_12427_),
    .X(_03812_));
 sky130_fd_sc_hd__mux2_1 _27951_ (.A0(_12369_),
    .A1(\datamem.data_ram[29][30] ),
    .S(_12421_),
    .X(_12428_));
 sky130_fd_sc_hd__clkbuf_1 _27952_ (.A(_12428_),
    .X(_03813_));
 sky130_fd_sc_hd__mux2_1 _27953_ (.A0(_12371_),
    .A1(\datamem.data_ram[29][31] ),
    .S(_12421_),
    .X(_12429_));
 sky130_fd_sc_hd__clkbuf_1 _27954_ (.A(_12429_),
    .X(_03814_));
 sky130_fd_sc_hd__clkbuf_2 _27955_ (.A(_09223_),
    .X(_12430_));
 sky130_fd_sc_hd__a21oi_4 _27956_ (.A1(_12178_),
    .A2(_12335_),
    .B1(_12356_),
    .Y(_12431_));
 sky130_fd_sc_hd__mux2_1 _27957_ (.A0(_12430_),
    .A1(\datamem.data_ram[29][16] ),
    .S(_12431_),
    .X(_12432_));
 sky130_fd_sc_hd__clkbuf_1 _27958_ (.A(_12432_),
    .X(_03815_));
 sky130_fd_sc_hd__clkbuf_2 _27959_ (.A(_09235_),
    .X(_12433_));
 sky130_fd_sc_hd__mux2_1 _27960_ (.A0(_12433_),
    .A1(\datamem.data_ram[29][17] ),
    .S(_12431_),
    .X(_12434_));
 sky130_fd_sc_hd__clkbuf_1 _27961_ (.A(_12434_),
    .X(_03816_));
 sky130_fd_sc_hd__clkbuf_2 _27962_ (.A(_09239_),
    .X(_12435_));
 sky130_fd_sc_hd__mux2_1 _27963_ (.A0(_12435_),
    .A1(\datamem.data_ram[29][18] ),
    .S(_12431_),
    .X(_12436_));
 sky130_fd_sc_hd__clkbuf_1 _27964_ (.A(_12436_),
    .X(_03817_));
 sky130_fd_sc_hd__clkbuf_2 _27965_ (.A(_09243_),
    .X(_12437_));
 sky130_fd_sc_hd__mux2_1 _27966_ (.A0(_12437_),
    .A1(\datamem.data_ram[29][19] ),
    .S(_12431_),
    .X(_12438_));
 sky130_fd_sc_hd__clkbuf_1 _27967_ (.A(_12438_),
    .X(_03818_));
 sky130_fd_sc_hd__clkbuf_2 _27968_ (.A(_09247_),
    .X(_12439_));
 sky130_fd_sc_hd__mux2_1 _27969_ (.A0(_12439_),
    .A1(\datamem.data_ram[29][20] ),
    .S(_12431_),
    .X(_12440_));
 sky130_fd_sc_hd__clkbuf_1 _27970_ (.A(_12440_),
    .X(_03819_));
 sky130_fd_sc_hd__clkbuf_2 _27971_ (.A(_09251_),
    .X(_12441_));
 sky130_fd_sc_hd__mux2_1 _27972_ (.A0(_12441_),
    .A1(\datamem.data_ram[29][21] ),
    .S(_12431_),
    .X(_12442_));
 sky130_fd_sc_hd__clkbuf_1 _27973_ (.A(_12442_),
    .X(_03820_));
 sky130_fd_sc_hd__clkbuf_2 _27974_ (.A(_09255_),
    .X(_12443_));
 sky130_fd_sc_hd__mux2_1 _27975_ (.A0(_12443_),
    .A1(\datamem.data_ram[29][22] ),
    .S(_12431_),
    .X(_12444_));
 sky130_fd_sc_hd__clkbuf_1 _27976_ (.A(_12444_),
    .X(_03821_));
 sky130_fd_sc_hd__clkbuf_2 _27977_ (.A(_09259_),
    .X(_12445_));
 sky130_fd_sc_hd__mux2_1 _27978_ (.A0(_12445_),
    .A1(\datamem.data_ram[29][23] ),
    .S(_12431_),
    .X(_12446_));
 sky130_fd_sc_hd__clkbuf_1 _27979_ (.A(_12446_),
    .X(_03822_));
 sky130_fd_sc_hd__clkbuf_2 _27980_ (.A(_09266_),
    .X(_12447_));
 sky130_fd_sc_hd__a21oi_1 _27981_ (.A1(_12178_),
    .A2(_12345_),
    .B1(_12356_),
    .Y(_12448_));
 sky130_fd_sc_hd__mux2_1 _27982_ (.A0(_12447_),
    .A1(\datamem.data_ram[29][8] ),
    .S(net76),
    .X(_12449_));
 sky130_fd_sc_hd__clkbuf_1 _27983_ (.A(_12449_),
    .X(_03823_));
 sky130_fd_sc_hd__clkbuf_2 _27984_ (.A(_09272_),
    .X(_12450_));
 sky130_fd_sc_hd__mux2_1 _27985_ (.A0(_12450_),
    .A1(\datamem.data_ram[29][9] ),
    .S(net76),
    .X(_12451_));
 sky130_fd_sc_hd__clkbuf_1 _27986_ (.A(_12451_),
    .X(_03824_));
 sky130_fd_sc_hd__clkbuf_2 _27987_ (.A(_09275_),
    .X(_12452_));
 sky130_fd_sc_hd__mux2_1 _27988_ (.A0(_12452_),
    .A1(\datamem.data_ram[29][10] ),
    .S(net76),
    .X(_12453_));
 sky130_fd_sc_hd__clkbuf_1 _27989_ (.A(_12453_),
    .X(_03825_));
 sky130_fd_sc_hd__clkbuf_2 _27990_ (.A(_09278_),
    .X(_12454_));
 sky130_fd_sc_hd__mux2_1 _27991_ (.A0(_12454_),
    .A1(\datamem.data_ram[29][11] ),
    .S(net76),
    .X(_12455_));
 sky130_fd_sc_hd__clkbuf_1 _27992_ (.A(_12455_),
    .X(_03826_));
 sky130_fd_sc_hd__buf_2 _27993_ (.A(_09281_),
    .X(_12456_));
 sky130_fd_sc_hd__mux2_1 _27994_ (.A0(_12456_),
    .A1(\datamem.data_ram[29][12] ),
    .S(net76),
    .X(_12457_));
 sky130_fd_sc_hd__clkbuf_1 _27995_ (.A(_12457_),
    .X(_03827_));
 sky130_fd_sc_hd__buf_2 _27996_ (.A(_09284_),
    .X(_12458_));
 sky130_fd_sc_hd__mux2_1 _27997_ (.A0(_12458_),
    .A1(\datamem.data_ram[29][13] ),
    .S(net76),
    .X(_12459_));
 sky130_fd_sc_hd__clkbuf_1 _27998_ (.A(_12459_),
    .X(_03828_));
 sky130_fd_sc_hd__clkbuf_2 _27999_ (.A(_09287_),
    .X(_12460_));
 sky130_fd_sc_hd__mux2_1 _28000_ (.A0(_12460_),
    .A1(\datamem.data_ram[29][14] ),
    .S(net76),
    .X(_12461_));
 sky130_fd_sc_hd__clkbuf_1 _28001_ (.A(_12461_),
    .X(_03829_));
 sky130_fd_sc_hd__clkbuf_2 _28002_ (.A(_09290_),
    .X(_12462_));
 sky130_fd_sc_hd__mux2_1 _28003_ (.A0(_12462_),
    .A1(\datamem.data_ram[29][15] ),
    .S(_12448_),
    .X(_12463_));
 sky130_fd_sc_hd__clkbuf_1 _28004_ (.A(_12463_),
    .X(_03830_));
 sky130_fd_sc_hd__a21oi_1 _28005_ (.A1(_10542_),
    .A2(_12325_),
    .B1(_12356_),
    .Y(_12464_));
 sky130_fd_sc_hd__mux2_1 _28006_ (.A0(_12355_),
    .A1(\datamem.data_ram[28][24] ),
    .S(net97),
    .X(_12465_));
 sky130_fd_sc_hd__clkbuf_1 _28007_ (.A(_12465_),
    .X(_03831_));
 sky130_fd_sc_hd__mux2_1 _28008_ (.A0(_12359_),
    .A1(\datamem.data_ram[28][25] ),
    .S(net97),
    .X(_12466_));
 sky130_fd_sc_hd__clkbuf_1 _28009_ (.A(_12466_),
    .X(_03832_));
 sky130_fd_sc_hd__mux2_1 _28010_ (.A0(_12361_),
    .A1(\datamem.data_ram[28][26] ),
    .S(net97),
    .X(_12467_));
 sky130_fd_sc_hd__clkbuf_1 _28011_ (.A(_12467_),
    .X(_03833_));
 sky130_fd_sc_hd__mux2_1 _28012_ (.A0(_12363_),
    .A1(\datamem.data_ram[28][27] ),
    .S(net97),
    .X(_12468_));
 sky130_fd_sc_hd__clkbuf_1 _28013_ (.A(_12468_),
    .X(_03834_));
 sky130_fd_sc_hd__mux2_1 _28014_ (.A0(_12365_),
    .A1(\datamem.data_ram[28][28] ),
    .S(net97),
    .X(_12469_));
 sky130_fd_sc_hd__clkbuf_1 _28015_ (.A(_12469_),
    .X(_03835_));
 sky130_fd_sc_hd__mux2_1 _28016_ (.A0(_12367_),
    .A1(\datamem.data_ram[28][29] ),
    .S(net97),
    .X(_12470_));
 sky130_fd_sc_hd__clkbuf_1 _28017_ (.A(_12470_),
    .X(_03836_));
 sky130_fd_sc_hd__mux2_1 _28018_ (.A0(_12369_),
    .A1(\datamem.data_ram[28][30] ),
    .S(net97),
    .X(_12471_));
 sky130_fd_sc_hd__clkbuf_1 _28019_ (.A(_12471_),
    .X(_03837_));
 sky130_fd_sc_hd__mux2_1 _28020_ (.A0(_12371_),
    .A1(\datamem.data_ram[28][31] ),
    .S(_12464_),
    .X(_12472_));
 sky130_fd_sc_hd__clkbuf_1 _28021_ (.A(_12472_),
    .X(_03838_));
 sky130_fd_sc_hd__a21oi_4 _28022_ (.A1(_09350_),
    .A2(_12335_),
    .B1(_12356_),
    .Y(_12473_));
 sky130_fd_sc_hd__mux2_1 _28023_ (.A0(_12430_),
    .A1(\datamem.data_ram[28][16] ),
    .S(_12473_),
    .X(_12474_));
 sky130_fd_sc_hd__clkbuf_1 _28024_ (.A(_12474_),
    .X(_03839_));
 sky130_fd_sc_hd__mux2_1 _28025_ (.A0(_12433_),
    .A1(\datamem.data_ram[28][17] ),
    .S(_12473_),
    .X(_12475_));
 sky130_fd_sc_hd__clkbuf_1 _28026_ (.A(_12475_),
    .X(_03840_));
 sky130_fd_sc_hd__mux2_1 _28027_ (.A0(_12435_),
    .A1(\datamem.data_ram[28][18] ),
    .S(_12473_),
    .X(_12476_));
 sky130_fd_sc_hd__clkbuf_1 _28028_ (.A(_12476_),
    .X(_03841_));
 sky130_fd_sc_hd__mux2_1 _28029_ (.A0(_12437_),
    .A1(\datamem.data_ram[28][19] ),
    .S(_12473_),
    .X(_12477_));
 sky130_fd_sc_hd__clkbuf_1 _28030_ (.A(_12477_),
    .X(_03842_));
 sky130_fd_sc_hd__mux2_1 _28031_ (.A0(_12439_),
    .A1(\datamem.data_ram[28][20] ),
    .S(_12473_),
    .X(_12478_));
 sky130_fd_sc_hd__clkbuf_1 _28032_ (.A(_12478_),
    .X(_03843_));
 sky130_fd_sc_hd__mux2_1 _28033_ (.A0(_12441_),
    .A1(\datamem.data_ram[28][21] ),
    .S(_12473_),
    .X(_12479_));
 sky130_fd_sc_hd__clkbuf_1 _28034_ (.A(_12479_),
    .X(_03844_));
 sky130_fd_sc_hd__mux2_1 _28035_ (.A0(_12443_),
    .A1(\datamem.data_ram[28][22] ),
    .S(_12473_),
    .X(_12480_));
 sky130_fd_sc_hd__clkbuf_1 _28036_ (.A(_12480_),
    .X(_03845_));
 sky130_fd_sc_hd__mux2_1 _28037_ (.A0(_12445_),
    .A1(\datamem.data_ram[28][23] ),
    .S(_12473_),
    .X(_12481_));
 sky130_fd_sc_hd__clkbuf_1 _28038_ (.A(_12481_),
    .X(_03846_));
 sky130_fd_sc_hd__clkbuf_8 _28039_ (.A(_10500_),
    .X(_12482_));
 sky130_fd_sc_hd__a21oi_1 _28040_ (.A1(_09350_),
    .A2(_12345_),
    .B1(_12482_),
    .Y(_12483_));
 sky130_fd_sc_hd__mux2_1 _28041_ (.A0(_12447_),
    .A1(\datamem.data_ram[28][8] ),
    .S(net96),
    .X(_12484_));
 sky130_fd_sc_hd__clkbuf_1 _28042_ (.A(_12484_),
    .X(_03847_));
 sky130_fd_sc_hd__mux2_1 _28043_ (.A0(_12450_),
    .A1(\datamem.data_ram[28][9] ),
    .S(net96),
    .X(_12485_));
 sky130_fd_sc_hd__clkbuf_1 _28044_ (.A(_12485_),
    .X(_03848_));
 sky130_fd_sc_hd__mux2_1 _28045_ (.A0(_12452_),
    .A1(\datamem.data_ram[28][10] ),
    .S(net96),
    .X(_12486_));
 sky130_fd_sc_hd__clkbuf_1 _28046_ (.A(_12486_),
    .X(_03849_));
 sky130_fd_sc_hd__mux2_1 _28047_ (.A0(_12454_),
    .A1(\datamem.data_ram[28][11] ),
    .S(net96),
    .X(_12487_));
 sky130_fd_sc_hd__clkbuf_1 _28048_ (.A(_12487_),
    .X(_03850_));
 sky130_fd_sc_hd__mux2_1 _28049_ (.A0(_12456_),
    .A1(\datamem.data_ram[28][12] ),
    .S(net96),
    .X(_12488_));
 sky130_fd_sc_hd__clkbuf_1 _28050_ (.A(_12488_),
    .X(_03851_));
 sky130_fd_sc_hd__mux2_1 _28051_ (.A0(_12458_),
    .A1(\datamem.data_ram[28][13] ),
    .S(net96),
    .X(_12489_));
 sky130_fd_sc_hd__clkbuf_1 _28052_ (.A(_12489_),
    .X(_03852_));
 sky130_fd_sc_hd__mux2_1 _28053_ (.A0(_12460_),
    .A1(\datamem.data_ram[28][14] ),
    .S(net96),
    .X(_12490_));
 sky130_fd_sc_hd__clkbuf_1 _28054_ (.A(_12490_),
    .X(_03853_));
 sky130_fd_sc_hd__mux2_1 _28055_ (.A0(_12462_),
    .A1(\datamem.data_ram[28][15] ),
    .S(_12483_),
    .X(_12491_));
 sky130_fd_sc_hd__clkbuf_1 _28056_ (.A(_12491_),
    .X(_03854_));
 sky130_fd_sc_hd__a21oi_4 _28057_ (.A1(_10141_),
    .A2(_12325_),
    .B1(_12482_),
    .Y(_12492_));
 sky130_fd_sc_hd__mux2_1 _28058_ (.A0(_12355_),
    .A1(\datamem.data_ram[27][24] ),
    .S(_12492_),
    .X(_12493_));
 sky130_fd_sc_hd__clkbuf_1 _28059_ (.A(_12493_),
    .X(_03855_));
 sky130_fd_sc_hd__mux2_1 _28060_ (.A0(_12359_),
    .A1(\datamem.data_ram[27][25] ),
    .S(_12492_),
    .X(_12494_));
 sky130_fd_sc_hd__clkbuf_1 _28061_ (.A(_12494_),
    .X(_03856_));
 sky130_fd_sc_hd__mux2_1 _28062_ (.A0(_12361_),
    .A1(\datamem.data_ram[27][26] ),
    .S(_12492_),
    .X(_12495_));
 sky130_fd_sc_hd__clkbuf_1 _28063_ (.A(_12495_),
    .X(_03857_));
 sky130_fd_sc_hd__mux2_1 _28064_ (.A0(_12363_),
    .A1(\datamem.data_ram[27][27] ),
    .S(_12492_),
    .X(_12496_));
 sky130_fd_sc_hd__clkbuf_1 _28065_ (.A(_12496_),
    .X(_03858_));
 sky130_fd_sc_hd__mux2_1 _28066_ (.A0(_12365_),
    .A1(\datamem.data_ram[27][28] ),
    .S(_12492_),
    .X(_12497_));
 sky130_fd_sc_hd__clkbuf_1 _28067_ (.A(_12497_),
    .X(_03859_));
 sky130_fd_sc_hd__mux2_1 _28068_ (.A0(_12367_),
    .A1(\datamem.data_ram[27][29] ),
    .S(_12492_),
    .X(_12498_));
 sky130_fd_sc_hd__clkbuf_1 _28069_ (.A(_12498_),
    .X(_03860_));
 sky130_fd_sc_hd__mux2_1 _28070_ (.A0(_12369_),
    .A1(\datamem.data_ram[27][30] ),
    .S(_12492_),
    .X(_12499_));
 sky130_fd_sc_hd__clkbuf_1 _28071_ (.A(_12499_),
    .X(_03861_));
 sky130_fd_sc_hd__mux2_1 _28072_ (.A0(_12371_),
    .A1(\datamem.data_ram[27][31] ),
    .S(_12492_),
    .X(_12500_));
 sky130_fd_sc_hd__clkbuf_1 _28073_ (.A(_12500_),
    .X(_03862_));
 sky130_fd_sc_hd__a21oi_4 _28074_ (.A1(_10141_),
    .A2(_12335_),
    .B1(_12482_),
    .Y(_12501_));
 sky130_fd_sc_hd__mux2_1 _28075_ (.A0(_12430_),
    .A1(\datamem.data_ram[27][16] ),
    .S(_12501_),
    .X(_12502_));
 sky130_fd_sc_hd__clkbuf_1 _28076_ (.A(_12502_),
    .X(_03863_));
 sky130_fd_sc_hd__mux2_1 _28077_ (.A0(_12433_),
    .A1(\datamem.data_ram[27][17] ),
    .S(_12501_),
    .X(_12503_));
 sky130_fd_sc_hd__clkbuf_1 _28078_ (.A(_12503_),
    .X(_03864_));
 sky130_fd_sc_hd__mux2_1 _28079_ (.A0(_12435_),
    .A1(\datamem.data_ram[27][18] ),
    .S(_12501_),
    .X(_12504_));
 sky130_fd_sc_hd__clkbuf_1 _28080_ (.A(_12504_),
    .X(_03865_));
 sky130_fd_sc_hd__mux2_1 _28081_ (.A0(_12437_),
    .A1(\datamem.data_ram[27][19] ),
    .S(_12501_),
    .X(_12505_));
 sky130_fd_sc_hd__clkbuf_1 _28082_ (.A(_12505_),
    .X(_03866_));
 sky130_fd_sc_hd__mux2_1 _28083_ (.A0(_12439_),
    .A1(\datamem.data_ram[27][20] ),
    .S(_12501_),
    .X(_12506_));
 sky130_fd_sc_hd__clkbuf_1 _28084_ (.A(_12506_),
    .X(_03867_));
 sky130_fd_sc_hd__mux2_1 _28085_ (.A0(_12441_),
    .A1(\datamem.data_ram[27][21] ),
    .S(_12501_),
    .X(_12507_));
 sky130_fd_sc_hd__clkbuf_1 _28086_ (.A(_12507_),
    .X(_03868_));
 sky130_fd_sc_hd__mux2_1 _28087_ (.A0(_12443_),
    .A1(\datamem.data_ram[27][22] ),
    .S(_12501_),
    .X(_12508_));
 sky130_fd_sc_hd__clkbuf_1 _28088_ (.A(_12508_),
    .X(_03869_));
 sky130_fd_sc_hd__mux2_1 _28089_ (.A0(_12445_),
    .A1(\datamem.data_ram[27][23] ),
    .S(_12501_),
    .X(_12509_));
 sky130_fd_sc_hd__clkbuf_1 _28090_ (.A(_12509_),
    .X(_03870_));
 sky130_fd_sc_hd__a21oi_1 _28091_ (.A1(_10141_),
    .A2(_12345_),
    .B1(_12482_),
    .Y(_12510_));
 sky130_fd_sc_hd__mux2_1 _28092_ (.A0(_12447_),
    .A1(\datamem.data_ram[27][8] ),
    .S(net75),
    .X(_12511_));
 sky130_fd_sc_hd__clkbuf_1 _28093_ (.A(_12511_),
    .X(_03871_));
 sky130_fd_sc_hd__mux2_1 _28094_ (.A0(_12450_),
    .A1(\datamem.data_ram[27][9] ),
    .S(net75),
    .X(_12512_));
 sky130_fd_sc_hd__clkbuf_1 _28095_ (.A(_12512_),
    .X(_03872_));
 sky130_fd_sc_hd__mux2_1 _28096_ (.A0(_12452_),
    .A1(\datamem.data_ram[27][10] ),
    .S(net75),
    .X(_12513_));
 sky130_fd_sc_hd__clkbuf_1 _28097_ (.A(_12513_),
    .X(_03873_));
 sky130_fd_sc_hd__mux2_1 _28098_ (.A0(_12454_),
    .A1(\datamem.data_ram[27][11] ),
    .S(net75),
    .X(_12514_));
 sky130_fd_sc_hd__clkbuf_1 _28099_ (.A(_12514_),
    .X(_03874_));
 sky130_fd_sc_hd__mux2_1 _28100_ (.A0(_12456_),
    .A1(\datamem.data_ram[27][12] ),
    .S(net75),
    .X(_12515_));
 sky130_fd_sc_hd__clkbuf_1 _28101_ (.A(_12515_),
    .X(_03875_));
 sky130_fd_sc_hd__mux2_1 _28102_ (.A0(_12458_),
    .A1(\datamem.data_ram[27][13] ),
    .S(net75),
    .X(_12516_));
 sky130_fd_sc_hd__clkbuf_1 _28103_ (.A(_12516_),
    .X(_03876_));
 sky130_fd_sc_hd__mux2_1 _28104_ (.A0(_12460_),
    .A1(\datamem.data_ram[27][14] ),
    .S(net75),
    .X(_12517_));
 sky130_fd_sc_hd__clkbuf_1 _28105_ (.A(_12517_),
    .X(_03877_));
 sky130_fd_sc_hd__mux2_1 _28106_ (.A0(_12462_),
    .A1(\datamem.data_ram[27][15] ),
    .S(_12510_),
    .X(_12518_));
 sky130_fd_sc_hd__clkbuf_1 _28107_ (.A(_12518_),
    .X(_03878_));
 sky130_fd_sc_hd__a21oi_2 _28108_ (.A1(_10777_),
    .A2(_12325_),
    .B1(_12482_),
    .Y(_12519_));
 sky130_fd_sc_hd__mux2_1 _28109_ (.A0(_12355_),
    .A1(\datamem.data_ram[26][24] ),
    .S(net74),
    .X(_12520_));
 sky130_fd_sc_hd__clkbuf_1 _28110_ (.A(_12520_),
    .X(_03879_));
 sky130_fd_sc_hd__mux2_1 _28111_ (.A0(_12359_),
    .A1(\datamem.data_ram[26][25] ),
    .S(net74),
    .X(_12521_));
 sky130_fd_sc_hd__clkbuf_1 _28112_ (.A(_12521_),
    .X(_03880_));
 sky130_fd_sc_hd__mux2_1 _28113_ (.A0(_12361_),
    .A1(\datamem.data_ram[26][26] ),
    .S(net74),
    .X(_12522_));
 sky130_fd_sc_hd__clkbuf_1 _28114_ (.A(_12522_),
    .X(_03881_));
 sky130_fd_sc_hd__mux2_1 _28115_ (.A0(_12363_),
    .A1(\datamem.data_ram[26][27] ),
    .S(net74),
    .X(_12523_));
 sky130_fd_sc_hd__clkbuf_1 _28116_ (.A(_12523_),
    .X(_03882_));
 sky130_fd_sc_hd__mux2_1 _28117_ (.A0(_12365_),
    .A1(\datamem.data_ram[26][28] ),
    .S(net74),
    .X(_12524_));
 sky130_fd_sc_hd__clkbuf_1 _28118_ (.A(_12524_),
    .X(_03883_));
 sky130_fd_sc_hd__mux2_1 _28119_ (.A0(_12367_),
    .A1(\datamem.data_ram[26][29] ),
    .S(net74),
    .X(_12525_));
 sky130_fd_sc_hd__clkbuf_1 _28120_ (.A(_12525_),
    .X(_03884_));
 sky130_fd_sc_hd__mux2_1 _28121_ (.A0(_12369_),
    .A1(\datamem.data_ram[26][30] ),
    .S(_12519_),
    .X(_12526_));
 sky130_fd_sc_hd__clkbuf_1 _28122_ (.A(_12526_),
    .X(_03885_));
 sky130_fd_sc_hd__mux2_1 _28123_ (.A0(_12371_),
    .A1(\datamem.data_ram[26][31] ),
    .S(_12519_),
    .X(_12527_));
 sky130_fd_sc_hd__clkbuf_1 _28124_ (.A(_12527_),
    .X(_03886_));
 sky130_fd_sc_hd__a21oi_4 _28125_ (.A1(_10777_),
    .A2(_12335_),
    .B1(_12482_),
    .Y(_12528_));
 sky130_fd_sc_hd__mux2_1 _28126_ (.A0(_12430_),
    .A1(\datamem.data_ram[26][16] ),
    .S(_12528_),
    .X(_12529_));
 sky130_fd_sc_hd__clkbuf_1 _28127_ (.A(_12529_),
    .X(_03887_));
 sky130_fd_sc_hd__mux2_1 _28128_ (.A0(_12433_),
    .A1(\datamem.data_ram[26][17] ),
    .S(_12528_),
    .X(_12530_));
 sky130_fd_sc_hd__clkbuf_1 _28129_ (.A(_12530_),
    .X(_03888_));
 sky130_fd_sc_hd__mux2_1 _28130_ (.A0(_12435_),
    .A1(\datamem.data_ram[26][18] ),
    .S(_12528_),
    .X(_12531_));
 sky130_fd_sc_hd__clkbuf_1 _28131_ (.A(_12531_),
    .X(_03889_));
 sky130_fd_sc_hd__mux2_1 _28132_ (.A0(_12437_),
    .A1(\datamem.data_ram[26][19] ),
    .S(_12528_),
    .X(_12532_));
 sky130_fd_sc_hd__clkbuf_1 _28133_ (.A(_12532_),
    .X(_03890_));
 sky130_fd_sc_hd__mux2_1 _28134_ (.A0(_12439_),
    .A1(\datamem.data_ram[26][20] ),
    .S(_12528_),
    .X(_12533_));
 sky130_fd_sc_hd__clkbuf_1 _28135_ (.A(_12533_),
    .X(_03891_));
 sky130_fd_sc_hd__mux2_1 _28136_ (.A0(_12441_),
    .A1(\datamem.data_ram[26][21] ),
    .S(_12528_),
    .X(_12534_));
 sky130_fd_sc_hd__clkbuf_1 _28137_ (.A(_12534_),
    .X(_03892_));
 sky130_fd_sc_hd__mux2_1 _28138_ (.A0(_12443_),
    .A1(\datamem.data_ram[26][22] ),
    .S(_12528_),
    .X(_12535_));
 sky130_fd_sc_hd__clkbuf_1 _28139_ (.A(_12535_),
    .X(_03893_));
 sky130_fd_sc_hd__mux2_1 _28140_ (.A0(_12445_),
    .A1(\datamem.data_ram[26][23] ),
    .S(_12528_),
    .X(_12536_));
 sky130_fd_sc_hd__clkbuf_1 _28141_ (.A(_12536_),
    .X(_03894_));
 sky130_fd_sc_hd__a21oi_1 _28142_ (.A1(_10777_),
    .A2(_12345_),
    .B1(_12482_),
    .Y(_12537_));
 sky130_fd_sc_hd__mux2_1 _28143_ (.A0(_12447_),
    .A1(\datamem.data_ram[26][8] ),
    .S(net73),
    .X(_12538_));
 sky130_fd_sc_hd__clkbuf_1 _28144_ (.A(_12538_),
    .X(_03895_));
 sky130_fd_sc_hd__mux2_1 _28145_ (.A0(_12450_),
    .A1(\datamem.data_ram[26][9] ),
    .S(net73),
    .X(_12539_));
 sky130_fd_sc_hd__clkbuf_1 _28146_ (.A(_12539_),
    .X(_03896_));
 sky130_fd_sc_hd__mux2_1 _28147_ (.A0(_12452_),
    .A1(\datamem.data_ram[26][10] ),
    .S(net73),
    .X(_12540_));
 sky130_fd_sc_hd__clkbuf_1 _28148_ (.A(_12540_),
    .X(_03897_));
 sky130_fd_sc_hd__mux2_1 _28149_ (.A0(_12454_),
    .A1(\datamem.data_ram[26][11] ),
    .S(net73),
    .X(_12541_));
 sky130_fd_sc_hd__clkbuf_1 _28150_ (.A(_12541_),
    .X(_03898_));
 sky130_fd_sc_hd__mux2_1 _28151_ (.A0(_12456_),
    .A1(\datamem.data_ram[26][12] ),
    .S(net73),
    .X(_12542_));
 sky130_fd_sc_hd__clkbuf_1 _28152_ (.A(_12542_),
    .X(_03899_));
 sky130_fd_sc_hd__mux2_1 _28153_ (.A0(_12458_),
    .A1(\datamem.data_ram[26][13] ),
    .S(net73),
    .X(_12543_));
 sky130_fd_sc_hd__clkbuf_1 _28154_ (.A(_12543_),
    .X(_03900_));
 sky130_fd_sc_hd__mux2_1 _28155_ (.A0(_12460_),
    .A1(\datamem.data_ram[26][14] ),
    .S(net73),
    .X(_12544_));
 sky130_fd_sc_hd__clkbuf_1 _28156_ (.A(_12544_),
    .X(_03901_));
 sky130_fd_sc_hd__mux2_1 _28157_ (.A0(_12462_),
    .A1(\datamem.data_ram[26][15] ),
    .S(_12537_),
    .X(_12545_));
 sky130_fd_sc_hd__clkbuf_1 _28158_ (.A(_12545_),
    .X(_03902_));
 sky130_fd_sc_hd__a21oi_4 _28159_ (.A1(_12279_),
    .A2(_12325_),
    .B1(_12482_),
    .Y(_12546_));
 sky130_fd_sc_hd__mux2_1 _28160_ (.A0(_12355_),
    .A1(\datamem.data_ram[25][24] ),
    .S(_12546_),
    .X(_12547_));
 sky130_fd_sc_hd__clkbuf_1 _28161_ (.A(_12547_),
    .X(_03903_));
 sky130_fd_sc_hd__mux2_1 _28162_ (.A0(_12359_),
    .A1(\datamem.data_ram[25][25] ),
    .S(_12546_),
    .X(_12548_));
 sky130_fd_sc_hd__clkbuf_1 _28163_ (.A(_12548_),
    .X(_03904_));
 sky130_fd_sc_hd__mux2_1 _28164_ (.A0(_12361_),
    .A1(\datamem.data_ram[25][26] ),
    .S(_12546_),
    .X(_12549_));
 sky130_fd_sc_hd__clkbuf_1 _28165_ (.A(_12549_),
    .X(_03905_));
 sky130_fd_sc_hd__mux2_1 _28166_ (.A0(_12363_),
    .A1(\datamem.data_ram[25][27] ),
    .S(_12546_),
    .X(_12550_));
 sky130_fd_sc_hd__clkbuf_1 _28167_ (.A(_12550_),
    .X(_03906_));
 sky130_fd_sc_hd__mux2_1 _28168_ (.A0(_12365_),
    .A1(\datamem.data_ram[25][28] ),
    .S(_12546_),
    .X(_12551_));
 sky130_fd_sc_hd__clkbuf_1 _28169_ (.A(_12551_),
    .X(_03907_));
 sky130_fd_sc_hd__mux2_1 _28170_ (.A0(_12367_),
    .A1(\datamem.data_ram[25][29] ),
    .S(_12546_),
    .X(_12552_));
 sky130_fd_sc_hd__clkbuf_1 _28171_ (.A(_12552_),
    .X(_03908_));
 sky130_fd_sc_hd__mux2_1 _28172_ (.A0(_12369_),
    .A1(\datamem.data_ram[25][30] ),
    .S(_12546_),
    .X(_12553_));
 sky130_fd_sc_hd__clkbuf_1 _28173_ (.A(_12553_),
    .X(_03909_));
 sky130_fd_sc_hd__mux2_1 _28174_ (.A0(_12371_),
    .A1(\datamem.data_ram[25][31] ),
    .S(_12546_),
    .X(_12554_));
 sky130_fd_sc_hd__clkbuf_1 _28175_ (.A(_12554_),
    .X(_03910_));
 sky130_fd_sc_hd__a21oi_4 _28176_ (.A1(_12279_),
    .A2(_12335_),
    .B1(_12482_),
    .Y(_12555_));
 sky130_fd_sc_hd__mux2_1 _28177_ (.A0(_12430_),
    .A1(\datamem.data_ram[25][16] ),
    .S(_12555_),
    .X(_12556_));
 sky130_fd_sc_hd__clkbuf_1 _28178_ (.A(_12556_),
    .X(_03911_));
 sky130_fd_sc_hd__mux2_1 _28179_ (.A0(_12433_),
    .A1(\datamem.data_ram[25][17] ),
    .S(_12555_),
    .X(_12557_));
 sky130_fd_sc_hd__clkbuf_1 _28180_ (.A(_12557_),
    .X(_03912_));
 sky130_fd_sc_hd__mux2_1 _28181_ (.A0(_12435_),
    .A1(\datamem.data_ram[25][18] ),
    .S(_12555_),
    .X(_12558_));
 sky130_fd_sc_hd__clkbuf_1 _28182_ (.A(_12558_),
    .X(_03913_));
 sky130_fd_sc_hd__mux2_1 _28183_ (.A0(_12437_),
    .A1(\datamem.data_ram[25][19] ),
    .S(_12555_),
    .X(_12559_));
 sky130_fd_sc_hd__clkbuf_1 _28184_ (.A(_12559_),
    .X(_03914_));
 sky130_fd_sc_hd__mux2_1 _28185_ (.A0(_12439_),
    .A1(\datamem.data_ram[25][20] ),
    .S(_12555_),
    .X(_12560_));
 sky130_fd_sc_hd__clkbuf_1 _28186_ (.A(_12560_),
    .X(_03915_));
 sky130_fd_sc_hd__mux2_1 _28187_ (.A0(_12441_),
    .A1(\datamem.data_ram[25][21] ),
    .S(_12555_),
    .X(_12561_));
 sky130_fd_sc_hd__clkbuf_1 _28188_ (.A(_12561_),
    .X(_03916_));
 sky130_fd_sc_hd__mux2_1 _28189_ (.A0(_12443_),
    .A1(\datamem.data_ram[25][22] ),
    .S(_12555_),
    .X(_12562_));
 sky130_fd_sc_hd__clkbuf_1 _28190_ (.A(_12562_),
    .X(_03917_));
 sky130_fd_sc_hd__mux2_1 _28191_ (.A0(_12445_),
    .A1(\datamem.data_ram[25][23] ),
    .S(_12555_),
    .X(_12563_));
 sky130_fd_sc_hd__clkbuf_1 _28192_ (.A(_12563_),
    .X(_03918_));
 sky130_fd_sc_hd__a21oi_1 _28193_ (.A1(_12279_),
    .A2(_12345_),
    .B1(_12482_),
    .Y(_12564_));
 sky130_fd_sc_hd__mux2_1 _28194_ (.A0(_12447_),
    .A1(\datamem.data_ram[25][8] ),
    .S(net46),
    .X(_12565_));
 sky130_fd_sc_hd__clkbuf_1 _28195_ (.A(_12565_),
    .X(_03919_));
 sky130_fd_sc_hd__mux2_1 _28196_ (.A0(_12450_),
    .A1(\datamem.data_ram[25][9] ),
    .S(net46),
    .X(_12566_));
 sky130_fd_sc_hd__clkbuf_1 _28197_ (.A(_12566_),
    .X(_03920_));
 sky130_fd_sc_hd__mux2_1 _28198_ (.A0(_12452_),
    .A1(\datamem.data_ram[25][10] ),
    .S(net46),
    .X(_12567_));
 sky130_fd_sc_hd__clkbuf_1 _28199_ (.A(_12567_),
    .X(_03921_));
 sky130_fd_sc_hd__mux2_1 _28200_ (.A0(_12454_),
    .A1(\datamem.data_ram[25][11] ),
    .S(net46),
    .X(_12568_));
 sky130_fd_sc_hd__clkbuf_1 _28201_ (.A(_12568_),
    .X(_03922_));
 sky130_fd_sc_hd__mux2_1 _28202_ (.A0(_12456_),
    .A1(\datamem.data_ram[25][12] ),
    .S(net46),
    .X(_12569_));
 sky130_fd_sc_hd__clkbuf_1 _28203_ (.A(_12569_),
    .X(_03923_));
 sky130_fd_sc_hd__mux2_1 _28204_ (.A0(_12458_),
    .A1(\datamem.data_ram[25][13] ),
    .S(net46),
    .X(_12570_));
 sky130_fd_sc_hd__clkbuf_1 _28205_ (.A(_12570_),
    .X(_03924_));
 sky130_fd_sc_hd__mux2_1 _28206_ (.A0(_12460_),
    .A1(\datamem.data_ram[25][14] ),
    .S(net46),
    .X(_12571_));
 sky130_fd_sc_hd__clkbuf_1 _28207_ (.A(_12571_),
    .X(_03925_));
 sky130_fd_sc_hd__mux2_1 _28208_ (.A0(_12462_),
    .A1(\datamem.data_ram[25][15] ),
    .S(_12564_),
    .X(_12572_));
 sky130_fd_sc_hd__clkbuf_1 _28209_ (.A(_12572_),
    .X(_03926_));
 sky130_fd_sc_hd__buf_6 _28210_ (.A(_06591_),
    .X(_12573_));
 sky130_fd_sc_hd__a21oi_1 _28211_ (.A1(_10838_),
    .A2(_12325_),
    .B1(_12573_),
    .Y(_12574_));
 sky130_fd_sc_hd__mux2_1 _28212_ (.A0(_12355_),
    .A1(\datamem.data_ram[24][24] ),
    .S(net45),
    .X(_12575_));
 sky130_fd_sc_hd__clkbuf_1 _28213_ (.A(_12575_),
    .X(_03927_));
 sky130_fd_sc_hd__mux2_1 _28214_ (.A0(_12359_),
    .A1(\datamem.data_ram[24][25] ),
    .S(net45),
    .X(_12576_));
 sky130_fd_sc_hd__clkbuf_1 _28215_ (.A(_12576_),
    .X(_03928_));
 sky130_fd_sc_hd__mux2_1 _28216_ (.A0(_12361_),
    .A1(\datamem.data_ram[24][26] ),
    .S(net45),
    .X(_12577_));
 sky130_fd_sc_hd__clkbuf_1 _28217_ (.A(_12577_),
    .X(_03929_));
 sky130_fd_sc_hd__mux2_1 _28218_ (.A0(_12363_),
    .A1(\datamem.data_ram[24][27] ),
    .S(net45),
    .X(_12578_));
 sky130_fd_sc_hd__clkbuf_1 _28219_ (.A(_12578_),
    .X(_03930_));
 sky130_fd_sc_hd__mux2_1 _28220_ (.A0(_12365_),
    .A1(\datamem.data_ram[24][28] ),
    .S(net45),
    .X(_12579_));
 sky130_fd_sc_hd__clkbuf_1 _28221_ (.A(_12579_),
    .X(_03931_));
 sky130_fd_sc_hd__mux2_1 _28222_ (.A0(_12367_),
    .A1(\datamem.data_ram[24][29] ),
    .S(net45),
    .X(_12580_));
 sky130_fd_sc_hd__clkbuf_1 _28223_ (.A(_12580_),
    .X(_03932_));
 sky130_fd_sc_hd__mux2_1 _28224_ (.A0(_12369_),
    .A1(\datamem.data_ram[24][30] ),
    .S(net45),
    .X(_12581_));
 sky130_fd_sc_hd__clkbuf_1 _28225_ (.A(_12581_),
    .X(_03933_));
 sky130_fd_sc_hd__mux2_1 _28226_ (.A0(_12371_),
    .A1(\datamem.data_ram[24][31] ),
    .S(_12574_),
    .X(_12582_));
 sky130_fd_sc_hd__clkbuf_1 _28227_ (.A(_12582_),
    .X(_03934_));
 sky130_fd_sc_hd__a21oi_4 _28228_ (.A1(_10979_),
    .A2(_12335_),
    .B1(_12573_),
    .Y(_12583_));
 sky130_fd_sc_hd__mux2_1 _28229_ (.A0(_12430_),
    .A1(\datamem.data_ram[24][16] ),
    .S(_12583_),
    .X(_12584_));
 sky130_fd_sc_hd__clkbuf_1 _28230_ (.A(_12584_),
    .X(_03935_));
 sky130_fd_sc_hd__mux2_1 _28231_ (.A0(_12433_),
    .A1(\datamem.data_ram[24][17] ),
    .S(_12583_),
    .X(_12585_));
 sky130_fd_sc_hd__clkbuf_1 _28232_ (.A(_12585_),
    .X(_03936_));
 sky130_fd_sc_hd__mux2_1 _28233_ (.A0(_12435_),
    .A1(\datamem.data_ram[24][18] ),
    .S(_12583_),
    .X(_12586_));
 sky130_fd_sc_hd__clkbuf_1 _28234_ (.A(_12586_),
    .X(_03937_));
 sky130_fd_sc_hd__mux2_1 _28235_ (.A0(_12437_),
    .A1(\datamem.data_ram[24][19] ),
    .S(_12583_),
    .X(_12587_));
 sky130_fd_sc_hd__clkbuf_1 _28236_ (.A(_12587_),
    .X(_03938_));
 sky130_fd_sc_hd__mux2_1 _28237_ (.A0(_12439_),
    .A1(\datamem.data_ram[24][20] ),
    .S(_12583_),
    .X(_12588_));
 sky130_fd_sc_hd__clkbuf_1 _28238_ (.A(_12588_),
    .X(_03939_));
 sky130_fd_sc_hd__mux2_1 _28239_ (.A0(_12441_),
    .A1(\datamem.data_ram[24][21] ),
    .S(_12583_),
    .X(_12589_));
 sky130_fd_sc_hd__clkbuf_1 _28240_ (.A(_12589_),
    .X(_03940_));
 sky130_fd_sc_hd__mux2_1 _28241_ (.A0(_12443_),
    .A1(\datamem.data_ram[24][22] ),
    .S(_12583_),
    .X(_12590_));
 sky130_fd_sc_hd__clkbuf_1 _28242_ (.A(_12590_),
    .X(_03941_));
 sky130_fd_sc_hd__mux2_1 _28243_ (.A0(_12445_),
    .A1(\datamem.data_ram[24][23] ),
    .S(_12583_),
    .X(_12591_));
 sky130_fd_sc_hd__clkbuf_1 _28244_ (.A(_12591_),
    .X(_03942_));
 sky130_fd_sc_hd__a21oi_1 _28245_ (.A1(_10979_),
    .A2(_12345_),
    .B1(_12573_),
    .Y(_12592_));
 sky130_fd_sc_hd__mux2_1 _28246_ (.A0(_12447_),
    .A1(\datamem.data_ram[24][8] ),
    .S(net44),
    .X(_12593_));
 sky130_fd_sc_hd__clkbuf_1 _28247_ (.A(_12593_),
    .X(_03943_));
 sky130_fd_sc_hd__mux2_1 _28248_ (.A0(_12450_),
    .A1(\datamem.data_ram[24][9] ),
    .S(net44),
    .X(_12594_));
 sky130_fd_sc_hd__clkbuf_1 _28249_ (.A(_12594_),
    .X(_03944_));
 sky130_fd_sc_hd__mux2_1 _28250_ (.A0(_12452_),
    .A1(\datamem.data_ram[24][10] ),
    .S(net44),
    .X(_12595_));
 sky130_fd_sc_hd__clkbuf_1 _28251_ (.A(_12595_),
    .X(_03945_));
 sky130_fd_sc_hd__mux2_1 _28252_ (.A0(_12454_),
    .A1(\datamem.data_ram[24][11] ),
    .S(net44),
    .X(_12596_));
 sky130_fd_sc_hd__clkbuf_1 _28253_ (.A(_12596_),
    .X(_03946_));
 sky130_fd_sc_hd__mux2_1 _28254_ (.A0(_12456_),
    .A1(\datamem.data_ram[24][12] ),
    .S(net44),
    .X(_12597_));
 sky130_fd_sc_hd__clkbuf_1 _28255_ (.A(_12597_),
    .X(_03947_));
 sky130_fd_sc_hd__mux2_1 _28256_ (.A0(_12458_),
    .A1(\datamem.data_ram[24][13] ),
    .S(net44),
    .X(_12598_));
 sky130_fd_sc_hd__clkbuf_1 _28257_ (.A(_12598_),
    .X(_03948_));
 sky130_fd_sc_hd__mux2_1 _28258_ (.A0(_12460_),
    .A1(\datamem.data_ram[24][14] ),
    .S(net44),
    .X(_12599_));
 sky130_fd_sc_hd__clkbuf_1 _28259_ (.A(_12599_),
    .X(_03949_));
 sky130_fd_sc_hd__mux2_1 _28260_ (.A0(_12462_),
    .A1(\datamem.data_ram[24][15] ),
    .S(_12592_),
    .X(_12600_));
 sky130_fd_sc_hd__clkbuf_1 _28261_ (.A(_12600_),
    .X(_03950_));
 sky130_fd_sc_hd__clkbuf_16 _28262_ (.A(_07125_),
    .X(_12601_));
 sky130_fd_sc_hd__nor2_8 _28263_ (.A(_08133_),
    .B(net106),
    .Y(_12602_));
 sky130_fd_sc_hd__a21oi_4 _28264_ (.A1(_12601_),
    .A2(_12602_),
    .B1(_12573_),
    .Y(_12603_));
 sky130_fd_sc_hd__mux2_1 _28265_ (.A0(_12355_),
    .A1(\datamem.data_ram[23][24] ),
    .S(_12603_),
    .X(_12604_));
 sky130_fd_sc_hd__clkbuf_1 _28266_ (.A(_12604_),
    .X(_03951_));
 sky130_fd_sc_hd__mux2_1 _28267_ (.A0(_12359_),
    .A1(\datamem.data_ram[23][25] ),
    .S(_12603_),
    .X(_12605_));
 sky130_fd_sc_hd__clkbuf_1 _28268_ (.A(_12605_),
    .X(_03952_));
 sky130_fd_sc_hd__mux2_1 _28269_ (.A0(_12361_),
    .A1(\datamem.data_ram[23][26] ),
    .S(_12603_),
    .X(_12606_));
 sky130_fd_sc_hd__clkbuf_1 _28270_ (.A(_12606_),
    .X(_03953_));
 sky130_fd_sc_hd__mux2_1 _28271_ (.A0(_12363_),
    .A1(\datamem.data_ram[23][27] ),
    .S(_12603_),
    .X(_12607_));
 sky130_fd_sc_hd__clkbuf_1 _28272_ (.A(_12607_),
    .X(_03954_));
 sky130_fd_sc_hd__mux2_1 _28273_ (.A0(_12365_),
    .A1(\datamem.data_ram[23][28] ),
    .S(_12603_),
    .X(_12608_));
 sky130_fd_sc_hd__clkbuf_1 _28274_ (.A(_12608_),
    .X(_03955_));
 sky130_fd_sc_hd__mux2_1 _28275_ (.A0(_12367_),
    .A1(\datamem.data_ram[23][29] ),
    .S(_12603_),
    .X(_12609_));
 sky130_fd_sc_hd__clkbuf_1 _28276_ (.A(_12609_),
    .X(_03956_));
 sky130_fd_sc_hd__mux2_1 _28277_ (.A0(_12369_),
    .A1(\datamem.data_ram[23][30] ),
    .S(_12603_),
    .X(_12610_));
 sky130_fd_sc_hd__clkbuf_1 _28278_ (.A(_12610_),
    .X(_03957_));
 sky130_fd_sc_hd__mux2_1 _28279_ (.A0(_12371_),
    .A1(\datamem.data_ram[23][31] ),
    .S(_12603_),
    .X(_12611_));
 sky130_fd_sc_hd__clkbuf_1 _28280_ (.A(_12611_),
    .X(_03958_));
 sky130_fd_sc_hd__nor2_8 _28281_ (.A(_08133_),
    .B(_09228_),
    .Y(_12612_));
 sky130_fd_sc_hd__a21oi_4 _28282_ (.A1(_12601_),
    .A2(_12612_),
    .B1(_12573_),
    .Y(_12613_));
 sky130_fd_sc_hd__mux2_1 _28283_ (.A0(_12430_),
    .A1(\datamem.data_ram[23][16] ),
    .S(_12613_),
    .X(_12614_));
 sky130_fd_sc_hd__clkbuf_1 _28284_ (.A(_12614_),
    .X(_03959_));
 sky130_fd_sc_hd__mux2_1 _28285_ (.A0(_12433_),
    .A1(\datamem.data_ram[23][17] ),
    .S(_12613_),
    .X(_12615_));
 sky130_fd_sc_hd__clkbuf_1 _28286_ (.A(_12615_),
    .X(_03960_));
 sky130_fd_sc_hd__mux2_1 _28287_ (.A0(_12435_),
    .A1(\datamem.data_ram[23][18] ),
    .S(_12613_),
    .X(_12616_));
 sky130_fd_sc_hd__clkbuf_1 _28288_ (.A(_12616_),
    .X(_03961_));
 sky130_fd_sc_hd__mux2_1 _28289_ (.A0(_12437_),
    .A1(\datamem.data_ram[23][19] ),
    .S(_12613_),
    .X(_12617_));
 sky130_fd_sc_hd__clkbuf_1 _28290_ (.A(_12617_),
    .X(_03962_));
 sky130_fd_sc_hd__mux2_1 _28291_ (.A0(_12439_),
    .A1(\datamem.data_ram[23][20] ),
    .S(_12613_),
    .X(_12618_));
 sky130_fd_sc_hd__clkbuf_1 _28292_ (.A(_12618_),
    .X(_03963_));
 sky130_fd_sc_hd__mux2_1 _28293_ (.A0(_12441_),
    .A1(\datamem.data_ram[23][21] ),
    .S(_12613_),
    .X(_12619_));
 sky130_fd_sc_hd__clkbuf_1 _28294_ (.A(_12619_),
    .X(_03964_));
 sky130_fd_sc_hd__mux2_1 _28295_ (.A0(_12443_),
    .A1(\datamem.data_ram[23][22] ),
    .S(_12613_),
    .X(_12620_));
 sky130_fd_sc_hd__clkbuf_1 _28296_ (.A(_12620_),
    .X(_03965_));
 sky130_fd_sc_hd__mux2_1 _28297_ (.A0(_12445_),
    .A1(\datamem.data_ram[23][23] ),
    .S(_12613_),
    .X(_12621_));
 sky130_fd_sc_hd__clkbuf_1 _28298_ (.A(_12621_),
    .X(_03966_));
 sky130_fd_sc_hd__nor2_4 _28299_ (.A(_08133_),
    .B(_09268_),
    .Y(_12622_));
 sky130_fd_sc_hd__a21oi_1 _28300_ (.A1(_12601_),
    .A2(_12622_),
    .B1(_12573_),
    .Y(_12623_));
 sky130_fd_sc_hd__mux2_1 _28301_ (.A0(_12447_),
    .A1(\datamem.data_ram[23][8] ),
    .S(net72),
    .X(_12624_));
 sky130_fd_sc_hd__clkbuf_1 _28302_ (.A(_12624_),
    .X(_03967_));
 sky130_fd_sc_hd__mux2_1 _28303_ (.A0(_12450_),
    .A1(\datamem.data_ram[23][9] ),
    .S(net72),
    .X(_12625_));
 sky130_fd_sc_hd__clkbuf_1 _28304_ (.A(_12625_),
    .X(_03968_));
 sky130_fd_sc_hd__mux2_1 _28305_ (.A0(_12452_),
    .A1(\datamem.data_ram[23][10] ),
    .S(net72),
    .X(_12626_));
 sky130_fd_sc_hd__clkbuf_1 _28306_ (.A(_12626_),
    .X(_03969_));
 sky130_fd_sc_hd__mux2_1 _28307_ (.A0(_12454_),
    .A1(\datamem.data_ram[23][11] ),
    .S(net72),
    .X(_12627_));
 sky130_fd_sc_hd__clkbuf_1 _28308_ (.A(_12627_),
    .X(_03970_));
 sky130_fd_sc_hd__mux2_1 _28309_ (.A0(_12456_),
    .A1(\datamem.data_ram[23][12] ),
    .S(net72),
    .X(_12628_));
 sky130_fd_sc_hd__clkbuf_1 _28310_ (.A(_12628_),
    .X(_03971_));
 sky130_fd_sc_hd__mux2_1 _28311_ (.A0(_12458_),
    .A1(\datamem.data_ram[23][13] ),
    .S(_12623_),
    .X(_12629_));
 sky130_fd_sc_hd__clkbuf_1 _28312_ (.A(_12629_),
    .X(_03972_));
 sky130_fd_sc_hd__mux2_1 _28313_ (.A0(_12460_),
    .A1(\datamem.data_ram[23][14] ),
    .S(net72),
    .X(_12630_));
 sky130_fd_sc_hd__clkbuf_1 _28314_ (.A(_12630_),
    .X(_03973_));
 sky130_fd_sc_hd__mux2_1 _28315_ (.A0(_12462_),
    .A1(\datamem.data_ram[23][15] ),
    .S(net72),
    .X(_12631_));
 sky130_fd_sc_hd__clkbuf_1 _28316_ (.A(_12631_),
    .X(_03974_));
 sky130_fd_sc_hd__a21oi_4 _28317_ (.A1(_10668_),
    .A2(_12602_),
    .B1(_12573_),
    .Y(_12632_));
 sky130_fd_sc_hd__mux2_1 _28318_ (.A0(_12355_),
    .A1(\datamem.data_ram[22][24] ),
    .S(_12632_),
    .X(_12633_));
 sky130_fd_sc_hd__clkbuf_1 _28319_ (.A(_12633_),
    .X(_03975_));
 sky130_fd_sc_hd__mux2_1 _28320_ (.A0(_12359_),
    .A1(\datamem.data_ram[22][25] ),
    .S(_12632_),
    .X(_12634_));
 sky130_fd_sc_hd__clkbuf_1 _28321_ (.A(_12634_),
    .X(_03976_));
 sky130_fd_sc_hd__mux2_1 _28322_ (.A0(_12361_),
    .A1(\datamem.data_ram[22][26] ),
    .S(_12632_),
    .X(_12635_));
 sky130_fd_sc_hd__clkbuf_1 _28323_ (.A(_12635_),
    .X(_03977_));
 sky130_fd_sc_hd__mux2_1 _28324_ (.A0(_12363_),
    .A1(\datamem.data_ram[22][27] ),
    .S(_12632_),
    .X(_12636_));
 sky130_fd_sc_hd__clkbuf_1 _28325_ (.A(_12636_),
    .X(_03978_));
 sky130_fd_sc_hd__mux2_1 _28326_ (.A0(_12365_),
    .A1(\datamem.data_ram[22][28] ),
    .S(_12632_),
    .X(_12637_));
 sky130_fd_sc_hd__clkbuf_1 _28327_ (.A(_12637_),
    .X(_03979_));
 sky130_fd_sc_hd__mux2_1 _28328_ (.A0(_12367_),
    .A1(\datamem.data_ram[22][29] ),
    .S(_12632_),
    .X(_12638_));
 sky130_fd_sc_hd__clkbuf_1 _28329_ (.A(_12638_),
    .X(_03980_));
 sky130_fd_sc_hd__mux2_1 _28330_ (.A0(_12369_),
    .A1(\datamem.data_ram[22][30] ),
    .S(_12632_),
    .X(_12639_));
 sky130_fd_sc_hd__clkbuf_1 _28331_ (.A(_12639_),
    .X(_03981_));
 sky130_fd_sc_hd__mux2_1 _28332_ (.A0(_12371_),
    .A1(\datamem.data_ram[22][31] ),
    .S(_12632_),
    .X(_12640_));
 sky130_fd_sc_hd__clkbuf_1 _28333_ (.A(_12640_),
    .X(_03982_));
 sky130_fd_sc_hd__a21oi_4 _28334_ (.A1(_10668_),
    .A2(_12612_),
    .B1(_12573_),
    .Y(_12641_));
 sky130_fd_sc_hd__mux2_1 _28335_ (.A0(_12430_),
    .A1(\datamem.data_ram[22][16] ),
    .S(_12641_),
    .X(_12642_));
 sky130_fd_sc_hd__clkbuf_1 _28336_ (.A(_12642_),
    .X(_03983_));
 sky130_fd_sc_hd__mux2_1 _28337_ (.A0(_12433_),
    .A1(\datamem.data_ram[22][17] ),
    .S(_12641_),
    .X(_12643_));
 sky130_fd_sc_hd__clkbuf_1 _28338_ (.A(_12643_),
    .X(_03984_));
 sky130_fd_sc_hd__mux2_1 _28339_ (.A0(_12435_),
    .A1(\datamem.data_ram[22][18] ),
    .S(_12641_),
    .X(_12644_));
 sky130_fd_sc_hd__clkbuf_1 _28340_ (.A(_12644_),
    .X(_03985_));
 sky130_fd_sc_hd__mux2_1 _28341_ (.A0(_12437_),
    .A1(\datamem.data_ram[22][19] ),
    .S(_12641_),
    .X(_12645_));
 sky130_fd_sc_hd__clkbuf_1 _28342_ (.A(_12645_),
    .X(_03986_));
 sky130_fd_sc_hd__mux2_1 _28343_ (.A0(_12439_),
    .A1(\datamem.data_ram[22][20] ),
    .S(_12641_),
    .X(_12646_));
 sky130_fd_sc_hd__clkbuf_1 _28344_ (.A(_12646_),
    .X(_03987_));
 sky130_fd_sc_hd__mux2_1 _28345_ (.A0(_12441_),
    .A1(\datamem.data_ram[22][21] ),
    .S(_12641_),
    .X(_12647_));
 sky130_fd_sc_hd__clkbuf_1 _28346_ (.A(_12647_),
    .X(_03988_));
 sky130_fd_sc_hd__mux2_1 _28347_ (.A0(_12443_),
    .A1(\datamem.data_ram[22][22] ),
    .S(_12641_),
    .X(_12648_));
 sky130_fd_sc_hd__clkbuf_1 _28348_ (.A(_12648_),
    .X(_03989_));
 sky130_fd_sc_hd__mux2_1 _28349_ (.A0(_12445_),
    .A1(\datamem.data_ram[22][23] ),
    .S(_12641_),
    .X(_12649_));
 sky130_fd_sc_hd__clkbuf_1 _28350_ (.A(_12649_),
    .X(_03990_));
 sky130_fd_sc_hd__a21oi_1 _28351_ (.A1(_09225_),
    .A2(_12622_),
    .B1(_12573_),
    .Y(_12650_));
 sky130_fd_sc_hd__mux2_1 _28352_ (.A0(_12447_),
    .A1(\datamem.data_ram[22][8] ),
    .S(net95),
    .X(_12651_));
 sky130_fd_sc_hd__clkbuf_1 _28353_ (.A(_12651_),
    .X(_03991_));
 sky130_fd_sc_hd__mux2_1 _28354_ (.A0(_12450_),
    .A1(\datamem.data_ram[22][9] ),
    .S(net95),
    .X(_12652_));
 sky130_fd_sc_hd__clkbuf_1 _28355_ (.A(_12652_),
    .X(_03992_));
 sky130_fd_sc_hd__mux2_1 _28356_ (.A0(_12452_),
    .A1(\datamem.data_ram[22][10] ),
    .S(net95),
    .X(_12653_));
 sky130_fd_sc_hd__clkbuf_1 _28357_ (.A(_12653_),
    .X(_03993_));
 sky130_fd_sc_hd__mux2_1 _28358_ (.A0(_12454_),
    .A1(\datamem.data_ram[22][11] ),
    .S(net95),
    .X(_12654_));
 sky130_fd_sc_hd__clkbuf_1 _28359_ (.A(_12654_),
    .X(_03994_));
 sky130_fd_sc_hd__mux2_1 _28360_ (.A0(_12456_),
    .A1(\datamem.data_ram[22][12] ),
    .S(net95),
    .X(_12655_));
 sky130_fd_sc_hd__clkbuf_1 _28361_ (.A(_12655_),
    .X(_03995_));
 sky130_fd_sc_hd__mux2_1 _28362_ (.A0(_12458_),
    .A1(\datamem.data_ram[22][13] ),
    .S(_12650_),
    .X(_12656_));
 sky130_fd_sc_hd__clkbuf_1 _28363_ (.A(_12656_),
    .X(_03996_));
 sky130_fd_sc_hd__mux2_1 _28364_ (.A0(_12460_),
    .A1(\datamem.data_ram[22][14] ),
    .S(net95),
    .X(_12657_));
 sky130_fd_sc_hd__clkbuf_1 _28365_ (.A(_12657_),
    .X(_03997_));
 sky130_fd_sc_hd__mux2_1 _28366_ (.A0(_12462_),
    .A1(\datamem.data_ram[22][15] ),
    .S(net95),
    .X(_12658_));
 sky130_fd_sc_hd__clkbuf_1 _28367_ (.A(_12658_),
    .X(_03998_));
 sky130_fd_sc_hd__a21oi_4 _28368_ (.A1(_12178_),
    .A2(_12602_),
    .B1(_12573_),
    .Y(_12659_));
 sky130_fd_sc_hd__mux2_1 _28369_ (.A0(_12355_),
    .A1(\datamem.data_ram[21][24] ),
    .S(_12659_),
    .X(_12660_));
 sky130_fd_sc_hd__clkbuf_1 _28370_ (.A(_12660_),
    .X(_03999_));
 sky130_fd_sc_hd__mux2_1 _28371_ (.A0(_12359_),
    .A1(\datamem.data_ram[21][25] ),
    .S(_12659_),
    .X(_12661_));
 sky130_fd_sc_hd__clkbuf_1 _28372_ (.A(_12661_),
    .X(_04000_));
 sky130_fd_sc_hd__mux2_1 _28373_ (.A0(_12361_),
    .A1(\datamem.data_ram[21][26] ),
    .S(_12659_),
    .X(_12662_));
 sky130_fd_sc_hd__clkbuf_1 _28374_ (.A(_12662_),
    .X(_04001_));
 sky130_fd_sc_hd__mux2_1 _28375_ (.A0(_12363_),
    .A1(\datamem.data_ram[21][27] ),
    .S(_12659_),
    .X(_12663_));
 sky130_fd_sc_hd__clkbuf_1 _28376_ (.A(_12663_),
    .X(_04002_));
 sky130_fd_sc_hd__mux2_1 _28377_ (.A0(_12365_),
    .A1(\datamem.data_ram[21][28] ),
    .S(_12659_),
    .X(_12664_));
 sky130_fd_sc_hd__clkbuf_1 _28378_ (.A(_12664_),
    .X(_04003_));
 sky130_fd_sc_hd__mux2_1 _28379_ (.A0(_12367_),
    .A1(\datamem.data_ram[21][29] ),
    .S(_12659_),
    .X(_12665_));
 sky130_fd_sc_hd__clkbuf_1 _28380_ (.A(_12665_),
    .X(_04004_));
 sky130_fd_sc_hd__mux2_1 _28381_ (.A0(_12369_),
    .A1(\datamem.data_ram[21][30] ),
    .S(_12659_),
    .X(_12666_));
 sky130_fd_sc_hd__clkbuf_1 _28382_ (.A(_12666_),
    .X(_04005_));
 sky130_fd_sc_hd__mux2_1 _28383_ (.A0(_12371_),
    .A1(\datamem.data_ram[21][31] ),
    .S(_12659_),
    .X(_12667_));
 sky130_fd_sc_hd__clkbuf_1 _28384_ (.A(_12667_),
    .X(_04006_));
 sky130_fd_sc_hd__clkbuf_16 _28385_ (.A(_06591_),
    .X(_12668_));
 sky130_fd_sc_hd__a21oi_4 _28386_ (.A1(_12178_),
    .A2(_12612_),
    .B1(_12668_),
    .Y(_12669_));
 sky130_fd_sc_hd__mux2_1 _28387_ (.A0(_12430_),
    .A1(\datamem.data_ram[21][16] ),
    .S(_12669_),
    .X(_12670_));
 sky130_fd_sc_hd__clkbuf_1 _28388_ (.A(_12670_),
    .X(_04007_));
 sky130_fd_sc_hd__mux2_1 _28389_ (.A0(_12433_),
    .A1(\datamem.data_ram[21][17] ),
    .S(_12669_),
    .X(_12671_));
 sky130_fd_sc_hd__clkbuf_1 _28390_ (.A(_12671_),
    .X(_04008_));
 sky130_fd_sc_hd__mux2_1 _28391_ (.A0(_12435_),
    .A1(\datamem.data_ram[21][18] ),
    .S(_12669_),
    .X(_12672_));
 sky130_fd_sc_hd__clkbuf_1 _28392_ (.A(_12672_),
    .X(_04009_));
 sky130_fd_sc_hd__mux2_1 _28393_ (.A0(_12437_),
    .A1(\datamem.data_ram[21][19] ),
    .S(_12669_),
    .X(_12673_));
 sky130_fd_sc_hd__clkbuf_1 _28394_ (.A(_12673_),
    .X(_04010_));
 sky130_fd_sc_hd__mux2_1 _28395_ (.A0(_12439_),
    .A1(\datamem.data_ram[21][20] ),
    .S(_12669_),
    .X(_12674_));
 sky130_fd_sc_hd__clkbuf_1 _28396_ (.A(_12674_),
    .X(_04011_));
 sky130_fd_sc_hd__mux2_1 _28397_ (.A0(_12441_),
    .A1(\datamem.data_ram[21][21] ),
    .S(_12669_),
    .X(_12675_));
 sky130_fd_sc_hd__clkbuf_1 _28398_ (.A(_12675_),
    .X(_04012_));
 sky130_fd_sc_hd__mux2_1 _28399_ (.A0(_12443_),
    .A1(\datamem.data_ram[21][22] ),
    .S(_12669_),
    .X(_12676_));
 sky130_fd_sc_hd__clkbuf_1 _28400_ (.A(_12676_),
    .X(_04013_));
 sky130_fd_sc_hd__mux2_1 _28401_ (.A0(_12445_),
    .A1(\datamem.data_ram[21][23] ),
    .S(_12669_),
    .X(_12677_));
 sky130_fd_sc_hd__clkbuf_1 _28402_ (.A(_12677_),
    .X(_04014_));
 sky130_fd_sc_hd__a21oi_4 _28403_ (.A1(_12178_),
    .A2(_12622_),
    .B1(_12668_),
    .Y(_12678_));
 sky130_fd_sc_hd__mux2_1 _28404_ (.A0(_12447_),
    .A1(\datamem.data_ram[21][8] ),
    .S(_12678_),
    .X(_12679_));
 sky130_fd_sc_hd__clkbuf_1 _28405_ (.A(_12679_),
    .X(_04015_));
 sky130_fd_sc_hd__mux2_1 _28406_ (.A0(_12450_),
    .A1(\datamem.data_ram[21][9] ),
    .S(_12678_),
    .X(_12680_));
 sky130_fd_sc_hd__clkbuf_1 _28407_ (.A(_12680_),
    .X(_04016_));
 sky130_fd_sc_hd__mux2_1 _28408_ (.A0(_12452_),
    .A1(\datamem.data_ram[21][10] ),
    .S(_12678_),
    .X(_12681_));
 sky130_fd_sc_hd__clkbuf_1 _28409_ (.A(_12681_),
    .X(_04017_));
 sky130_fd_sc_hd__mux2_1 _28410_ (.A0(_12454_),
    .A1(\datamem.data_ram[21][11] ),
    .S(_12678_),
    .X(_12682_));
 sky130_fd_sc_hd__clkbuf_1 _28411_ (.A(_12682_),
    .X(_04018_));
 sky130_fd_sc_hd__mux2_1 _28412_ (.A0(_12456_),
    .A1(\datamem.data_ram[21][12] ),
    .S(_12678_),
    .X(_12683_));
 sky130_fd_sc_hd__clkbuf_1 _28413_ (.A(_12683_),
    .X(_04019_));
 sky130_fd_sc_hd__mux2_1 _28414_ (.A0(_12458_),
    .A1(\datamem.data_ram[21][13] ),
    .S(_12678_),
    .X(_12684_));
 sky130_fd_sc_hd__clkbuf_1 _28415_ (.A(_12684_),
    .X(_04020_));
 sky130_fd_sc_hd__mux2_1 _28416_ (.A0(_12460_),
    .A1(\datamem.data_ram[21][14] ),
    .S(_12678_),
    .X(_12685_));
 sky130_fd_sc_hd__clkbuf_1 _28417_ (.A(_12685_),
    .X(_04021_));
 sky130_fd_sc_hd__mux2_1 _28418_ (.A0(_12462_),
    .A1(\datamem.data_ram[21][15] ),
    .S(_12678_),
    .X(_12686_));
 sky130_fd_sc_hd__clkbuf_1 _28419_ (.A(_12686_),
    .X(_04022_));
 sky130_fd_sc_hd__clkbuf_2 _28420_ (.A(_09297_),
    .X(_12687_));
 sky130_fd_sc_hd__a21oi_4 _28421_ (.A1(_09350_),
    .A2(_12602_),
    .B1(_12668_),
    .Y(_12688_));
 sky130_fd_sc_hd__mux2_1 _28422_ (.A0(_12687_),
    .A1(\datamem.data_ram[20][24] ),
    .S(_12688_),
    .X(_12689_));
 sky130_fd_sc_hd__clkbuf_1 _28423_ (.A(_12689_),
    .X(_04023_));
 sky130_fd_sc_hd__clkbuf_2 _28424_ (.A(_09305_),
    .X(_12690_));
 sky130_fd_sc_hd__mux2_1 _28425_ (.A0(_12690_),
    .A1(\datamem.data_ram[20][25] ),
    .S(_12688_),
    .X(_12691_));
 sky130_fd_sc_hd__clkbuf_1 _28426_ (.A(_12691_),
    .X(_04024_));
 sky130_fd_sc_hd__clkbuf_2 _28427_ (.A(_09309_),
    .X(_12692_));
 sky130_fd_sc_hd__mux2_1 _28428_ (.A0(_12692_),
    .A1(\datamem.data_ram[20][26] ),
    .S(_12688_),
    .X(_12693_));
 sky130_fd_sc_hd__clkbuf_1 _28429_ (.A(_12693_),
    .X(_04025_));
 sky130_fd_sc_hd__clkbuf_2 _28430_ (.A(_09313_),
    .X(_12694_));
 sky130_fd_sc_hd__mux2_1 _28431_ (.A0(_12694_),
    .A1(\datamem.data_ram[20][27] ),
    .S(_12688_),
    .X(_12695_));
 sky130_fd_sc_hd__clkbuf_1 _28432_ (.A(_12695_),
    .X(_04026_));
 sky130_fd_sc_hd__clkbuf_2 _28433_ (.A(_09317_),
    .X(_12696_));
 sky130_fd_sc_hd__mux2_1 _28434_ (.A0(_12696_),
    .A1(\datamem.data_ram[20][28] ),
    .S(_12688_),
    .X(_12697_));
 sky130_fd_sc_hd__clkbuf_1 _28435_ (.A(_12697_),
    .X(_04027_));
 sky130_fd_sc_hd__clkbuf_2 _28436_ (.A(_09321_),
    .X(_12698_));
 sky130_fd_sc_hd__mux2_1 _28437_ (.A0(_12698_),
    .A1(\datamem.data_ram[20][29] ),
    .S(_12688_),
    .X(_12699_));
 sky130_fd_sc_hd__clkbuf_1 _28438_ (.A(_12699_),
    .X(_04028_));
 sky130_fd_sc_hd__clkbuf_2 _28439_ (.A(_09325_),
    .X(_12700_));
 sky130_fd_sc_hd__mux2_1 _28440_ (.A0(_12700_),
    .A1(\datamem.data_ram[20][30] ),
    .S(_12688_),
    .X(_12701_));
 sky130_fd_sc_hd__clkbuf_1 _28441_ (.A(_12701_),
    .X(_04029_));
 sky130_fd_sc_hd__clkbuf_2 _28442_ (.A(_09329_),
    .X(_12702_));
 sky130_fd_sc_hd__mux2_1 _28443_ (.A0(_12702_),
    .A1(\datamem.data_ram[20][31] ),
    .S(_12688_),
    .X(_12703_));
 sky130_fd_sc_hd__clkbuf_1 _28444_ (.A(_12703_),
    .X(_04030_));
 sky130_fd_sc_hd__a21oi_4 _28445_ (.A1(_09350_),
    .A2(_12612_),
    .B1(_12668_),
    .Y(_12704_));
 sky130_fd_sc_hd__mux2_1 _28446_ (.A0(_12430_),
    .A1(\datamem.data_ram[20][16] ),
    .S(_12704_),
    .X(_12705_));
 sky130_fd_sc_hd__clkbuf_1 _28447_ (.A(_12705_),
    .X(_04031_));
 sky130_fd_sc_hd__mux2_1 _28448_ (.A0(_12433_),
    .A1(\datamem.data_ram[20][17] ),
    .S(_12704_),
    .X(_12706_));
 sky130_fd_sc_hd__clkbuf_1 _28449_ (.A(_12706_),
    .X(_04032_));
 sky130_fd_sc_hd__mux2_1 _28450_ (.A0(_12435_),
    .A1(\datamem.data_ram[20][18] ),
    .S(_12704_),
    .X(_12707_));
 sky130_fd_sc_hd__clkbuf_1 _28451_ (.A(_12707_),
    .X(_04033_));
 sky130_fd_sc_hd__mux2_1 _28452_ (.A0(_12437_),
    .A1(\datamem.data_ram[20][19] ),
    .S(_12704_),
    .X(_12708_));
 sky130_fd_sc_hd__clkbuf_1 _28453_ (.A(_12708_),
    .X(_04034_));
 sky130_fd_sc_hd__mux2_1 _28454_ (.A0(_12439_),
    .A1(\datamem.data_ram[20][20] ),
    .S(_12704_),
    .X(_12709_));
 sky130_fd_sc_hd__clkbuf_1 _28455_ (.A(_12709_),
    .X(_04035_));
 sky130_fd_sc_hd__mux2_1 _28456_ (.A0(_12441_),
    .A1(\datamem.data_ram[20][21] ),
    .S(_12704_),
    .X(_12710_));
 sky130_fd_sc_hd__clkbuf_1 _28457_ (.A(_12710_),
    .X(_04036_));
 sky130_fd_sc_hd__mux2_1 _28458_ (.A0(_12443_),
    .A1(\datamem.data_ram[20][22] ),
    .S(_12704_),
    .X(_12711_));
 sky130_fd_sc_hd__clkbuf_1 _28459_ (.A(_12711_),
    .X(_04037_));
 sky130_fd_sc_hd__mux2_1 _28460_ (.A0(_12445_),
    .A1(\datamem.data_ram[20][23] ),
    .S(_12704_),
    .X(_12712_));
 sky130_fd_sc_hd__clkbuf_1 _28461_ (.A(_12712_),
    .X(_04038_));
 sky130_fd_sc_hd__a21oi_4 _28462_ (.A1(_09350_),
    .A2(_12622_),
    .B1(_12668_),
    .Y(_12713_));
 sky130_fd_sc_hd__mux2_1 _28463_ (.A0(_12447_),
    .A1(\datamem.data_ram[20][8] ),
    .S(_12713_),
    .X(_12714_));
 sky130_fd_sc_hd__clkbuf_1 _28464_ (.A(_12714_),
    .X(_04039_));
 sky130_fd_sc_hd__mux2_1 _28465_ (.A0(_12450_),
    .A1(\datamem.data_ram[20][9] ),
    .S(_12713_),
    .X(_12715_));
 sky130_fd_sc_hd__clkbuf_1 _28466_ (.A(_12715_),
    .X(_04040_));
 sky130_fd_sc_hd__mux2_1 _28467_ (.A0(_12452_),
    .A1(\datamem.data_ram[20][10] ),
    .S(_12713_),
    .X(_12716_));
 sky130_fd_sc_hd__clkbuf_1 _28468_ (.A(_12716_),
    .X(_04041_));
 sky130_fd_sc_hd__mux2_1 _28469_ (.A0(_12454_),
    .A1(\datamem.data_ram[20][11] ),
    .S(_12713_),
    .X(_12717_));
 sky130_fd_sc_hd__clkbuf_1 _28470_ (.A(_12717_),
    .X(_04042_));
 sky130_fd_sc_hd__mux2_1 _28471_ (.A0(_12456_),
    .A1(\datamem.data_ram[20][12] ),
    .S(_12713_),
    .X(_12718_));
 sky130_fd_sc_hd__clkbuf_1 _28472_ (.A(_12718_),
    .X(_04043_));
 sky130_fd_sc_hd__mux2_1 _28473_ (.A0(_12458_),
    .A1(\datamem.data_ram[20][13] ),
    .S(_12713_),
    .X(_12719_));
 sky130_fd_sc_hd__clkbuf_1 _28474_ (.A(_12719_),
    .X(_04044_));
 sky130_fd_sc_hd__mux2_1 _28475_ (.A0(_12460_),
    .A1(\datamem.data_ram[20][14] ),
    .S(_12713_),
    .X(_12720_));
 sky130_fd_sc_hd__clkbuf_1 _28476_ (.A(_12720_),
    .X(_04045_));
 sky130_fd_sc_hd__mux2_1 _28477_ (.A0(_12462_),
    .A1(\datamem.data_ram[20][15] ),
    .S(_12713_),
    .X(_12721_));
 sky130_fd_sc_hd__clkbuf_1 _28478_ (.A(_12721_),
    .X(_04046_));
 sky130_fd_sc_hd__or3_1 _28479_ (.A(_07808_),
    .B(_10042_),
    .C(_10044_),
    .X(_12722_));
 sky130_fd_sc_hd__buf_2 _28480_ (.A(_12722_),
    .X(_12723_));
 sky130_fd_sc_hd__and3_2 _28481_ (.A(_06997_),
    .B(_10049_),
    .C(_10921_),
    .X(_12724_));
 sky130_fd_sc_hd__and2_1 _28482_ (.A(_11965_),
    .B(_12724_),
    .X(_12725_));
 sky130_fd_sc_hd__a31o_1 _28483_ (.A1(_12391_),
    .A2(\datamem.data_ram[1][0] ),
    .A3(_12723_),
    .B1(_12725_),
    .X(_04047_));
 sky130_fd_sc_hd__and2_1 _28484_ (.A(_11968_),
    .B(_12724_),
    .X(_12726_));
 sky130_fd_sc_hd__a31o_1 _28485_ (.A1(_12391_),
    .A2(\datamem.data_ram[1][1] ),
    .A3(_12723_),
    .B1(_12726_),
    .X(_04048_));
 sky130_fd_sc_hd__buf_2 _28486_ (.A(_06587_),
    .X(_12727_));
 sky130_fd_sc_hd__and2_1 _28487_ (.A(_11970_),
    .B(_12724_),
    .X(_12728_));
 sky130_fd_sc_hd__a31o_1 _28488_ (.A1(_12727_),
    .A2(\datamem.data_ram[1][2] ),
    .A3(_12723_),
    .B1(_12728_),
    .X(_04049_));
 sky130_fd_sc_hd__and2_1 _28489_ (.A(_11972_),
    .B(_12724_),
    .X(_12729_));
 sky130_fd_sc_hd__a31o_1 _28490_ (.A1(_12727_),
    .A2(\datamem.data_ram[1][3] ),
    .A3(_12723_),
    .B1(_12729_),
    .X(_04050_));
 sky130_fd_sc_hd__or3_1 _28491_ (.A(_09231_),
    .B(\datamem.data_ram[1][4] ),
    .C(_12724_),
    .X(_12730_));
 sky130_fd_sc_hd__o21a_1 _28492_ (.A1(_10782_),
    .A2(_12723_),
    .B1(_12730_),
    .X(_04051_));
 sky130_fd_sc_hd__and2_1 _28493_ (.A(_11976_),
    .B(_12724_),
    .X(_12731_));
 sky130_fd_sc_hd__a31o_1 _28494_ (.A1(_12727_),
    .A2(\datamem.data_ram[1][5] ),
    .A3(_12723_),
    .B1(_12731_),
    .X(_04052_));
 sky130_fd_sc_hd__and2_1 _28495_ (.A(_11978_),
    .B(_12724_),
    .X(_12732_));
 sky130_fd_sc_hd__a31o_1 _28496_ (.A1(_12727_),
    .A2(\datamem.data_ram[1][6] ),
    .A3(_12723_),
    .B1(_12732_),
    .X(_04053_));
 sky130_fd_sc_hd__and2_1 _28497_ (.A(_11980_),
    .B(_12724_),
    .X(_12733_));
 sky130_fd_sc_hd__a31o_1 _28498_ (.A1(_12727_),
    .A2(\datamem.data_ram[1][7] ),
    .A3(_12723_),
    .B1(_12733_),
    .X(_04054_));
 sky130_fd_sc_hd__clkbuf_2 _28499_ (.A(_09266_),
    .X(_12734_));
 sky130_fd_sc_hd__a21oi_4 _28500_ (.A1(_12279_),
    .A2(_10092_),
    .B1(_12668_),
    .Y(_12735_));
 sky130_fd_sc_hd__mux2_1 _28501_ (.A0(_12734_),
    .A1(\datamem.data_ram[1][8] ),
    .S(net43),
    .X(_12736_));
 sky130_fd_sc_hd__clkbuf_1 _28502_ (.A(_12736_),
    .X(_04055_));
 sky130_fd_sc_hd__clkbuf_2 _28503_ (.A(_09272_),
    .X(_12737_));
 sky130_fd_sc_hd__mux2_1 _28504_ (.A0(_12737_),
    .A1(\datamem.data_ram[1][9] ),
    .S(net43),
    .X(_12738_));
 sky130_fd_sc_hd__clkbuf_1 _28505_ (.A(_12738_),
    .X(_04056_));
 sky130_fd_sc_hd__clkbuf_2 _28506_ (.A(_09275_),
    .X(_12739_));
 sky130_fd_sc_hd__mux2_1 _28507_ (.A0(_12739_),
    .A1(\datamem.data_ram[1][10] ),
    .S(net43),
    .X(_12740_));
 sky130_fd_sc_hd__clkbuf_1 _28508_ (.A(_12740_),
    .X(_04057_));
 sky130_fd_sc_hd__clkbuf_2 _28509_ (.A(_09278_),
    .X(_12741_));
 sky130_fd_sc_hd__mux2_1 _28510_ (.A0(_12741_),
    .A1(\datamem.data_ram[1][11] ),
    .S(net43),
    .X(_12742_));
 sky130_fd_sc_hd__clkbuf_1 _28511_ (.A(_12742_),
    .X(_04058_));
 sky130_fd_sc_hd__clkbuf_2 _28512_ (.A(_09281_),
    .X(_12743_));
 sky130_fd_sc_hd__mux2_1 _28513_ (.A0(_12743_),
    .A1(\datamem.data_ram[1][12] ),
    .S(net43),
    .X(_12744_));
 sky130_fd_sc_hd__clkbuf_1 _28514_ (.A(_12744_),
    .X(_04059_));
 sky130_fd_sc_hd__clkbuf_2 _28515_ (.A(_09284_),
    .X(_12745_));
 sky130_fd_sc_hd__mux2_1 _28516_ (.A0(_12745_),
    .A1(\datamem.data_ram[1][13] ),
    .S(_12735_),
    .X(_12746_));
 sky130_fd_sc_hd__clkbuf_1 _28517_ (.A(_12746_),
    .X(_04060_));
 sky130_fd_sc_hd__clkbuf_2 _28518_ (.A(_09287_),
    .X(_12747_));
 sky130_fd_sc_hd__mux2_1 _28519_ (.A0(_12747_),
    .A1(\datamem.data_ram[1][14] ),
    .S(_12735_),
    .X(_12748_));
 sky130_fd_sc_hd__clkbuf_1 _28520_ (.A(_12748_),
    .X(_04061_));
 sky130_fd_sc_hd__clkbuf_2 _28521_ (.A(_09290_),
    .X(_12749_));
 sky130_fd_sc_hd__mux2_1 _28522_ (.A0(_12749_),
    .A1(\datamem.data_ram[1][15] ),
    .S(_12735_),
    .X(_12750_));
 sky130_fd_sc_hd__clkbuf_1 _28523_ (.A(_12750_),
    .X(_04062_));
 sky130_fd_sc_hd__buf_2 _28524_ (.A(_09223_),
    .X(_12751_));
 sky130_fd_sc_hd__a21oi_4 _28525_ (.A1(_12279_),
    .A2(_10114_),
    .B1(_12668_),
    .Y(_12752_));
 sky130_fd_sc_hd__mux2_1 _28526_ (.A0(_12751_),
    .A1(\datamem.data_ram[1][16] ),
    .S(_12752_),
    .X(_12753_));
 sky130_fd_sc_hd__clkbuf_1 _28527_ (.A(_12753_),
    .X(_04063_));
 sky130_fd_sc_hd__buf_2 _28528_ (.A(_09235_),
    .X(_12754_));
 sky130_fd_sc_hd__mux2_1 _28529_ (.A0(_12754_),
    .A1(\datamem.data_ram[1][17] ),
    .S(_12752_),
    .X(_12755_));
 sky130_fd_sc_hd__clkbuf_1 _28530_ (.A(_12755_),
    .X(_04064_));
 sky130_fd_sc_hd__buf_2 _28531_ (.A(_09239_),
    .X(_12756_));
 sky130_fd_sc_hd__mux2_1 _28532_ (.A0(_12756_),
    .A1(\datamem.data_ram[1][18] ),
    .S(_12752_),
    .X(_12757_));
 sky130_fd_sc_hd__clkbuf_1 _28533_ (.A(_12757_),
    .X(_04065_));
 sky130_fd_sc_hd__buf_2 _28534_ (.A(_09243_),
    .X(_12758_));
 sky130_fd_sc_hd__mux2_1 _28535_ (.A0(_12758_),
    .A1(\datamem.data_ram[1][19] ),
    .S(_12752_),
    .X(_12759_));
 sky130_fd_sc_hd__clkbuf_1 _28536_ (.A(_12759_),
    .X(_04066_));
 sky130_fd_sc_hd__buf_2 _28537_ (.A(_09247_),
    .X(_12760_));
 sky130_fd_sc_hd__mux2_1 _28538_ (.A0(_12760_),
    .A1(\datamem.data_ram[1][20] ),
    .S(_12752_),
    .X(_12761_));
 sky130_fd_sc_hd__clkbuf_1 _28539_ (.A(_12761_),
    .X(_04067_));
 sky130_fd_sc_hd__buf_2 _28540_ (.A(_09251_),
    .X(_12762_));
 sky130_fd_sc_hd__mux2_1 _28541_ (.A0(_12762_),
    .A1(\datamem.data_ram[1][21] ),
    .S(_12752_),
    .X(_12763_));
 sky130_fd_sc_hd__clkbuf_1 _28542_ (.A(_12763_),
    .X(_04068_));
 sky130_fd_sc_hd__buf_2 _28543_ (.A(_09255_),
    .X(_12764_));
 sky130_fd_sc_hd__mux2_1 _28544_ (.A0(_12764_),
    .A1(\datamem.data_ram[1][22] ),
    .S(_12752_),
    .X(_12765_));
 sky130_fd_sc_hd__clkbuf_1 _28545_ (.A(_12765_),
    .X(_04069_));
 sky130_fd_sc_hd__buf_2 _28546_ (.A(_09259_),
    .X(_12766_));
 sky130_fd_sc_hd__mux2_1 _28547_ (.A0(_12766_),
    .A1(\datamem.data_ram[1][23] ),
    .S(_12752_),
    .X(_12767_));
 sky130_fd_sc_hd__clkbuf_1 _28548_ (.A(_12767_),
    .X(_04070_));
 sky130_fd_sc_hd__a21oi_4 _28549_ (.A1(_10141_),
    .A2(_12602_),
    .B1(_12668_),
    .Y(_12768_));
 sky130_fd_sc_hd__mux2_1 _28550_ (.A0(_12687_),
    .A1(\datamem.data_ram[19][24] ),
    .S(_12768_),
    .X(_12769_));
 sky130_fd_sc_hd__clkbuf_1 _28551_ (.A(_12769_),
    .X(_04071_));
 sky130_fd_sc_hd__mux2_1 _28552_ (.A0(_12690_),
    .A1(\datamem.data_ram[19][25] ),
    .S(_12768_),
    .X(_12770_));
 sky130_fd_sc_hd__clkbuf_1 _28553_ (.A(_12770_),
    .X(_04072_));
 sky130_fd_sc_hd__mux2_1 _28554_ (.A0(_12692_),
    .A1(\datamem.data_ram[19][26] ),
    .S(_12768_),
    .X(_12771_));
 sky130_fd_sc_hd__clkbuf_1 _28555_ (.A(_12771_),
    .X(_04073_));
 sky130_fd_sc_hd__mux2_1 _28556_ (.A0(_12694_),
    .A1(\datamem.data_ram[19][27] ),
    .S(_12768_),
    .X(_12772_));
 sky130_fd_sc_hd__clkbuf_1 _28557_ (.A(_12772_),
    .X(_04074_));
 sky130_fd_sc_hd__mux2_1 _28558_ (.A0(_12696_),
    .A1(\datamem.data_ram[19][28] ),
    .S(_12768_),
    .X(_12773_));
 sky130_fd_sc_hd__clkbuf_1 _28559_ (.A(_12773_),
    .X(_04075_));
 sky130_fd_sc_hd__mux2_1 _28560_ (.A0(_12698_),
    .A1(\datamem.data_ram[19][29] ),
    .S(_12768_),
    .X(_12774_));
 sky130_fd_sc_hd__clkbuf_1 _28561_ (.A(_12774_),
    .X(_04076_));
 sky130_fd_sc_hd__mux2_1 _28562_ (.A0(_12700_),
    .A1(\datamem.data_ram[19][30] ),
    .S(_12768_),
    .X(_12775_));
 sky130_fd_sc_hd__clkbuf_1 _28563_ (.A(_12775_),
    .X(_04077_));
 sky130_fd_sc_hd__mux2_1 _28564_ (.A0(_12702_),
    .A1(\datamem.data_ram[19][31] ),
    .S(_12768_),
    .X(_12776_));
 sky130_fd_sc_hd__clkbuf_1 _28565_ (.A(_12776_),
    .X(_04078_));
 sky130_fd_sc_hd__a21oi_4 _28566_ (.A1(_10141_),
    .A2(_12612_),
    .B1(_12668_),
    .Y(_12777_));
 sky130_fd_sc_hd__mux2_1 _28567_ (.A0(_12751_),
    .A1(\datamem.data_ram[19][16] ),
    .S(_12777_),
    .X(_12778_));
 sky130_fd_sc_hd__clkbuf_1 _28568_ (.A(_12778_),
    .X(_04079_));
 sky130_fd_sc_hd__mux2_1 _28569_ (.A0(_12754_),
    .A1(\datamem.data_ram[19][17] ),
    .S(_12777_),
    .X(_12779_));
 sky130_fd_sc_hd__clkbuf_1 _28570_ (.A(_12779_),
    .X(_04080_));
 sky130_fd_sc_hd__mux2_1 _28571_ (.A0(_12756_),
    .A1(\datamem.data_ram[19][18] ),
    .S(_12777_),
    .X(_12780_));
 sky130_fd_sc_hd__clkbuf_1 _28572_ (.A(_12780_),
    .X(_04081_));
 sky130_fd_sc_hd__mux2_1 _28573_ (.A0(_12758_),
    .A1(\datamem.data_ram[19][19] ),
    .S(_12777_),
    .X(_12781_));
 sky130_fd_sc_hd__clkbuf_1 _28574_ (.A(_12781_),
    .X(_04082_));
 sky130_fd_sc_hd__mux2_1 _28575_ (.A0(_12760_),
    .A1(\datamem.data_ram[19][20] ),
    .S(_12777_),
    .X(_12782_));
 sky130_fd_sc_hd__clkbuf_1 _28576_ (.A(_12782_),
    .X(_04083_));
 sky130_fd_sc_hd__mux2_1 _28577_ (.A0(_12762_),
    .A1(\datamem.data_ram[19][21] ),
    .S(_12777_),
    .X(_12783_));
 sky130_fd_sc_hd__clkbuf_1 _28578_ (.A(_12783_),
    .X(_04084_));
 sky130_fd_sc_hd__mux2_1 _28579_ (.A0(_12764_),
    .A1(\datamem.data_ram[19][22] ),
    .S(_12777_),
    .X(_12784_));
 sky130_fd_sc_hd__clkbuf_1 _28580_ (.A(_12784_),
    .X(_04085_));
 sky130_fd_sc_hd__mux2_1 _28581_ (.A0(_12766_),
    .A1(\datamem.data_ram[19][23] ),
    .S(_12777_),
    .X(_12785_));
 sky130_fd_sc_hd__clkbuf_1 _28582_ (.A(_12785_),
    .X(_04086_));
 sky130_fd_sc_hd__a21oi_4 _28583_ (.A1(_10141_),
    .A2(_12622_),
    .B1(_12668_),
    .Y(_12786_));
 sky130_fd_sc_hd__mux2_1 _28584_ (.A0(_12734_),
    .A1(\datamem.data_ram[19][8] ),
    .S(_12786_),
    .X(_12787_));
 sky130_fd_sc_hd__clkbuf_1 _28585_ (.A(_12787_),
    .X(_04087_));
 sky130_fd_sc_hd__mux2_1 _28586_ (.A0(_12737_),
    .A1(\datamem.data_ram[19][9] ),
    .S(_12786_),
    .X(_12788_));
 sky130_fd_sc_hd__clkbuf_1 _28587_ (.A(_12788_),
    .X(_04088_));
 sky130_fd_sc_hd__mux2_1 _28588_ (.A0(_12739_),
    .A1(\datamem.data_ram[19][10] ),
    .S(_12786_),
    .X(_12789_));
 sky130_fd_sc_hd__clkbuf_1 _28589_ (.A(_12789_),
    .X(_04089_));
 sky130_fd_sc_hd__mux2_1 _28590_ (.A0(_12741_),
    .A1(\datamem.data_ram[19][11] ),
    .S(_12786_),
    .X(_12790_));
 sky130_fd_sc_hd__clkbuf_1 _28591_ (.A(_12790_),
    .X(_04090_));
 sky130_fd_sc_hd__mux2_1 _28592_ (.A0(_12743_),
    .A1(\datamem.data_ram[19][12] ),
    .S(_12786_),
    .X(_12791_));
 sky130_fd_sc_hd__clkbuf_1 _28593_ (.A(_12791_),
    .X(_04091_));
 sky130_fd_sc_hd__mux2_1 _28594_ (.A0(_12745_),
    .A1(\datamem.data_ram[19][13] ),
    .S(_12786_),
    .X(_12792_));
 sky130_fd_sc_hd__clkbuf_1 _28595_ (.A(_12792_),
    .X(_04092_));
 sky130_fd_sc_hd__mux2_1 _28596_ (.A0(_12747_),
    .A1(\datamem.data_ram[19][14] ),
    .S(_12786_),
    .X(_12793_));
 sky130_fd_sc_hd__clkbuf_1 _28597_ (.A(_12793_),
    .X(_04093_));
 sky130_fd_sc_hd__mux2_1 _28598_ (.A0(_12749_),
    .A1(\datamem.data_ram[19][15] ),
    .S(_12786_),
    .X(_12794_));
 sky130_fd_sc_hd__clkbuf_1 _28599_ (.A(_12794_),
    .X(_04094_));
 sky130_fd_sc_hd__buf_8 _28600_ (.A(_06591_),
    .X(_12795_));
 sky130_fd_sc_hd__a21oi_4 _28601_ (.A1(_10777_),
    .A2(_12602_),
    .B1(_12795_),
    .Y(_12796_));
 sky130_fd_sc_hd__mux2_1 _28602_ (.A0(_12687_),
    .A1(\datamem.data_ram[18][24] ),
    .S(_12796_),
    .X(_12797_));
 sky130_fd_sc_hd__clkbuf_1 _28603_ (.A(_12797_),
    .X(_04095_));
 sky130_fd_sc_hd__mux2_1 _28604_ (.A0(_12690_),
    .A1(\datamem.data_ram[18][25] ),
    .S(_12796_),
    .X(_12798_));
 sky130_fd_sc_hd__clkbuf_1 _28605_ (.A(_12798_),
    .X(_04096_));
 sky130_fd_sc_hd__mux2_1 _28606_ (.A0(_12692_),
    .A1(\datamem.data_ram[18][26] ),
    .S(_12796_),
    .X(_12799_));
 sky130_fd_sc_hd__clkbuf_1 _28607_ (.A(_12799_),
    .X(_04097_));
 sky130_fd_sc_hd__mux2_1 _28608_ (.A0(_12694_),
    .A1(\datamem.data_ram[18][27] ),
    .S(_12796_),
    .X(_12800_));
 sky130_fd_sc_hd__clkbuf_1 _28609_ (.A(_12800_),
    .X(_04098_));
 sky130_fd_sc_hd__mux2_1 _28610_ (.A0(_12696_),
    .A1(\datamem.data_ram[18][28] ),
    .S(_12796_),
    .X(_12801_));
 sky130_fd_sc_hd__clkbuf_1 _28611_ (.A(_12801_),
    .X(_04099_));
 sky130_fd_sc_hd__mux2_1 _28612_ (.A0(_12698_),
    .A1(\datamem.data_ram[18][29] ),
    .S(_12796_),
    .X(_12802_));
 sky130_fd_sc_hd__clkbuf_1 _28613_ (.A(_12802_),
    .X(_04100_));
 sky130_fd_sc_hd__mux2_1 _28614_ (.A0(_12700_),
    .A1(\datamem.data_ram[18][30] ),
    .S(_12796_),
    .X(_12803_));
 sky130_fd_sc_hd__clkbuf_1 _28615_ (.A(_12803_),
    .X(_04101_));
 sky130_fd_sc_hd__mux2_1 _28616_ (.A0(_12702_),
    .A1(\datamem.data_ram[18][31] ),
    .S(_12796_),
    .X(_12804_));
 sky130_fd_sc_hd__clkbuf_1 _28617_ (.A(_12804_),
    .X(_04102_));
 sky130_fd_sc_hd__a21oi_4 _28618_ (.A1(_10777_),
    .A2(_12612_),
    .B1(_12795_),
    .Y(_12805_));
 sky130_fd_sc_hd__mux2_1 _28619_ (.A0(_12751_),
    .A1(\datamem.data_ram[18][16] ),
    .S(_12805_),
    .X(_12806_));
 sky130_fd_sc_hd__clkbuf_1 _28620_ (.A(_12806_),
    .X(_04103_));
 sky130_fd_sc_hd__mux2_1 _28621_ (.A0(_12754_),
    .A1(\datamem.data_ram[18][17] ),
    .S(_12805_),
    .X(_12807_));
 sky130_fd_sc_hd__clkbuf_1 _28622_ (.A(_12807_),
    .X(_04104_));
 sky130_fd_sc_hd__mux2_1 _28623_ (.A0(_12756_),
    .A1(\datamem.data_ram[18][18] ),
    .S(_12805_),
    .X(_12808_));
 sky130_fd_sc_hd__clkbuf_1 _28624_ (.A(_12808_),
    .X(_04105_));
 sky130_fd_sc_hd__mux2_1 _28625_ (.A0(_12758_),
    .A1(\datamem.data_ram[18][19] ),
    .S(_12805_),
    .X(_12809_));
 sky130_fd_sc_hd__clkbuf_1 _28626_ (.A(_12809_),
    .X(_04106_));
 sky130_fd_sc_hd__mux2_1 _28627_ (.A0(_12760_),
    .A1(\datamem.data_ram[18][20] ),
    .S(_12805_),
    .X(_12810_));
 sky130_fd_sc_hd__clkbuf_1 _28628_ (.A(_12810_),
    .X(_04107_));
 sky130_fd_sc_hd__mux2_1 _28629_ (.A0(_12762_),
    .A1(\datamem.data_ram[18][21] ),
    .S(_12805_),
    .X(_12811_));
 sky130_fd_sc_hd__clkbuf_1 _28630_ (.A(_12811_),
    .X(_04108_));
 sky130_fd_sc_hd__mux2_1 _28631_ (.A0(_12764_),
    .A1(\datamem.data_ram[18][22] ),
    .S(_12805_),
    .X(_12812_));
 sky130_fd_sc_hd__clkbuf_1 _28632_ (.A(_12812_),
    .X(_04109_));
 sky130_fd_sc_hd__mux2_1 _28633_ (.A0(_12766_),
    .A1(\datamem.data_ram[18][23] ),
    .S(_12805_),
    .X(_12813_));
 sky130_fd_sc_hd__clkbuf_1 _28634_ (.A(_12813_),
    .X(_04110_));
 sky130_fd_sc_hd__a21oi_2 _28635_ (.A1(_10777_),
    .A2(_12622_),
    .B1(_12795_),
    .Y(_12814_));
 sky130_fd_sc_hd__mux2_1 _28636_ (.A0(_12734_),
    .A1(\datamem.data_ram[18][8] ),
    .S(net71),
    .X(_12815_));
 sky130_fd_sc_hd__clkbuf_1 _28637_ (.A(_12815_),
    .X(_04111_));
 sky130_fd_sc_hd__mux2_1 _28638_ (.A0(_12737_),
    .A1(\datamem.data_ram[18][9] ),
    .S(net71),
    .X(_12816_));
 sky130_fd_sc_hd__clkbuf_1 _28639_ (.A(_12816_),
    .X(_04112_));
 sky130_fd_sc_hd__mux2_1 _28640_ (.A0(_12739_),
    .A1(\datamem.data_ram[18][10] ),
    .S(net71),
    .X(_12817_));
 sky130_fd_sc_hd__clkbuf_1 _28641_ (.A(_12817_),
    .X(_04113_));
 sky130_fd_sc_hd__mux2_1 _28642_ (.A0(_12741_),
    .A1(\datamem.data_ram[18][11] ),
    .S(net71),
    .X(_12818_));
 sky130_fd_sc_hd__clkbuf_1 _28643_ (.A(_12818_),
    .X(_04114_));
 sky130_fd_sc_hd__mux2_1 _28644_ (.A0(_12743_),
    .A1(\datamem.data_ram[18][12] ),
    .S(net71),
    .X(_12819_));
 sky130_fd_sc_hd__clkbuf_1 _28645_ (.A(_12819_),
    .X(_04115_));
 sky130_fd_sc_hd__mux2_1 _28646_ (.A0(_12745_),
    .A1(\datamem.data_ram[18][13] ),
    .S(_12814_),
    .X(_12820_));
 sky130_fd_sc_hd__clkbuf_1 _28647_ (.A(_12820_),
    .X(_04116_));
 sky130_fd_sc_hd__mux2_1 _28648_ (.A0(_12747_),
    .A1(\datamem.data_ram[18][14] ),
    .S(net71),
    .X(_12821_));
 sky130_fd_sc_hd__clkbuf_1 _28649_ (.A(_12821_),
    .X(_04117_));
 sky130_fd_sc_hd__mux2_1 _28650_ (.A0(_12749_),
    .A1(\datamem.data_ram[18][15] ),
    .S(_12814_),
    .X(_12822_));
 sky130_fd_sc_hd__clkbuf_1 _28651_ (.A(_12822_),
    .X(_04118_));
 sky130_fd_sc_hd__a21oi_4 _28652_ (.A1(_12279_),
    .A2(_12602_),
    .B1(_12795_),
    .Y(_12823_));
 sky130_fd_sc_hd__mux2_1 _28653_ (.A0(_12687_),
    .A1(\datamem.data_ram[17][24] ),
    .S(_12823_),
    .X(_12824_));
 sky130_fd_sc_hd__clkbuf_1 _28654_ (.A(_12824_),
    .X(_04119_));
 sky130_fd_sc_hd__mux2_1 _28655_ (.A0(_12690_),
    .A1(\datamem.data_ram[17][25] ),
    .S(_12823_),
    .X(_12825_));
 sky130_fd_sc_hd__clkbuf_1 _28656_ (.A(_12825_),
    .X(_04120_));
 sky130_fd_sc_hd__mux2_1 _28657_ (.A0(_12692_),
    .A1(\datamem.data_ram[17][26] ),
    .S(_12823_),
    .X(_12826_));
 sky130_fd_sc_hd__clkbuf_1 _28658_ (.A(_12826_),
    .X(_04121_));
 sky130_fd_sc_hd__mux2_1 _28659_ (.A0(_12694_),
    .A1(\datamem.data_ram[17][27] ),
    .S(_12823_),
    .X(_12827_));
 sky130_fd_sc_hd__clkbuf_1 _28660_ (.A(_12827_),
    .X(_04122_));
 sky130_fd_sc_hd__mux2_1 _28661_ (.A0(_12696_),
    .A1(\datamem.data_ram[17][28] ),
    .S(_12823_),
    .X(_12828_));
 sky130_fd_sc_hd__clkbuf_1 _28662_ (.A(_12828_),
    .X(_04123_));
 sky130_fd_sc_hd__mux2_1 _28663_ (.A0(_12698_),
    .A1(\datamem.data_ram[17][29] ),
    .S(_12823_),
    .X(_12829_));
 sky130_fd_sc_hd__clkbuf_1 _28664_ (.A(_12829_),
    .X(_04124_));
 sky130_fd_sc_hd__mux2_1 _28665_ (.A0(_12700_),
    .A1(\datamem.data_ram[17][30] ),
    .S(_12823_),
    .X(_12830_));
 sky130_fd_sc_hd__clkbuf_1 _28666_ (.A(_12830_),
    .X(_04125_));
 sky130_fd_sc_hd__mux2_1 _28667_ (.A0(_12702_),
    .A1(\datamem.data_ram[17][31] ),
    .S(_12823_),
    .X(_12831_));
 sky130_fd_sc_hd__clkbuf_1 _28668_ (.A(_12831_),
    .X(_04126_));
 sky130_fd_sc_hd__a21oi_4 _28669_ (.A1(_12279_),
    .A2(_12612_),
    .B1(_12795_),
    .Y(_12832_));
 sky130_fd_sc_hd__mux2_1 _28670_ (.A0(_12751_),
    .A1(\datamem.data_ram[17][16] ),
    .S(_12832_),
    .X(_12833_));
 sky130_fd_sc_hd__clkbuf_1 _28671_ (.A(_12833_),
    .X(_04127_));
 sky130_fd_sc_hd__mux2_1 _28672_ (.A0(_12754_),
    .A1(\datamem.data_ram[17][17] ),
    .S(_12832_),
    .X(_12834_));
 sky130_fd_sc_hd__clkbuf_1 _28673_ (.A(_12834_),
    .X(_04128_));
 sky130_fd_sc_hd__mux2_1 _28674_ (.A0(_12756_),
    .A1(\datamem.data_ram[17][18] ),
    .S(_12832_),
    .X(_12835_));
 sky130_fd_sc_hd__clkbuf_1 _28675_ (.A(_12835_),
    .X(_04129_));
 sky130_fd_sc_hd__mux2_1 _28676_ (.A0(_12758_),
    .A1(\datamem.data_ram[17][19] ),
    .S(_12832_),
    .X(_12836_));
 sky130_fd_sc_hd__clkbuf_1 _28677_ (.A(_12836_),
    .X(_04130_));
 sky130_fd_sc_hd__mux2_1 _28678_ (.A0(_12760_),
    .A1(\datamem.data_ram[17][20] ),
    .S(_12832_),
    .X(_12837_));
 sky130_fd_sc_hd__clkbuf_1 _28679_ (.A(_12837_),
    .X(_04131_));
 sky130_fd_sc_hd__mux2_1 _28680_ (.A0(_12762_),
    .A1(\datamem.data_ram[17][21] ),
    .S(_12832_),
    .X(_12838_));
 sky130_fd_sc_hd__clkbuf_1 _28681_ (.A(_12838_),
    .X(_04132_));
 sky130_fd_sc_hd__mux2_1 _28682_ (.A0(_12764_),
    .A1(\datamem.data_ram[17][22] ),
    .S(_12832_),
    .X(_12839_));
 sky130_fd_sc_hd__clkbuf_1 _28683_ (.A(_12839_),
    .X(_04133_));
 sky130_fd_sc_hd__mux2_1 _28684_ (.A0(_12766_),
    .A1(\datamem.data_ram[17][23] ),
    .S(_12832_),
    .X(_12840_));
 sky130_fd_sc_hd__clkbuf_1 _28685_ (.A(_12840_),
    .X(_04134_));
 sky130_fd_sc_hd__a21oi_1 _28686_ (.A1(_12279_),
    .A2(_12622_),
    .B1(_12795_),
    .Y(_12841_));
 sky130_fd_sc_hd__mux2_1 _28687_ (.A0(_12734_),
    .A1(\datamem.data_ram[17][8] ),
    .S(net42),
    .X(_12842_));
 sky130_fd_sc_hd__clkbuf_1 _28688_ (.A(_12842_),
    .X(_04135_));
 sky130_fd_sc_hd__mux2_1 _28689_ (.A0(_12737_),
    .A1(\datamem.data_ram[17][9] ),
    .S(net42),
    .X(_12843_));
 sky130_fd_sc_hd__clkbuf_1 _28690_ (.A(_12843_),
    .X(_04136_));
 sky130_fd_sc_hd__mux2_1 _28691_ (.A0(_12739_),
    .A1(\datamem.data_ram[17][10] ),
    .S(net42),
    .X(_12844_));
 sky130_fd_sc_hd__clkbuf_1 _28692_ (.A(_12844_),
    .X(_04137_));
 sky130_fd_sc_hd__mux2_1 _28693_ (.A0(_12741_),
    .A1(\datamem.data_ram[17][11] ),
    .S(net42),
    .X(_12845_));
 sky130_fd_sc_hd__clkbuf_1 _28694_ (.A(_12845_),
    .X(_04138_));
 sky130_fd_sc_hd__mux2_1 _28695_ (.A0(_12743_),
    .A1(\datamem.data_ram[17][12] ),
    .S(net42),
    .X(_12846_));
 sky130_fd_sc_hd__clkbuf_1 _28696_ (.A(_12846_),
    .X(_04139_));
 sky130_fd_sc_hd__mux2_1 _28697_ (.A0(_12745_),
    .A1(\datamem.data_ram[17][13] ),
    .S(net42),
    .X(_12847_));
 sky130_fd_sc_hd__clkbuf_1 _28698_ (.A(_12847_),
    .X(_04140_));
 sky130_fd_sc_hd__mux2_1 _28699_ (.A0(_12747_),
    .A1(\datamem.data_ram[17][14] ),
    .S(net42),
    .X(_12848_));
 sky130_fd_sc_hd__clkbuf_1 _28700_ (.A(_12848_),
    .X(_04141_));
 sky130_fd_sc_hd__mux2_1 _28701_ (.A0(_12749_),
    .A1(\datamem.data_ram[17][15] ),
    .S(net42),
    .X(_12849_));
 sky130_fd_sc_hd__clkbuf_1 _28702_ (.A(_12849_),
    .X(_04142_));
 sky130_fd_sc_hd__a21oi_4 _28703_ (.A1(_10979_),
    .A2(_12602_),
    .B1(_12795_),
    .Y(_12850_));
 sky130_fd_sc_hd__mux2_1 _28704_ (.A0(_12687_),
    .A1(\datamem.data_ram[16][24] ),
    .S(_12850_),
    .X(_12851_));
 sky130_fd_sc_hd__clkbuf_1 _28705_ (.A(_12851_),
    .X(_04143_));
 sky130_fd_sc_hd__mux2_1 _28706_ (.A0(_12690_),
    .A1(\datamem.data_ram[16][25] ),
    .S(_12850_),
    .X(_12852_));
 sky130_fd_sc_hd__clkbuf_1 _28707_ (.A(_12852_),
    .X(_04144_));
 sky130_fd_sc_hd__mux2_1 _28708_ (.A0(_12692_),
    .A1(\datamem.data_ram[16][26] ),
    .S(_12850_),
    .X(_12853_));
 sky130_fd_sc_hd__clkbuf_1 _28709_ (.A(_12853_),
    .X(_04145_));
 sky130_fd_sc_hd__mux2_1 _28710_ (.A0(_12694_),
    .A1(\datamem.data_ram[16][27] ),
    .S(_12850_),
    .X(_12854_));
 sky130_fd_sc_hd__clkbuf_1 _28711_ (.A(_12854_),
    .X(_04146_));
 sky130_fd_sc_hd__mux2_1 _28712_ (.A0(_12696_),
    .A1(\datamem.data_ram[16][28] ),
    .S(_12850_),
    .X(_12855_));
 sky130_fd_sc_hd__clkbuf_1 _28713_ (.A(_12855_),
    .X(_04147_));
 sky130_fd_sc_hd__mux2_1 _28714_ (.A0(_12698_),
    .A1(\datamem.data_ram[16][29] ),
    .S(_12850_),
    .X(_12856_));
 sky130_fd_sc_hd__clkbuf_1 _28715_ (.A(_12856_),
    .X(_04148_));
 sky130_fd_sc_hd__mux2_1 _28716_ (.A0(_12700_),
    .A1(\datamem.data_ram[16][30] ),
    .S(_12850_),
    .X(_12857_));
 sky130_fd_sc_hd__clkbuf_1 _28717_ (.A(_12857_),
    .X(_04149_));
 sky130_fd_sc_hd__mux2_1 _28718_ (.A0(_12702_),
    .A1(\datamem.data_ram[16][31] ),
    .S(_12850_),
    .X(_12858_));
 sky130_fd_sc_hd__clkbuf_1 _28719_ (.A(_12858_),
    .X(_04150_));
 sky130_fd_sc_hd__a21oi_4 _28720_ (.A1(_10979_),
    .A2(_12612_),
    .B1(_12795_),
    .Y(_12859_));
 sky130_fd_sc_hd__mux2_1 _28721_ (.A0(_12751_),
    .A1(\datamem.data_ram[16][16] ),
    .S(_12859_),
    .X(_12860_));
 sky130_fd_sc_hd__clkbuf_1 _28722_ (.A(_12860_),
    .X(_04151_));
 sky130_fd_sc_hd__mux2_1 _28723_ (.A0(_12754_),
    .A1(\datamem.data_ram[16][17] ),
    .S(_12859_),
    .X(_12861_));
 sky130_fd_sc_hd__clkbuf_1 _28724_ (.A(_12861_),
    .X(_04152_));
 sky130_fd_sc_hd__mux2_1 _28725_ (.A0(_12756_),
    .A1(\datamem.data_ram[16][18] ),
    .S(_12859_),
    .X(_12862_));
 sky130_fd_sc_hd__clkbuf_1 _28726_ (.A(_12862_),
    .X(_04153_));
 sky130_fd_sc_hd__mux2_1 _28727_ (.A0(_12758_),
    .A1(\datamem.data_ram[16][19] ),
    .S(_12859_),
    .X(_12863_));
 sky130_fd_sc_hd__clkbuf_1 _28728_ (.A(_12863_),
    .X(_04154_));
 sky130_fd_sc_hd__mux2_1 _28729_ (.A0(_12760_),
    .A1(\datamem.data_ram[16][20] ),
    .S(_12859_),
    .X(_12864_));
 sky130_fd_sc_hd__clkbuf_1 _28730_ (.A(_12864_),
    .X(_04155_));
 sky130_fd_sc_hd__mux2_1 _28731_ (.A0(_12762_),
    .A1(\datamem.data_ram[16][21] ),
    .S(_12859_),
    .X(_12865_));
 sky130_fd_sc_hd__clkbuf_1 _28732_ (.A(_12865_),
    .X(_04156_));
 sky130_fd_sc_hd__mux2_1 _28733_ (.A0(_12764_),
    .A1(\datamem.data_ram[16][22] ),
    .S(_12859_),
    .X(_12866_));
 sky130_fd_sc_hd__clkbuf_1 _28734_ (.A(_12866_),
    .X(_04157_));
 sky130_fd_sc_hd__mux2_1 _28735_ (.A0(_12766_),
    .A1(\datamem.data_ram[16][23] ),
    .S(_12859_),
    .X(_12867_));
 sky130_fd_sc_hd__clkbuf_1 _28736_ (.A(_12867_),
    .X(_04158_));
 sky130_fd_sc_hd__a21oi_1 _28737_ (.A1(_10979_),
    .A2(_12622_),
    .B1(_12795_),
    .Y(_12868_));
 sky130_fd_sc_hd__mux2_1 _28738_ (.A0(_12734_),
    .A1(\datamem.data_ram[16][8] ),
    .S(net41),
    .X(_12869_));
 sky130_fd_sc_hd__clkbuf_1 _28739_ (.A(_12869_),
    .X(_04159_));
 sky130_fd_sc_hd__mux2_1 _28740_ (.A0(_12737_),
    .A1(\datamem.data_ram[16][9] ),
    .S(net41),
    .X(_12870_));
 sky130_fd_sc_hd__clkbuf_1 _28741_ (.A(_12870_),
    .X(_04160_));
 sky130_fd_sc_hd__mux2_1 _28742_ (.A0(_12739_),
    .A1(\datamem.data_ram[16][10] ),
    .S(net41),
    .X(_12871_));
 sky130_fd_sc_hd__clkbuf_1 _28743_ (.A(_12871_),
    .X(_04161_));
 sky130_fd_sc_hd__mux2_1 _28744_ (.A0(_12741_),
    .A1(\datamem.data_ram[16][11] ),
    .S(net41),
    .X(_12872_));
 sky130_fd_sc_hd__clkbuf_1 _28745_ (.A(_12872_),
    .X(_04162_));
 sky130_fd_sc_hd__mux2_1 _28746_ (.A0(_12743_),
    .A1(\datamem.data_ram[16][12] ),
    .S(net41),
    .X(_12873_));
 sky130_fd_sc_hd__clkbuf_1 _28747_ (.A(_12873_),
    .X(_04163_));
 sky130_fd_sc_hd__mux2_1 _28748_ (.A0(_12745_),
    .A1(\datamem.data_ram[16][13] ),
    .S(net41),
    .X(_12874_));
 sky130_fd_sc_hd__clkbuf_1 _28749_ (.A(_12874_),
    .X(_04164_));
 sky130_fd_sc_hd__mux2_1 _28750_ (.A0(_12747_),
    .A1(\datamem.data_ram[16][14] ),
    .S(net41),
    .X(_12875_));
 sky130_fd_sc_hd__clkbuf_1 _28751_ (.A(_12875_),
    .X(_04165_));
 sky130_fd_sc_hd__mux2_1 _28752_ (.A0(_12749_),
    .A1(\datamem.data_ram[16][15] ),
    .S(net41),
    .X(_12876_));
 sky130_fd_sc_hd__clkbuf_1 _28753_ (.A(_12876_),
    .X(_04166_));
 sky130_fd_sc_hd__a21oi_4 _28754_ (.A1(_12601_),
    .A2(_10997_),
    .B1(_12795_),
    .Y(_12877_));
 sky130_fd_sc_hd__mux2_1 _28755_ (.A0(_12687_),
    .A1(\datamem.data_ram[15][24] ),
    .S(_12877_),
    .X(_12878_));
 sky130_fd_sc_hd__clkbuf_1 _28756_ (.A(_12878_),
    .X(_04167_));
 sky130_fd_sc_hd__mux2_1 _28757_ (.A0(_12690_),
    .A1(\datamem.data_ram[15][25] ),
    .S(_12877_),
    .X(_12879_));
 sky130_fd_sc_hd__clkbuf_1 _28758_ (.A(_12879_),
    .X(_04168_));
 sky130_fd_sc_hd__mux2_1 _28759_ (.A0(_12692_),
    .A1(\datamem.data_ram[15][26] ),
    .S(_12877_),
    .X(_12880_));
 sky130_fd_sc_hd__clkbuf_1 _28760_ (.A(_12880_),
    .X(_04169_));
 sky130_fd_sc_hd__mux2_1 _28761_ (.A0(_12694_),
    .A1(\datamem.data_ram[15][27] ),
    .S(_12877_),
    .X(_12881_));
 sky130_fd_sc_hd__clkbuf_1 _28762_ (.A(_12881_),
    .X(_04170_));
 sky130_fd_sc_hd__mux2_1 _28763_ (.A0(_12696_),
    .A1(\datamem.data_ram[15][28] ),
    .S(_12877_),
    .X(_12882_));
 sky130_fd_sc_hd__clkbuf_1 _28764_ (.A(_12882_),
    .X(_04171_));
 sky130_fd_sc_hd__mux2_1 _28765_ (.A0(_12698_),
    .A1(\datamem.data_ram[15][29] ),
    .S(_12877_),
    .X(_12883_));
 sky130_fd_sc_hd__clkbuf_1 _28766_ (.A(_12883_),
    .X(_04172_));
 sky130_fd_sc_hd__mux2_1 _28767_ (.A0(_12700_),
    .A1(\datamem.data_ram[15][30] ),
    .S(_12877_),
    .X(_12884_));
 sky130_fd_sc_hd__clkbuf_1 _28768_ (.A(_12884_),
    .X(_04173_));
 sky130_fd_sc_hd__mux2_1 _28769_ (.A0(_12702_),
    .A1(\datamem.data_ram[15][31] ),
    .S(_12877_),
    .X(_12885_));
 sky130_fd_sc_hd__clkbuf_1 _28770_ (.A(_12885_),
    .X(_04174_));
 sky130_fd_sc_hd__buf_8 _28771_ (.A(_06591_),
    .X(_12886_));
 sky130_fd_sc_hd__a21oi_4 _28772_ (.A1(_12601_),
    .A2(_10960_),
    .B1(_12886_),
    .Y(_12887_));
 sky130_fd_sc_hd__mux2_1 _28773_ (.A0(_12751_),
    .A1(\datamem.data_ram[15][16] ),
    .S(_12887_),
    .X(_12888_));
 sky130_fd_sc_hd__clkbuf_1 _28774_ (.A(_12888_),
    .X(_04175_));
 sky130_fd_sc_hd__mux2_1 _28775_ (.A0(_12754_),
    .A1(\datamem.data_ram[15][17] ),
    .S(_12887_),
    .X(_12889_));
 sky130_fd_sc_hd__clkbuf_1 _28776_ (.A(_12889_),
    .X(_04176_));
 sky130_fd_sc_hd__mux2_1 _28777_ (.A0(_12756_),
    .A1(\datamem.data_ram[15][18] ),
    .S(_12887_),
    .X(_12890_));
 sky130_fd_sc_hd__clkbuf_1 _28778_ (.A(_12890_),
    .X(_04177_));
 sky130_fd_sc_hd__mux2_1 _28779_ (.A0(_12758_),
    .A1(\datamem.data_ram[15][19] ),
    .S(_12887_),
    .X(_12891_));
 sky130_fd_sc_hd__clkbuf_1 _28780_ (.A(_12891_),
    .X(_04178_));
 sky130_fd_sc_hd__mux2_1 _28781_ (.A0(_12760_),
    .A1(\datamem.data_ram[15][20] ),
    .S(_12887_),
    .X(_12892_));
 sky130_fd_sc_hd__clkbuf_1 _28782_ (.A(_12892_),
    .X(_04179_));
 sky130_fd_sc_hd__mux2_1 _28783_ (.A0(_12762_),
    .A1(\datamem.data_ram[15][21] ),
    .S(_12887_),
    .X(_12893_));
 sky130_fd_sc_hd__clkbuf_1 _28784_ (.A(_12893_),
    .X(_04180_));
 sky130_fd_sc_hd__mux2_1 _28785_ (.A0(_12764_),
    .A1(\datamem.data_ram[15][22] ),
    .S(_12887_),
    .X(_12894_));
 sky130_fd_sc_hd__clkbuf_1 _28786_ (.A(_12894_),
    .X(_04181_));
 sky130_fd_sc_hd__mux2_1 _28787_ (.A0(_12766_),
    .A1(\datamem.data_ram[15][23] ),
    .S(_12887_),
    .X(_12895_));
 sky130_fd_sc_hd__clkbuf_1 _28788_ (.A(_12895_),
    .X(_04182_));
 sky130_fd_sc_hd__a21oi_2 _28789_ (.A1(_12601_),
    .A2(_11020_),
    .B1(_12886_),
    .Y(_12896_));
 sky130_fd_sc_hd__mux2_1 _28790_ (.A0(_12734_),
    .A1(\datamem.data_ram[15][8] ),
    .S(net70),
    .X(_12897_));
 sky130_fd_sc_hd__clkbuf_1 _28791_ (.A(_12897_),
    .X(_04183_));
 sky130_fd_sc_hd__mux2_1 _28792_ (.A0(_12737_),
    .A1(\datamem.data_ram[15][9] ),
    .S(net70),
    .X(_12898_));
 sky130_fd_sc_hd__clkbuf_1 _28793_ (.A(_12898_),
    .X(_04184_));
 sky130_fd_sc_hd__mux2_1 _28794_ (.A0(_12739_),
    .A1(\datamem.data_ram[15][10] ),
    .S(net70),
    .X(_12899_));
 sky130_fd_sc_hd__clkbuf_1 _28795_ (.A(_12899_),
    .X(_04185_));
 sky130_fd_sc_hd__mux2_1 _28796_ (.A0(_12741_),
    .A1(\datamem.data_ram[15][11] ),
    .S(net70),
    .X(_12900_));
 sky130_fd_sc_hd__clkbuf_1 _28797_ (.A(_12900_),
    .X(_04186_));
 sky130_fd_sc_hd__mux2_1 _28798_ (.A0(_12743_),
    .A1(\datamem.data_ram[15][12] ),
    .S(net70),
    .X(_12901_));
 sky130_fd_sc_hd__clkbuf_1 _28799_ (.A(_12901_),
    .X(_04187_));
 sky130_fd_sc_hd__mux2_1 _28800_ (.A0(_12745_),
    .A1(\datamem.data_ram[15][13] ),
    .S(_12896_),
    .X(_12902_));
 sky130_fd_sc_hd__clkbuf_1 _28801_ (.A(_12902_),
    .X(_04188_));
 sky130_fd_sc_hd__mux2_1 _28802_ (.A0(_12747_),
    .A1(\datamem.data_ram[15][14] ),
    .S(_12896_),
    .X(_12903_));
 sky130_fd_sc_hd__clkbuf_1 _28803_ (.A(_12903_),
    .X(_04189_));
 sky130_fd_sc_hd__mux2_1 _28804_ (.A0(_12749_),
    .A1(\datamem.data_ram[15][15] ),
    .S(_12896_),
    .X(_12904_));
 sky130_fd_sc_hd__clkbuf_1 _28805_ (.A(_12904_),
    .X(_04190_));
 sky130_fd_sc_hd__a21oi_4 _28806_ (.A1(_09225_),
    .A2(_10997_),
    .B1(_12886_),
    .Y(_12905_));
 sky130_fd_sc_hd__mux2_1 _28807_ (.A0(_12687_),
    .A1(\datamem.data_ram[14][24] ),
    .S(_12905_),
    .X(_12906_));
 sky130_fd_sc_hd__clkbuf_1 _28808_ (.A(_12906_),
    .X(_04191_));
 sky130_fd_sc_hd__mux2_1 _28809_ (.A0(_12690_),
    .A1(\datamem.data_ram[14][25] ),
    .S(_12905_),
    .X(_12907_));
 sky130_fd_sc_hd__clkbuf_1 _28810_ (.A(_12907_),
    .X(_04192_));
 sky130_fd_sc_hd__mux2_1 _28811_ (.A0(_12692_),
    .A1(\datamem.data_ram[14][26] ),
    .S(_12905_),
    .X(_12908_));
 sky130_fd_sc_hd__clkbuf_1 _28812_ (.A(_12908_),
    .X(_04193_));
 sky130_fd_sc_hd__mux2_1 _28813_ (.A0(_12694_),
    .A1(\datamem.data_ram[14][27] ),
    .S(_12905_),
    .X(_12909_));
 sky130_fd_sc_hd__clkbuf_1 _28814_ (.A(_12909_),
    .X(_04194_));
 sky130_fd_sc_hd__mux2_1 _28815_ (.A0(_12696_),
    .A1(\datamem.data_ram[14][28] ),
    .S(_12905_),
    .X(_12910_));
 sky130_fd_sc_hd__clkbuf_1 _28816_ (.A(_12910_),
    .X(_04195_));
 sky130_fd_sc_hd__mux2_1 _28817_ (.A0(_12698_),
    .A1(\datamem.data_ram[14][29] ),
    .S(_12905_),
    .X(_12911_));
 sky130_fd_sc_hd__clkbuf_1 _28818_ (.A(_12911_),
    .X(_04196_));
 sky130_fd_sc_hd__mux2_1 _28819_ (.A0(_12700_),
    .A1(\datamem.data_ram[14][30] ),
    .S(_12905_),
    .X(_12912_));
 sky130_fd_sc_hd__clkbuf_1 _28820_ (.A(_12912_),
    .X(_04197_));
 sky130_fd_sc_hd__mux2_1 _28821_ (.A0(_12702_),
    .A1(\datamem.data_ram[14][31] ),
    .S(_12905_),
    .X(_12913_));
 sky130_fd_sc_hd__clkbuf_1 _28822_ (.A(_12913_),
    .X(_04198_));
 sky130_fd_sc_hd__a21oi_4 _28823_ (.A1(_09225_),
    .A2(_10960_),
    .B1(_12886_),
    .Y(_12914_));
 sky130_fd_sc_hd__mux2_1 _28824_ (.A0(_12751_),
    .A1(\datamem.data_ram[14][16] ),
    .S(_12914_),
    .X(_12915_));
 sky130_fd_sc_hd__clkbuf_1 _28825_ (.A(_12915_),
    .X(_04199_));
 sky130_fd_sc_hd__mux2_1 _28826_ (.A0(_12754_),
    .A1(\datamem.data_ram[14][17] ),
    .S(_12914_),
    .X(_12916_));
 sky130_fd_sc_hd__clkbuf_1 _28827_ (.A(_12916_),
    .X(_04200_));
 sky130_fd_sc_hd__mux2_1 _28828_ (.A0(_12756_),
    .A1(\datamem.data_ram[14][18] ),
    .S(_12914_),
    .X(_12917_));
 sky130_fd_sc_hd__clkbuf_1 _28829_ (.A(_12917_),
    .X(_04201_));
 sky130_fd_sc_hd__mux2_1 _28830_ (.A0(_12758_),
    .A1(\datamem.data_ram[14][19] ),
    .S(_12914_),
    .X(_12918_));
 sky130_fd_sc_hd__clkbuf_1 _28831_ (.A(_12918_),
    .X(_04202_));
 sky130_fd_sc_hd__mux2_1 _28832_ (.A0(_12760_),
    .A1(\datamem.data_ram[14][20] ),
    .S(_12914_),
    .X(_12919_));
 sky130_fd_sc_hd__clkbuf_1 _28833_ (.A(_12919_),
    .X(_04203_));
 sky130_fd_sc_hd__mux2_1 _28834_ (.A0(_12762_),
    .A1(\datamem.data_ram[14][21] ),
    .S(_12914_),
    .X(_12920_));
 sky130_fd_sc_hd__clkbuf_1 _28835_ (.A(_12920_),
    .X(_04204_));
 sky130_fd_sc_hd__mux2_1 _28836_ (.A0(_12764_),
    .A1(\datamem.data_ram[14][22] ),
    .S(_12914_),
    .X(_12921_));
 sky130_fd_sc_hd__clkbuf_1 _28837_ (.A(_12921_),
    .X(_04205_));
 sky130_fd_sc_hd__mux2_1 _28838_ (.A0(_12766_),
    .A1(\datamem.data_ram[14][23] ),
    .S(_12914_),
    .X(_12922_));
 sky130_fd_sc_hd__clkbuf_1 _28839_ (.A(_12922_),
    .X(_04206_));
 sky130_fd_sc_hd__a21oi_2 _28840_ (.A1(_09225_),
    .A2(_11020_),
    .B1(_12886_),
    .Y(_12923_));
 sky130_fd_sc_hd__mux2_1 _28841_ (.A0(_12734_),
    .A1(\datamem.data_ram[14][8] ),
    .S(net69),
    .X(_12924_));
 sky130_fd_sc_hd__clkbuf_1 _28842_ (.A(_12924_),
    .X(_04207_));
 sky130_fd_sc_hd__mux2_1 _28843_ (.A0(_12737_),
    .A1(\datamem.data_ram[14][9] ),
    .S(net69),
    .X(_12925_));
 sky130_fd_sc_hd__clkbuf_1 _28844_ (.A(_12925_),
    .X(_04208_));
 sky130_fd_sc_hd__mux2_1 _28845_ (.A0(_12739_),
    .A1(\datamem.data_ram[14][10] ),
    .S(net69),
    .X(_12926_));
 sky130_fd_sc_hd__clkbuf_1 _28846_ (.A(_12926_),
    .X(_04209_));
 sky130_fd_sc_hd__mux2_1 _28847_ (.A0(_12741_),
    .A1(\datamem.data_ram[14][11] ),
    .S(net69),
    .X(_12927_));
 sky130_fd_sc_hd__clkbuf_1 _28848_ (.A(_12927_),
    .X(_04210_));
 sky130_fd_sc_hd__mux2_1 _28849_ (.A0(_12743_),
    .A1(\datamem.data_ram[14][12] ),
    .S(net69),
    .X(_12928_));
 sky130_fd_sc_hd__clkbuf_1 _28850_ (.A(_12928_),
    .X(_04211_));
 sky130_fd_sc_hd__mux2_1 _28851_ (.A0(_12745_),
    .A1(\datamem.data_ram[14][13] ),
    .S(_12923_),
    .X(_12929_));
 sky130_fd_sc_hd__clkbuf_1 _28852_ (.A(_12929_),
    .X(_04212_));
 sky130_fd_sc_hd__mux2_1 _28853_ (.A0(_12747_),
    .A1(\datamem.data_ram[14][14] ),
    .S(_12923_),
    .X(_12930_));
 sky130_fd_sc_hd__clkbuf_1 _28854_ (.A(_12930_),
    .X(_04213_));
 sky130_fd_sc_hd__mux2_1 _28855_ (.A0(_12749_),
    .A1(\datamem.data_ram[14][15] ),
    .S(_12923_),
    .X(_12931_));
 sky130_fd_sc_hd__clkbuf_1 _28856_ (.A(_12931_),
    .X(_04214_));
 sky130_fd_sc_hd__a21oi_4 _28857_ (.A1(_12178_),
    .A2(_10997_),
    .B1(_12886_),
    .Y(_12932_));
 sky130_fd_sc_hd__mux2_1 _28858_ (.A0(_12687_),
    .A1(\datamem.data_ram[13][24] ),
    .S(_12932_),
    .X(_12933_));
 sky130_fd_sc_hd__clkbuf_1 _28859_ (.A(_12933_),
    .X(_04215_));
 sky130_fd_sc_hd__mux2_1 _28860_ (.A0(_12690_),
    .A1(\datamem.data_ram[13][25] ),
    .S(_12932_),
    .X(_12934_));
 sky130_fd_sc_hd__clkbuf_1 _28861_ (.A(_12934_),
    .X(_04216_));
 sky130_fd_sc_hd__mux2_1 _28862_ (.A0(_12692_),
    .A1(\datamem.data_ram[13][26] ),
    .S(_12932_),
    .X(_12935_));
 sky130_fd_sc_hd__clkbuf_1 _28863_ (.A(_12935_),
    .X(_04217_));
 sky130_fd_sc_hd__mux2_1 _28864_ (.A0(_12694_),
    .A1(\datamem.data_ram[13][27] ),
    .S(_12932_),
    .X(_12936_));
 sky130_fd_sc_hd__clkbuf_1 _28865_ (.A(_12936_),
    .X(_04218_));
 sky130_fd_sc_hd__mux2_1 _28866_ (.A0(_12696_),
    .A1(\datamem.data_ram[13][28] ),
    .S(_12932_),
    .X(_12937_));
 sky130_fd_sc_hd__clkbuf_1 _28867_ (.A(_12937_),
    .X(_04219_));
 sky130_fd_sc_hd__mux2_1 _28868_ (.A0(_12698_),
    .A1(\datamem.data_ram[13][29] ),
    .S(_12932_),
    .X(_12938_));
 sky130_fd_sc_hd__clkbuf_1 _28869_ (.A(_12938_),
    .X(_04220_));
 sky130_fd_sc_hd__mux2_1 _28870_ (.A0(_12700_),
    .A1(\datamem.data_ram[13][30] ),
    .S(_12932_),
    .X(_12939_));
 sky130_fd_sc_hd__clkbuf_1 _28871_ (.A(_12939_),
    .X(_04221_));
 sky130_fd_sc_hd__mux2_1 _28872_ (.A0(_12702_),
    .A1(\datamem.data_ram[13][31] ),
    .S(_12932_),
    .X(_12940_));
 sky130_fd_sc_hd__clkbuf_1 _28873_ (.A(_12940_),
    .X(_04222_));
 sky130_fd_sc_hd__a21oi_4 _28874_ (.A1(_12178_),
    .A2(_10960_),
    .B1(_12886_),
    .Y(_12941_));
 sky130_fd_sc_hd__mux2_1 _28875_ (.A0(_12751_),
    .A1(\datamem.data_ram[13][16] ),
    .S(_12941_),
    .X(_12942_));
 sky130_fd_sc_hd__clkbuf_1 _28876_ (.A(_12942_),
    .X(_04223_));
 sky130_fd_sc_hd__mux2_1 _28877_ (.A0(_12754_),
    .A1(\datamem.data_ram[13][17] ),
    .S(_12941_),
    .X(_12943_));
 sky130_fd_sc_hd__clkbuf_1 _28878_ (.A(_12943_),
    .X(_04224_));
 sky130_fd_sc_hd__mux2_1 _28879_ (.A0(_12756_),
    .A1(\datamem.data_ram[13][18] ),
    .S(_12941_),
    .X(_12944_));
 sky130_fd_sc_hd__clkbuf_1 _28880_ (.A(_12944_),
    .X(_04225_));
 sky130_fd_sc_hd__mux2_1 _28881_ (.A0(_12758_),
    .A1(\datamem.data_ram[13][19] ),
    .S(_12941_),
    .X(_12945_));
 sky130_fd_sc_hd__clkbuf_1 _28882_ (.A(_12945_),
    .X(_04226_));
 sky130_fd_sc_hd__mux2_1 _28883_ (.A0(_12760_),
    .A1(\datamem.data_ram[13][20] ),
    .S(_12941_),
    .X(_12946_));
 sky130_fd_sc_hd__clkbuf_1 _28884_ (.A(_12946_),
    .X(_04227_));
 sky130_fd_sc_hd__mux2_1 _28885_ (.A0(_12762_),
    .A1(\datamem.data_ram[13][21] ),
    .S(_12941_),
    .X(_12947_));
 sky130_fd_sc_hd__clkbuf_1 _28886_ (.A(_12947_),
    .X(_04228_));
 sky130_fd_sc_hd__mux2_1 _28887_ (.A0(_12764_),
    .A1(\datamem.data_ram[13][22] ),
    .S(_12941_),
    .X(_12948_));
 sky130_fd_sc_hd__clkbuf_1 _28888_ (.A(_12948_),
    .X(_04229_));
 sky130_fd_sc_hd__mux2_1 _28889_ (.A0(_12766_),
    .A1(\datamem.data_ram[13][23] ),
    .S(_12941_),
    .X(_12949_));
 sky130_fd_sc_hd__clkbuf_1 _28890_ (.A(_12949_),
    .X(_04230_));
 sky130_fd_sc_hd__a21oi_1 _28891_ (.A1(_12178_),
    .A2(_11020_),
    .B1(_12886_),
    .Y(_12950_));
 sky130_fd_sc_hd__mux2_1 _28892_ (.A0(_12734_),
    .A1(\datamem.data_ram[13][8] ),
    .S(net68),
    .X(_12951_));
 sky130_fd_sc_hd__clkbuf_1 _28893_ (.A(_12951_),
    .X(_04231_));
 sky130_fd_sc_hd__mux2_1 _28894_ (.A0(_12737_),
    .A1(\datamem.data_ram[13][9] ),
    .S(net68),
    .X(_12952_));
 sky130_fd_sc_hd__clkbuf_1 _28895_ (.A(_12952_),
    .X(_04232_));
 sky130_fd_sc_hd__mux2_1 _28896_ (.A0(_12739_),
    .A1(\datamem.data_ram[13][10] ),
    .S(net68),
    .X(_12953_));
 sky130_fd_sc_hd__clkbuf_1 _28897_ (.A(_12953_),
    .X(_04233_));
 sky130_fd_sc_hd__mux2_1 _28898_ (.A0(_12741_),
    .A1(\datamem.data_ram[13][11] ),
    .S(net68),
    .X(_12954_));
 sky130_fd_sc_hd__clkbuf_1 _28899_ (.A(_12954_),
    .X(_04234_));
 sky130_fd_sc_hd__mux2_1 _28900_ (.A0(_12743_),
    .A1(\datamem.data_ram[13][12] ),
    .S(net68),
    .X(_12955_));
 sky130_fd_sc_hd__clkbuf_1 _28901_ (.A(_12955_),
    .X(_04235_));
 sky130_fd_sc_hd__mux2_1 _28902_ (.A0(_12745_),
    .A1(\datamem.data_ram[13][13] ),
    .S(net68),
    .X(_12956_));
 sky130_fd_sc_hd__clkbuf_1 _28903_ (.A(_12956_),
    .X(_04236_));
 sky130_fd_sc_hd__mux2_1 _28904_ (.A0(_12747_),
    .A1(\datamem.data_ram[13][14] ),
    .S(net68),
    .X(_12957_));
 sky130_fd_sc_hd__clkbuf_1 _28905_ (.A(_12957_),
    .X(_04237_));
 sky130_fd_sc_hd__mux2_1 _28906_ (.A0(_12749_),
    .A1(\datamem.data_ram[13][15] ),
    .S(net68),
    .X(_12958_));
 sky130_fd_sc_hd__clkbuf_1 _28907_ (.A(_12958_),
    .X(_04238_));
 sky130_fd_sc_hd__a21oi_4 _28908_ (.A1(_09350_),
    .A2(_10997_),
    .B1(_12886_),
    .Y(_12959_));
 sky130_fd_sc_hd__mux2_1 _28909_ (.A0(_12687_),
    .A1(\datamem.data_ram[12][24] ),
    .S(_12959_),
    .X(_12960_));
 sky130_fd_sc_hd__clkbuf_1 _28910_ (.A(_12960_),
    .X(_04239_));
 sky130_fd_sc_hd__mux2_1 _28911_ (.A0(_12690_),
    .A1(\datamem.data_ram[12][25] ),
    .S(_12959_),
    .X(_12961_));
 sky130_fd_sc_hd__clkbuf_1 _28912_ (.A(_12961_),
    .X(_04240_));
 sky130_fd_sc_hd__mux2_1 _28913_ (.A0(_12692_),
    .A1(\datamem.data_ram[12][26] ),
    .S(_12959_),
    .X(_12962_));
 sky130_fd_sc_hd__clkbuf_1 _28914_ (.A(_12962_),
    .X(_04241_));
 sky130_fd_sc_hd__mux2_1 _28915_ (.A0(_12694_),
    .A1(\datamem.data_ram[12][27] ),
    .S(_12959_),
    .X(_12963_));
 sky130_fd_sc_hd__clkbuf_1 _28916_ (.A(_12963_),
    .X(_04242_));
 sky130_fd_sc_hd__mux2_1 _28917_ (.A0(_12696_),
    .A1(\datamem.data_ram[12][28] ),
    .S(_12959_),
    .X(_12964_));
 sky130_fd_sc_hd__clkbuf_1 _28918_ (.A(_12964_),
    .X(_04243_));
 sky130_fd_sc_hd__mux2_1 _28919_ (.A0(_12698_),
    .A1(\datamem.data_ram[12][29] ),
    .S(_12959_),
    .X(_12965_));
 sky130_fd_sc_hd__clkbuf_1 _28920_ (.A(_12965_),
    .X(_04244_));
 sky130_fd_sc_hd__mux2_1 _28921_ (.A0(_12700_),
    .A1(\datamem.data_ram[12][30] ),
    .S(_12959_),
    .X(_12966_));
 sky130_fd_sc_hd__clkbuf_1 _28922_ (.A(_12966_),
    .X(_04245_));
 sky130_fd_sc_hd__mux2_1 _28923_ (.A0(_12702_),
    .A1(\datamem.data_ram[12][31] ),
    .S(_12959_),
    .X(_12967_));
 sky130_fd_sc_hd__clkbuf_1 _28924_ (.A(_12967_),
    .X(_04246_));
 sky130_fd_sc_hd__a21oi_4 _28925_ (.A1(_09350_),
    .A2(_10960_),
    .B1(_12886_),
    .Y(_12968_));
 sky130_fd_sc_hd__mux2_1 _28926_ (.A0(_12751_),
    .A1(\datamem.data_ram[12][16] ),
    .S(_12968_),
    .X(_12969_));
 sky130_fd_sc_hd__clkbuf_1 _28927_ (.A(_12969_),
    .X(_04247_));
 sky130_fd_sc_hd__mux2_1 _28928_ (.A0(_12754_),
    .A1(\datamem.data_ram[12][17] ),
    .S(_12968_),
    .X(_12970_));
 sky130_fd_sc_hd__clkbuf_1 _28929_ (.A(_12970_),
    .X(_04248_));
 sky130_fd_sc_hd__mux2_1 _28930_ (.A0(_12756_),
    .A1(\datamem.data_ram[12][18] ),
    .S(_12968_),
    .X(_12971_));
 sky130_fd_sc_hd__clkbuf_1 _28931_ (.A(_12971_),
    .X(_04249_));
 sky130_fd_sc_hd__mux2_1 _28932_ (.A0(_12758_),
    .A1(\datamem.data_ram[12][19] ),
    .S(_12968_),
    .X(_12972_));
 sky130_fd_sc_hd__clkbuf_1 _28933_ (.A(_12972_),
    .X(_04250_));
 sky130_fd_sc_hd__mux2_1 _28934_ (.A0(_12760_),
    .A1(\datamem.data_ram[12][20] ),
    .S(_12968_),
    .X(_12973_));
 sky130_fd_sc_hd__clkbuf_1 _28935_ (.A(_12973_),
    .X(_04251_));
 sky130_fd_sc_hd__mux2_1 _28936_ (.A0(_12762_),
    .A1(\datamem.data_ram[12][21] ),
    .S(_12968_),
    .X(_12974_));
 sky130_fd_sc_hd__clkbuf_1 _28937_ (.A(_12974_),
    .X(_04252_));
 sky130_fd_sc_hd__mux2_1 _28938_ (.A0(_12764_),
    .A1(\datamem.data_ram[12][22] ),
    .S(_12968_),
    .X(_12975_));
 sky130_fd_sc_hd__clkbuf_1 _28939_ (.A(_12975_),
    .X(_04253_));
 sky130_fd_sc_hd__mux2_1 _28940_ (.A0(_12766_),
    .A1(\datamem.data_ram[12][23] ),
    .S(_12968_),
    .X(_12976_));
 sky130_fd_sc_hd__clkbuf_1 _28941_ (.A(_12976_),
    .X(_04254_));
 sky130_fd_sc_hd__buf_8 _28942_ (.A(_06591_),
    .X(_12977_));
 sky130_fd_sc_hd__a21oi_2 _28943_ (.A1(_09350_),
    .A2(_11020_),
    .B1(_12977_),
    .Y(_12978_));
 sky130_fd_sc_hd__mux2_1 _28944_ (.A0(_12734_),
    .A1(\datamem.data_ram[12][8] ),
    .S(net67),
    .X(_12979_));
 sky130_fd_sc_hd__clkbuf_1 _28945_ (.A(_12979_),
    .X(_04255_));
 sky130_fd_sc_hd__mux2_1 _28946_ (.A0(_12737_),
    .A1(\datamem.data_ram[12][9] ),
    .S(net67),
    .X(_12980_));
 sky130_fd_sc_hd__clkbuf_1 _28947_ (.A(_12980_),
    .X(_04256_));
 sky130_fd_sc_hd__mux2_1 _28948_ (.A0(_12739_),
    .A1(\datamem.data_ram[12][10] ),
    .S(net67),
    .X(_12981_));
 sky130_fd_sc_hd__clkbuf_1 _28949_ (.A(_12981_),
    .X(_04257_));
 sky130_fd_sc_hd__mux2_1 _28950_ (.A0(_12741_),
    .A1(\datamem.data_ram[12][11] ),
    .S(net67),
    .X(_12982_));
 sky130_fd_sc_hd__clkbuf_1 _28951_ (.A(_12982_),
    .X(_04258_));
 sky130_fd_sc_hd__mux2_1 _28952_ (.A0(_12743_),
    .A1(\datamem.data_ram[12][12] ),
    .S(net67),
    .X(_12983_));
 sky130_fd_sc_hd__clkbuf_1 _28953_ (.A(_12983_),
    .X(_04259_));
 sky130_fd_sc_hd__mux2_1 _28954_ (.A0(_12745_),
    .A1(\datamem.data_ram[12][13] ),
    .S(net67),
    .X(_12984_));
 sky130_fd_sc_hd__clkbuf_1 _28955_ (.A(_12984_),
    .X(_04260_));
 sky130_fd_sc_hd__mux2_1 _28956_ (.A0(_12747_),
    .A1(\datamem.data_ram[12][14] ),
    .S(_12978_),
    .X(_12985_));
 sky130_fd_sc_hd__clkbuf_1 _28957_ (.A(_12985_),
    .X(_04261_));
 sky130_fd_sc_hd__mux2_1 _28958_ (.A0(_12749_),
    .A1(\datamem.data_ram[12][15] ),
    .S(_12978_),
    .X(_12986_));
 sky130_fd_sc_hd__clkbuf_1 _28959_ (.A(_12986_),
    .X(_04262_));
 sky130_fd_sc_hd__or3_1 _28960_ (.A(_07791_),
    .B(_10042_),
    .C(_10918_),
    .X(_12987_));
 sky130_fd_sc_hd__buf_2 _28961_ (.A(_12987_),
    .X(_12988_));
 sky130_fd_sc_hd__and3_2 _28962_ (.A(_10325_),
    .B(_10049_),
    .C(_11898_),
    .X(_12989_));
 sky130_fd_sc_hd__and2_1 _28963_ (.A(_10047_),
    .B(_12989_),
    .X(_12990_));
 sky130_fd_sc_hd__a31o_1 _28964_ (.A1(_12727_),
    .A2(\datamem.data_ram[7][0] ),
    .A3(_12988_),
    .B1(_12990_),
    .X(_04263_));
 sky130_fd_sc_hd__and2_1 _28965_ (.A(_10057_),
    .B(_12989_),
    .X(_12991_));
 sky130_fd_sc_hd__a31o_1 _28966_ (.A1(_12727_),
    .A2(\datamem.data_ram[7][1] ),
    .A3(_12988_),
    .B1(_12991_),
    .X(_04264_));
 sky130_fd_sc_hd__and2_1 _28967_ (.A(_10060_),
    .B(_12989_),
    .X(_12992_));
 sky130_fd_sc_hd__a31o_1 _28968_ (.A1(_12727_),
    .A2(\datamem.data_ram[7][2] ),
    .A3(_12988_),
    .B1(_12992_),
    .X(_04265_));
 sky130_fd_sc_hd__and2_1 _28969_ (.A(_10063_),
    .B(_12989_),
    .X(_12993_));
 sky130_fd_sc_hd__a31o_1 _28970_ (.A1(_12727_),
    .A2(\datamem.data_ram[7][3] ),
    .A3(_12988_),
    .B1(_12993_),
    .X(_04266_));
 sky130_fd_sc_hd__and2_1 _28971_ (.A(_10066_),
    .B(_12989_),
    .X(_12994_));
 sky130_fd_sc_hd__a31o_1 _28972_ (.A1(_12727_),
    .A2(\datamem.data_ram[7][4] ),
    .A3(_12988_),
    .B1(_12994_),
    .X(_04267_));
 sky130_fd_sc_hd__clkbuf_4 _28973_ (.A(_06587_),
    .X(_12995_));
 sky130_fd_sc_hd__and2_1 _28974_ (.A(_10069_),
    .B(_12989_),
    .X(_12996_));
 sky130_fd_sc_hd__a31o_1 _28975_ (.A1(_12995_),
    .A2(\datamem.data_ram[7][5] ),
    .A3(_12988_),
    .B1(_12996_),
    .X(_04268_));
 sky130_fd_sc_hd__and2_1 _28976_ (.A(_10072_),
    .B(_12989_),
    .X(_12997_));
 sky130_fd_sc_hd__a31o_1 _28977_ (.A1(_12995_),
    .A2(\datamem.data_ram[7][6] ),
    .A3(_12988_),
    .B1(_12997_),
    .X(_04269_));
 sky130_fd_sc_hd__and2_1 _28978_ (.A(_10075_),
    .B(_12989_),
    .X(_12998_));
 sky130_fd_sc_hd__a31o_1 _28979_ (.A1(_12995_),
    .A2(\datamem.data_ram[7][7] ),
    .A3(_12988_),
    .B1(_12998_),
    .X(_04270_));
 sky130_fd_sc_hd__a21oi_4 _28980_ (.A1(_10141_),
    .A2(_10997_),
    .B1(_12977_),
    .Y(_12999_));
 sky130_fd_sc_hd__mux2_1 _28981_ (.A0(_12687_),
    .A1(\datamem.data_ram[11][24] ),
    .S(_12999_),
    .X(_13000_));
 sky130_fd_sc_hd__clkbuf_1 _28982_ (.A(_13000_),
    .X(_04271_));
 sky130_fd_sc_hd__mux2_1 _28983_ (.A0(_12690_),
    .A1(\datamem.data_ram[11][25] ),
    .S(_12999_),
    .X(_13001_));
 sky130_fd_sc_hd__clkbuf_1 _28984_ (.A(_13001_),
    .X(_04272_));
 sky130_fd_sc_hd__mux2_1 _28985_ (.A0(_12692_),
    .A1(\datamem.data_ram[11][26] ),
    .S(_12999_),
    .X(_13002_));
 sky130_fd_sc_hd__clkbuf_1 _28986_ (.A(_13002_),
    .X(_04273_));
 sky130_fd_sc_hd__mux2_1 _28987_ (.A0(_12694_),
    .A1(\datamem.data_ram[11][27] ),
    .S(_12999_),
    .X(_13003_));
 sky130_fd_sc_hd__clkbuf_1 _28988_ (.A(_13003_),
    .X(_04274_));
 sky130_fd_sc_hd__mux2_1 _28989_ (.A0(_12696_),
    .A1(\datamem.data_ram[11][28] ),
    .S(_12999_),
    .X(_13004_));
 sky130_fd_sc_hd__clkbuf_1 _28990_ (.A(_13004_),
    .X(_04275_));
 sky130_fd_sc_hd__mux2_1 _28991_ (.A0(_12698_),
    .A1(\datamem.data_ram[11][29] ),
    .S(_12999_),
    .X(_13005_));
 sky130_fd_sc_hd__clkbuf_1 _28992_ (.A(_13005_),
    .X(_04276_));
 sky130_fd_sc_hd__mux2_1 _28993_ (.A0(_12700_),
    .A1(\datamem.data_ram[11][30] ),
    .S(_12999_),
    .X(_13006_));
 sky130_fd_sc_hd__clkbuf_1 _28994_ (.A(_13006_),
    .X(_04277_));
 sky130_fd_sc_hd__mux2_1 _28995_ (.A0(_12702_),
    .A1(\datamem.data_ram[11][31] ),
    .S(_12999_),
    .X(_13007_));
 sky130_fd_sc_hd__clkbuf_1 _28996_ (.A(_13007_),
    .X(_04278_));
 sky130_fd_sc_hd__or3_1 _28997_ (.A(_07077_),
    .B(_10932_),
    .C(_10918_),
    .X(_13008_));
 sky130_fd_sc_hd__clkbuf_2 _28998_ (.A(_13008_),
    .X(_13009_));
 sky130_fd_sc_hd__and3_2 _28999_ (.A(_10142_),
    .B(_10935_),
    .C(_10921_),
    .X(_13010_));
 sky130_fd_sc_hd__and2_1 _29000_ (.A(_10047_),
    .B(_13010_),
    .X(_13011_));
 sky130_fd_sc_hd__a31o_1 _29001_ (.A1(_12995_),
    .A2(\datamem.data_ram[11][0] ),
    .A3(_13009_),
    .B1(_13011_),
    .X(_04279_));
 sky130_fd_sc_hd__and2_1 _29002_ (.A(_10057_),
    .B(_13010_),
    .X(_13012_));
 sky130_fd_sc_hd__a31o_1 _29003_ (.A1(_12995_),
    .A2(\datamem.data_ram[11][1] ),
    .A3(_13009_),
    .B1(_13012_),
    .X(_04280_));
 sky130_fd_sc_hd__and2_1 _29004_ (.A(_10060_),
    .B(_13010_),
    .X(_13013_));
 sky130_fd_sc_hd__a31o_1 _29005_ (.A1(_12995_),
    .A2(\datamem.data_ram[11][2] ),
    .A3(_13009_),
    .B1(_13013_),
    .X(_04281_));
 sky130_fd_sc_hd__and2_1 _29006_ (.A(_10063_),
    .B(_13010_),
    .X(_13014_));
 sky130_fd_sc_hd__a31o_1 _29007_ (.A1(_12995_),
    .A2(\datamem.data_ram[11][3] ),
    .A3(_13009_),
    .B1(_13014_),
    .X(_04282_));
 sky130_fd_sc_hd__and2_1 _29008_ (.A(_10066_),
    .B(_13010_),
    .X(_13015_));
 sky130_fd_sc_hd__a31o_1 _29009_ (.A1(_12995_),
    .A2(\datamem.data_ram[11][4] ),
    .A3(_13009_),
    .B1(_13015_),
    .X(_04283_));
 sky130_fd_sc_hd__and2_1 _29010_ (.A(_10069_),
    .B(_13010_),
    .X(_13016_));
 sky130_fd_sc_hd__a31o_1 _29011_ (.A1(_12995_),
    .A2(\datamem.data_ram[11][5] ),
    .A3(_13009_),
    .B1(_13016_),
    .X(_04284_));
 sky130_fd_sc_hd__and2_1 _29012_ (.A(_10072_),
    .B(_13010_),
    .X(_13017_));
 sky130_fd_sc_hd__a31o_1 _29013_ (.A1(_12995_),
    .A2(\datamem.data_ram[11][6] ),
    .A3(_13009_),
    .B1(_13017_),
    .X(_04285_));
 sky130_fd_sc_hd__clkbuf_4 _29014_ (.A(_06587_),
    .X(_13018_));
 sky130_fd_sc_hd__and2_1 _29015_ (.A(_10075_),
    .B(_13010_),
    .X(_13019_));
 sky130_fd_sc_hd__a31o_1 _29016_ (.A1(_13018_),
    .A2(\datamem.data_ram[11][7] ),
    .A3(_13009_),
    .B1(_13019_),
    .X(_04286_));
 sky130_fd_sc_hd__a21oi_2 _29017_ (.A1(_10141_),
    .A2(_11020_),
    .B1(_12977_),
    .Y(_13020_));
 sky130_fd_sc_hd__mux2_1 _29018_ (.A0(_12734_),
    .A1(\datamem.data_ram[11][8] ),
    .S(net66),
    .X(_13021_));
 sky130_fd_sc_hd__clkbuf_1 _29019_ (.A(_13021_),
    .X(_04287_));
 sky130_fd_sc_hd__mux2_1 _29020_ (.A0(_12737_),
    .A1(\datamem.data_ram[11][9] ),
    .S(net66),
    .X(_13022_));
 sky130_fd_sc_hd__clkbuf_1 _29021_ (.A(_13022_),
    .X(_04288_));
 sky130_fd_sc_hd__mux2_1 _29022_ (.A0(_12739_),
    .A1(\datamem.data_ram[11][10] ),
    .S(net66),
    .X(_13023_));
 sky130_fd_sc_hd__clkbuf_1 _29023_ (.A(_13023_),
    .X(_04289_));
 sky130_fd_sc_hd__mux2_1 _29024_ (.A0(_12741_),
    .A1(\datamem.data_ram[11][11] ),
    .S(net66),
    .X(_13024_));
 sky130_fd_sc_hd__clkbuf_1 _29025_ (.A(_13024_),
    .X(_04290_));
 sky130_fd_sc_hd__mux2_1 _29026_ (.A0(_12743_),
    .A1(\datamem.data_ram[11][12] ),
    .S(net66),
    .X(_13025_));
 sky130_fd_sc_hd__clkbuf_1 _29027_ (.A(_13025_),
    .X(_04291_));
 sky130_fd_sc_hd__mux2_1 _29028_ (.A0(_12745_),
    .A1(\datamem.data_ram[11][13] ),
    .S(_13020_),
    .X(_13026_));
 sky130_fd_sc_hd__clkbuf_1 _29029_ (.A(_13026_),
    .X(_04292_));
 sky130_fd_sc_hd__mux2_1 _29030_ (.A0(_12747_),
    .A1(\datamem.data_ram[11][14] ),
    .S(_13020_),
    .X(_13027_));
 sky130_fd_sc_hd__clkbuf_1 _29031_ (.A(_13027_),
    .X(_04293_));
 sky130_fd_sc_hd__mux2_1 _29032_ (.A0(_12749_),
    .A1(\datamem.data_ram[11][15] ),
    .S(_13020_),
    .X(_13028_));
 sky130_fd_sc_hd__clkbuf_1 _29033_ (.A(_13028_),
    .X(_04294_));
 sky130_fd_sc_hd__or2_1 _29034_ (.A(_10932_),
    .B(_10778_),
    .X(_13029_));
 sky130_fd_sc_hd__clkbuf_2 _29035_ (.A(_13029_),
    .X(_13030_));
 sky130_fd_sc_hd__nor2_1 _29036_ (.A(_10932_),
    .B(_10778_),
    .Y(_13031_));
 sky130_fd_sc_hd__and2_1 _29037_ (.A(_10047_),
    .B(_13031_),
    .X(_13032_));
 sky130_fd_sc_hd__a31o_1 _29038_ (.A1(_13018_),
    .A2(\datamem.data_ram[10][0] ),
    .A3(_13030_),
    .B1(_13032_),
    .X(_04295_));
 sky130_fd_sc_hd__and2_1 _29039_ (.A(_10057_),
    .B(_13031_),
    .X(_13033_));
 sky130_fd_sc_hd__a31o_1 _29040_ (.A1(_13018_),
    .A2(\datamem.data_ram[10][1] ),
    .A3(_13030_),
    .B1(_13033_),
    .X(_04296_));
 sky130_fd_sc_hd__and2_1 _29041_ (.A(_10060_),
    .B(_13031_),
    .X(_13034_));
 sky130_fd_sc_hd__a31o_1 _29042_ (.A1(_13018_),
    .A2(\datamem.data_ram[10][2] ),
    .A3(_13030_),
    .B1(_13034_),
    .X(_04297_));
 sky130_fd_sc_hd__and2_1 _29043_ (.A(_10063_),
    .B(_13031_),
    .X(_13035_));
 sky130_fd_sc_hd__a31o_1 _29044_ (.A1(_13018_),
    .A2(\datamem.data_ram[10][3] ),
    .A3(_13030_),
    .B1(_13035_),
    .X(_04298_));
 sky130_fd_sc_hd__and2_1 _29045_ (.A(_10066_),
    .B(_13031_),
    .X(_13036_));
 sky130_fd_sc_hd__a31o_1 _29046_ (.A1(_13018_),
    .A2(\datamem.data_ram[10][4] ),
    .A3(_13030_),
    .B1(_13036_),
    .X(_04299_));
 sky130_fd_sc_hd__and2_1 _29047_ (.A(_10069_),
    .B(_13031_),
    .X(_13037_));
 sky130_fd_sc_hd__a31o_1 _29048_ (.A1(_13018_),
    .A2(\datamem.data_ram[10][5] ),
    .A3(_13030_),
    .B1(_13037_),
    .X(_04300_));
 sky130_fd_sc_hd__and2_1 _29049_ (.A(_10072_),
    .B(_13031_),
    .X(_13038_));
 sky130_fd_sc_hd__a31o_1 _29050_ (.A1(_13018_),
    .A2(\datamem.data_ram[10][6] ),
    .A3(_13030_),
    .B1(_13038_),
    .X(_04301_));
 sky130_fd_sc_hd__and2_1 _29051_ (.A(_10075_),
    .B(_13031_),
    .X(_13039_));
 sky130_fd_sc_hd__a31o_1 _29052_ (.A1(_13018_),
    .A2(\datamem.data_ram[10][7] ),
    .A3(_13030_),
    .B1(_13039_),
    .X(_04302_));
 sky130_fd_sc_hd__a21oi_2 _29053_ (.A1(_10777_),
    .A2(_11020_),
    .B1(_12977_),
    .Y(_13040_));
 sky130_fd_sc_hd__mux2_1 _29054_ (.A0(_09266_),
    .A1(\datamem.data_ram[10][8] ),
    .S(net65),
    .X(_13041_));
 sky130_fd_sc_hd__clkbuf_1 _29055_ (.A(_13041_),
    .X(_04303_));
 sky130_fd_sc_hd__mux2_1 _29056_ (.A0(_09272_),
    .A1(\datamem.data_ram[10][9] ),
    .S(net65),
    .X(_13042_));
 sky130_fd_sc_hd__clkbuf_1 _29057_ (.A(_13042_),
    .X(_04304_));
 sky130_fd_sc_hd__mux2_1 _29058_ (.A0(_09275_),
    .A1(\datamem.data_ram[10][10] ),
    .S(net65),
    .X(_13043_));
 sky130_fd_sc_hd__clkbuf_1 _29059_ (.A(_13043_),
    .X(_04305_));
 sky130_fd_sc_hd__mux2_1 _29060_ (.A0(_09278_),
    .A1(\datamem.data_ram[10][11] ),
    .S(net65),
    .X(_13044_));
 sky130_fd_sc_hd__clkbuf_1 _29061_ (.A(_13044_),
    .X(_04306_));
 sky130_fd_sc_hd__mux2_1 _29062_ (.A0(_09281_),
    .A1(\datamem.data_ram[10][12] ),
    .S(net65),
    .X(_13045_));
 sky130_fd_sc_hd__clkbuf_1 _29063_ (.A(_13045_),
    .X(_04307_));
 sky130_fd_sc_hd__mux2_1 _29064_ (.A0(_09284_),
    .A1(\datamem.data_ram[10][13] ),
    .S(net65),
    .X(_13046_));
 sky130_fd_sc_hd__clkbuf_1 _29065_ (.A(_13046_),
    .X(_04308_));
 sky130_fd_sc_hd__mux2_1 _29066_ (.A0(_09287_),
    .A1(\datamem.data_ram[10][14] ),
    .S(_13040_),
    .X(_13047_));
 sky130_fd_sc_hd__clkbuf_1 _29067_ (.A(_13047_),
    .X(_04309_));
 sky130_fd_sc_hd__mux2_1 _29068_ (.A0(_09290_),
    .A1(\datamem.data_ram[10][15] ),
    .S(_13040_),
    .X(_13048_));
 sky130_fd_sc_hd__clkbuf_1 _29069_ (.A(_13048_),
    .X(_04310_));
 sky130_fd_sc_hd__a21oi_4 _29070_ (.A1(_10777_),
    .A2(_10960_),
    .B1(_12977_),
    .Y(_13049_));
 sky130_fd_sc_hd__mux2_1 _29071_ (.A0(_12751_),
    .A1(\datamem.data_ram[10][16] ),
    .S(_13049_),
    .X(_13050_));
 sky130_fd_sc_hd__clkbuf_1 _29072_ (.A(_13050_),
    .X(_04311_));
 sky130_fd_sc_hd__mux2_1 _29073_ (.A0(_12754_),
    .A1(\datamem.data_ram[10][17] ),
    .S(_13049_),
    .X(_13051_));
 sky130_fd_sc_hd__clkbuf_1 _29074_ (.A(_13051_),
    .X(_04312_));
 sky130_fd_sc_hd__mux2_1 _29075_ (.A0(_12756_),
    .A1(\datamem.data_ram[10][18] ),
    .S(_13049_),
    .X(_13052_));
 sky130_fd_sc_hd__clkbuf_1 _29076_ (.A(_13052_),
    .X(_04313_));
 sky130_fd_sc_hd__mux2_1 _29077_ (.A0(_12758_),
    .A1(\datamem.data_ram[10][19] ),
    .S(_13049_),
    .X(_13053_));
 sky130_fd_sc_hd__clkbuf_1 _29078_ (.A(_13053_),
    .X(_04314_));
 sky130_fd_sc_hd__mux2_1 _29079_ (.A0(_12760_),
    .A1(\datamem.data_ram[10][20] ),
    .S(_13049_),
    .X(_13054_));
 sky130_fd_sc_hd__clkbuf_1 _29080_ (.A(_13054_),
    .X(_04315_));
 sky130_fd_sc_hd__mux2_1 _29081_ (.A0(_12762_),
    .A1(\datamem.data_ram[10][21] ),
    .S(_13049_),
    .X(_13055_));
 sky130_fd_sc_hd__clkbuf_1 _29082_ (.A(_13055_),
    .X(_04316_));
 sky130_fd_sc_hd__mux2_1 _29083_ (.A0(_12764_),
    .A1(\datamem.data_ram[10][22] ),
    .S(_13049_),
    .X(_13056_));
 sky130_fd_sc_hd__clkbuf_1 _29084_ (.A(_13056_),
    .X(_04317_));
 sky130_fd_sc_hd__mux2_1 _29085_ (.A0(_12766_),
    .A1(\datamem.data_ram[10][23] ),
    .S(_13049_),
    .X(_13057_));
 sky130_fd_sc_hd__clkbuf_1 _29086_ (.A(_13057_),
    .X(_04318_));
 sky130_fd_sc_hd__a21oi_4 _29087_ (.A1(_10979_),
    .A2(_11123_),
    .B1(_12977_),
    .Y(_13058_));
 sky130_fd_sc_hd__mux2_1 _29088_ (.A0(_09297_),
    .A1(\datamem.data_ram[0][24] ),
    .S(net40),
    .X(_13059_));
 sky130_fd_sc_hd__clkbuf_1 _29089_ (.A(_13059_),
    .X(_04319_));
 sky130_fd_sc_hd__mux2_1 _29090_ (.A0(_09305_),
    .A1(\datamem.data_ram[0][25] ),
    .S(net40),
    .X(_13060_));
 sky130_fd_sc_hd__clkbuf_1 _29091_ (.A(_13060_),
    .X(_04320_));
 sky130_fd_sc_hd__mux2_1 _29092_ (.A0(_09309_),
    .A1(\datamem.data_ram[0][26] ),
    .S(_13058_),
    .X(_13061_));
 sky130_fd_sc_hd__clkbuf_1 _29093_ (.A(_13061_),
    .X(_04321_));
 sky130_fd_sc_hd__mux2_1 _29094_ (.A0(_09313_),
    .A1(\datamem.data_ram[0][27] ),
    .S(net40),
    .X(_13062_));
 sky130_fd_sc_hd__clkbuf_1 _29095_ (.A(_13062_),
    .X(_04322_));
 sky130_fd_sc_hd__mux2_1 _29096_ (.A0(_09317_),
    .A1(\datamem.data_ram[0][28] ),
    .S(net40),
    .X(_13063_));
 sky130_fd_sc_hd__clkbuf_1 _29097_ (.A(_13063_),
    .X(_04323_));
 sky130_fd_sc_hd__mux2_1 _29098_ (.A0(_09321_),
    .A1(\datamem.data_ram[0][29] ),
    .S(net40),
    .X(_13064_));
 sky130_fd_sc_hd__clkbuf_1 _29099_ (.A(_13064_),
    .X(_04324_));
 sky130_fd_sc_hd__mux2_1 _29100_ (.A0(_09325_),
    .A1(\datamem.data_ram[0][30] ),
    .S(_13058_),
    .X(_13065_));
 sky130_fd_sc_hd__clkbuf_1 _29101_ (.A(_13065_),
    .X(_04325_));
 sky130_fd_sc_hd__mux2_1 _29102_ (.A0(_09329_),
    .A1(\datamem.data_ram[0][31] ),
    .S(_13058_),
    .X(_13066_));
 sky130_fd_sc_hd__clkbuf_1 _29103_ (.A(_13066_),
    .X(_04326_));
 sky130_fd_sc_hd__a21oi_4 _29104_ (.A1(_12601_),
    .A2(_10092_),
    .B1(_12977_),
    .Y(_13067_));
 sky130_fd_sc_hd__mux2_1 _29105_ (.A0(_09266_),
    .A1(\datamem.data_ram[7][8] ),
    .S(_13067_),
    .X(_13068_));
 sky130_fd_sc_hd__clkbuf_1 _29106_ (.A(_13068_),
    .X(_04327_));
 sky130_fd_sc_hd__mux2_1 _29107_ (.A0(_09272_),
    .A1(\datamem.data_ram[7][9] ),
    .S(_13067_),
    .X(_13069_));
 sky130_fd_sc_hd__clkbuf_1 _29108_ (.A(_13069_),
    .X(_04328_));
 sky130_fd_sc_hd__mux2_1 _29109_ (.A0(_09275_),
    .A1(\datamem.data_ram[7][10] ),
    .S(_13067_),
    .X(_13070_));
 sky130_fd_sc_hd__clkbuf_1 _29110_ (.A(_13070_),
    .X(_04329_));
 sky130_fd_sc_hd__mux2_1 _29111_ (.A0(_09278_),
    .A1(\datamem.data_ram[7][11] ),
    .S(_13067_),
    .X(_13071_));
 sky130_fd_sc_hd__clkbuf_1 _29112_ (.A(_13071_),
    .X(_04330_));
 sky130_fd_sc_hd__mux2_1 _29113_ (.A0(_09281_),
    .A1(\datamem.data_ram[7][12] ),
    .S(_13067_),
    .X(_13072_));
 sky130_fd_sc_hd__clkbuf_1 _29114_ (.A(_13072_),
    .X(_04331_));
 sky130_fd_sc_hd__mux2_1 _29115_ (.A0(_09284_),
    .A1(\datamem.data_ram[7][13] ),
    .S(_13067_),
    .X(_13073_));
 sky130_fd_sc_hd__clkbuf_1 _29116_ (.A(_13073_),
    .X(_04332_));
 sky130_fd_sc_hd__mux2_1 _29117_ (.A0(_09287_),
    .A1(\datamem.data_ram[7][14] ),
    .S(_13067_),
    .X(_13074_));
 sky130_fd_sc_hd__clkbuf_1 _29118_ (.A(_13074_),
    .X(_04333_));
 sky130_fd_sc_hd__mux2_1 _29119_ (.A0(_09290_),
    .A1(\datamem.data_ram[7][15] ),
    .S(_13067_),
    .X(_13075_));
 sky130_fd_sc_hd__clkbuf_1 _29120_ (.A(_13075_),
    .X(_04334_));
 sky130_fd_sc_hd__a21oi_4 _29121_ (.A1(_10979_),
    .A2(_10114_),
    .B1(_12977_),
    .Y(_13076_));
 sky130_fd_sc_hd__mux2_1 _29122_ (.A0(_09223_),
    .A1(\datamem.data_ram[0][16] ),
    .S(_13076_),
    .X(_13077_));
 sky130_fd_sc_hd__clkbuf_1 _29123_ (.A(_13077_),
    .X(_04335_));
 sky130_fd_sc_hd__mux2_1 _29124_ (.A0(_09235_),
    .A1(\datamem.data_ram[0][17] ),
    .S(_13076_),
    .X(_13078_));
 sky130_fd_sc_hd__clkbuf_1 _29125_ (.A(_13078_),
    .X(_04336_));
 sky130_fd_sc_hd__mux2_1 _29126_ (.A0(_09239_),
    .A1(\datamem.data_ram[0][18] ),
    .S(_13076_),
    .X(_13079_));
 sky130_fd_sc_hd__clkbuf_1 _29127_ (.A(_13079_),
    .X(_04337_));
 sky130_fd_sc_hd__mux2_1 _29128_ (.A0(_09243_),
    .A1(\datamem.data_ram[0][19] ),
    .S(_13076_),
    .X(_13080_));
 sky130_fd_sc_hd__clkbuf_1 _29129_ (.A(_13080_),
    .X(_04338_));
 sky130_fd_sc_hd__mux2_1 _29130_ (.A0(_09247_),
    .A1(\datamem.data_ram[0][20] ),
    .S(_13076_),
    .X(_13081_));
 sky130_fd_sc_hd__clkbuf_1 _29131_ (.A(_13081_),
    .X(_04339_));
 sky130_fd_sc_hd__mux2_1 _29132_ (.A0(_09251_),
    .A1(\datamem.data_ram[0][21] ),
    .S(_13076_),
    .X(_13082_));
 sky130_fd_sc_hd__clkbuf_1 _29133_ (.A(_13082_),
    .X(_04340_));
 sky130_fd_sc_hd__mux2_1 _29134_ (.A0(_09255_),
    .A1(\datamem.data_ram[0][22] ),
    .S(_13076_),
    .X(_13083_));
 sky130_fd_sc_hd__clkbuf_1 _29135_ (.A(_13083_),
    .X(_04341_));
 sky130_fd_sc_hd__mux2_1 _29136_ (.A0(_09259_),
    .A1(\datamem.data_ram[0][23] ),
    .S(_13076_),
    .X(_13084_));
 sky130_fd_sc_hd__clkbuf_1 _29137_ (.A(_13084_),
    .X(_04342_));
 sky130_fd_sc_hd__a21oi_4 _29138_ (.A1(_10979_),
    .A2(_10092_),
    .B1(_12977_),
    .Y(_13085_));
 sky130_fd_sc_hd__mux2_1 _29139_ (.A0(_09266_),
    .A1(\datamem.data_ram[0][8] ),
    .S(net39),
    .X(_13086_));
 sky130_fd_sc_hd__clkbuf_1 _29140_ (.A(_13086_),
    .X(_04343_));
 sky130_fd_sc_hd__mux2_1 _29141_ (.A0(_09272_),
    .A1(\datamem.data_ram[0][9] ),
    .S(net39),
    .X(_13087_));
 sky130_fd_sc_hd__clkbuf_1 _29142_ (.A(_13087_),
    .X(_04344_));
 sky130_fd_sc_hd__mux2_1 _29143_ (.A0(_09275_),
    .A1(\datamem.data_ram[0][10] ),
    .S(net39),
    .X(_13088_));
 sky130_fd_sc_hd__clkbuf_1 _29144_ (.A(_13088_),
    .X(_04345_));
 sky130_fd_sc_hd__mux2_1 _29145_ (.A0(_09278_),
    .A1(\datamem.data_ram[0][11] ),
    .S(net39),
    .X(_13089_));
 sky130_fd_sc_hd__clkbuf_1 _29146_ (.A(_13089_),
    .X(_04346_));
 sky130_fd_sc_hd__mux2_1 _29147_ (.A0(_09281_),
    .A1(\datamem.data_ram[0][12] ),
    .S(net39),
    .X(_13090_));
 sky130_fd_sc_hd__clkbuf_1 _29148_ (.A(_13090_),
    .X(_04347_));
 sky130_fd_sc_hd__mux2_1 _29149_ (.A0(_09284_),
    .A1(\datamem.data_ram[0][13] ),
    .S(_13085_),
    .X(_13091_));
 sky130_fd_sc_hd__clkbuf_1 _29150_ (.A(_13091_),
    .X(_04348_));
 sky130_fd_sc_hd__mux2_1 _29151_ (.A0(_09287_),
    .A1(\datamem.data_ram[0][14] ),
    .S(_13085_),
    .X(_13092_));
 sky130_fd_sc_hd__clkbuf_1 _29152_ (.A(_13092_),
    .X(_04349_));
 sky130_fd_sc_hd__mux2_1 _29153_ (.A0(_09290_),
    .A1(\datamem.data_ram[0][15] ),
    .S(_13085_),
    .X(_13093_));
 sky130_fd_sc_hd__clkbuf_1 _29154_ (.A(_13093_),
    .X(_04350_));
 sky130_fd_sc_hd__a21oi_4 _29155_ (.A1(_12601_),
    .A2(_10114_),
    .B1(_12977_),
    .Y(_13094_));
 sky130_fd_sc_hd__mux2_1 _29156_ (.A0(_09223_),
    .A1(\datamem.data_ram[7][16] ),
    .S(net64),
    .X(_13095_));
 sky130_fd_sc_hd__clkbuf_1 _29157_ (.A(_13095_),
    .X(_04351_));
 sky130_fd_sc_hd__mux2_1 _29158_ (.A0(_09235_),
    .A1(\datamem.data_ram[7][17] ),
    .S(_13094_),
    .X(_13096_));
 sky130_fd_sc_hd__clkbuf_1 _29159_ (.A(_13096_),
    .X(_04352_));
 sky130_fd_sc_hd__mux2_1 _29160_ (.A0(_09239_),
    .A1(\datamem.data_ram[7][18] ),
    .S(net64),
    .X(_13097_));
 sky130_fd_sc_hd__clkbuf_1 _29161_ (.A(_13097_),
    .X(_04353_));
 sky130_fd_sc_hd__mux2_1 _29162_ (.A0(_09243_),
    .A1(\datamem.data_ram[7][19] ),
    .S(_13094_),
    .X(_13098_));
 sky130_fd_sc_hd__clkbuf_1 _29163_ (.A(_13098_),
    .X(_04354_));
 sky130_fd_sc_hd__mux2_1 _29164_ (.A0(_09247_),
    .A1(\datamem.data_ram[7][20] ),
    .S(net64),
    .X(_13099_));
 sky130_fd_sc_hd__clkbuf_1 _29165_ (.A(_13099_),
    .X(_04355_));
 sky130_fd_sc_hd__mux2_1 _29166_ (.A0(_09251_),
    .A1(\datamem.data_ram[7][21] ),
    .S(_13094_),
    .X(_13100_));
 sky130_fd_sc_hd__clkbuf_1 _29167_ (.A(_13100_),
    .X(_04356_));
 sky130_fd_sc_hd__mux2_1 _29168_ (.A0(_09255_),
    .A1(\datamem.data_ram[7][22] ),
    .S(net64),
    .X(_13101_));
 sky130_fd_sc_hd__clkbuf_1 _29169_ (.A(_13101_),
    .X(_04357_));
 sky130_fd_sc_hd__mux2_1 _29170_ (.A0(_09259_),
    .A1(\datamem.data_ram[7][23] ),
    .S(net64),
    .X(_13102_));
 sky130_fd_sc_hd__clkbuf_1 _29171_ (.A(_13102_),
    .X(_04358_));
 sky130_fd_sc_hd__a21oi_2 _29172_ (.A1(_09225_),
    .A2(_10114_),
    .B1(_09230_),
    .Y(_13103_));
 sky130_fd_sc_hd__mux2_1 _29173_ (.A0(_09223_),
    .A1(\datamem.data_ram[6][16] ),
    .S(net63),
    .X(_13104_));
 sky130_fd_sc_hd__clkbuf_1 _29174_ (.A(_13104_),
    .X(_04359_));
 sky130_fd_sc_hd__mux2_1 _29175_ (.A0(_09235_),
    .A1(\datamem.data_ram[6][17] ),
    .S(net63),
    .X(_13105_));
 sky130_fd_sc_hd__clkbuf_1 _29176_ (.A(_13105_),
    .X(_04360_));
 sky130_fd_sc_hd__mux2_1 _29177_ (.A0(_09239_),
    .A1(\datamem.data_ram[6][18] ),
    .S(net63),
    .X(_13106_));
 sky130_fd_sc_hd__clkbuf_1 _29178_ (.A(_13106_),
    .X(_04361_));
 sky130_fd_sc_hd__mux2_1 _29179_ (.A0(_09243_),
    .A1(\datamem.data_ram[6][19] ),
    .S(net63),
    .X(_13107_));
 sky130_fd_sc_hd__clkbuf_1 _29180_ (.A(_13107_),
    .X(_04362_));
 sky130_fd_sc_hd__mux2_1 _29181_ (.A0(_09247_),
    .A1(\datamem.data_ram[6][20] ),
    .S(net63),
    .X(_13108_));
 sky130_fd_sc_hd__clkbuf_1 _29182_ (.A(_13108_),
    .X(_04363_));
 sky130_fd_sc_hd__mux2_1 _29183_ (.A0(_09251_),
    .A1(\datamem.data_ram[6][21] ),
    .S(net63),
    .X(_13109_));
 sky130_fd_sc_hd__clkbuf_1 _29184_ (.A(_13109_),
    .X(_04364_));
 sky130_fd_sc_hd__mux2_1 _29185_ (.A0(_09255_),
    .A1(\datamem.data_ram[6][22] ),
    .S(net63),
    .X(_13110_));
 sky130_fd_sc_hd__clkbuf_1 _29186_ (.A(_13110_),
    .X(_04365_));
 sky130_fd_sc_hd__mux2_1 _29187_ (.A0(_09259_),
    .A1(\datamem.data_ram[6][23] ),
    .S(_13103_),
    .X(_13111_));
 sky130_fd_sc_hd__clkbuf_1 _29188_ (.A(_13111_),
    .X(_04366_));
 sky130_fd_sc_hd__a21oi_4 _29189_ (.A1(_09225_),
    .A2(_11123_),
    .B1(_09230_),
    .Y(_13112_));
 sky130_fd_sc_hd__mux2_1 _29190_ (.A0(_09297_),
    .A1(\datamem.data_ram[6][24] ),
    .S(_13112_),
    .X(_13113_));
 sky130_fd_sc_hd__clkbuf_1 _29191_ (.A(_13113_),
    .X(_04367_));
 sky130_fd_sc_hd__mux2_1 _29192_ (.A0(_09305_),
    .A1(\datamem.data_ram[6][25] ),
    .S(_13112_),
    .X(_13114_));
 sky130_fd_sc_hd__clkbuf_1 _29193_ (.A(_13114_),
    .X(_04368_));
 sky130_fd_sc_hd__mux2_1 _29194_ (.A0(_09309_),
    .A1(\datamem.data_ram[6][26] ),
    .S(_13112_),
    .X(_13115_));
 sky130_fd_sc_hd__clkbuf_1 _29195_ (.A(_13115_),
    .X(_04369_));
 sky130_fd_sc_hd__mux2_1 _29196_ (.A0(_09313_),
    .A1(\datamem.data_ram[6][27] ),
    .S(_13112_),
    .X(_13116_));
 sky130_fd_sc_hd__clkbuf_1 _29197_ (.A(_13116_),
    .X(_04370_));
 sky130_fd_sc_hd__mux2_1 _29198_ (.A0(_09317_),
    .A1(\datamem.data_ram[6][28] ),
    .S(_13112_),
    .X(_13117_));
 sky130_fd_sc_hd__clkbuf_1 _29199_ (.A(_13117_),
    .X(_04371_));
 sky130_fd_sc_hd__mux2_1 _29200_ (.A0(_09321_),
    .A1(\datamem.data_ram[6][29] ),
    .S(_13112_),
    .X(_13118_));
 sky130_fd_sc_hd__clkbuf_1 _29201_ (.A(_13118_),
    .X(_04372_));
 sky130_fd_sc_hd__mux2_1 _29202_ (.A0(_09325_),
    .A1(\datamem.data_ram[6][30] ),
    .S(_13112_),
    .X(_13119_));
 sky130_fd_sc_hd__clkbuf_1 _29203_ (.A(_13119_),
    .X(_04373_));
 sky130_fd_sc_hd__mux2_1 _29204_ (.A0(_09329_),
    .A1(\datamem.data_ram[6][31] ),
    .S(_13112_),
    .X(_13120_));
 sky130_fd_sc_hd__clkbuf_1 _29205_ (.A(_13120_),
    .X(_04374_));
 sky130_fd_sc_hd__or2_1 _29206_ (.A(_10042_),
    .B(_10947_),
    .X(_13121_));
 sky130_fd_sc_hd__buf_2 _29207_ (.A(_13121_),
    .X(_13122_));
 sky130_fd_sc_hd__nor2_2 _29208_ (.A(_10042_),
    .B(_10947_),
    .Y(_13123_));
 sky130_fd_sc_hd__and2_1 _29209_ (.A(_10047_),
    .B(_13123_),
    .X(_13124_));
 sky130_fd_sc_hd__a31o_1 _29210_ (.A1(_13018_),
    .A2(\datamem.data_ram[6][0] ),
    .A3(_13122_),
    .B1(_13124_),
    .X(_04375_));
 sky130_fd_sc_hd__and2_1 _29211_ (.A(_10057_),
    .B(_13123_),
    .X(_13125_));
 sky130_fd_sc_hd__a31o_1 _29212_ (.A1(_11533_),
    .A2(\datamem.data_ram[6][1] ),
    .A3(_13122_),
    .B1(_13125_),
    .X(_04376_));
 sky130_fd_sc_hd__and2_1 _29213_ (.A(_10060_),
    .B(_13123_),
    .X(_13126_));
 sky130_fd_sc_hd__a31o_1 _29214_ (.A1(_11533_),
    .A2(\datamem.data_ram[6][2] ),
    .A3(_13122_),
    .B1(_13126_),
    .X(_04377_));
 sky130_fd_sc_hd__and2_1 _29215_ (.A(_10063_),
    .B(_13123_),
    .X(_13127_));
 sky130_fd_sc_hd__a31o_1 _29216_ (.A1(_11533_),
    .A2(\datamem.data_ram[6][3] ),
    .A3(_13122_),
    .B1(_13127_),
    .X(_04378_));
 sky130_fd_sc_hd__and2_1 _29217_ (.A(_10066_),
    .B(_13123_),
    .X(_13128_));
 sky130_fd_sc_hd__a31o_1 _29218_ (.A1(_11533_),
    .A2(\datamem.data_ram[6][4] ),
    .A3(_13122_),
    .B1(_13128_),
    .X(_04379_));
 sky130_fd_sc_hd__and2_1 _29219_ (.A(_10069_),
    .B(_13123_),
    .X(_13129_));
 sky130_fd_sc_hd__a31o_1 _29220_ (.A1(_11533_),
    .A2(\datamem.data_ram[6][5] ),
    .A3(_13122_),
    .B1(_13129_),
    .X(_04380_));
 sky130_fd_sc_hd__and2_1 _29221_ (.A(_10072_),
    .B(_13123_),
    .X(_13130_));
 sky130_fd_sc_hd__a31o_1 _29222_ (.A1(_11533_),
    .A2(\datamem.data_ram[6][6] ),
    .A3(_13122_),
    .B1(_13130_),
    .X(_04381_));
 sky130_fd_sc_hd__and2_1 _29223_ (.A(_10075_),
    .B(_13123_),
    .X(_13131_));
 sky130_fd_sc_hd__a31o_1 _29224_ (.A1(_11533_),
    .A2(\datamem.data_ram[6][7] ),
    .A3(_13122_),
    .B1(_13131_),
    .X(_04382_));
 sky130_fd_sc_hd__a21oi_4 _29225_ (.A1(_12601_),
    .A2(_09301_),
    .B1(_09230_),
    .Y(_13132_));
 sky130_fd_sc_hd__mux2_1 _29226_ (.A0(_09297_),
    .A1(\datamem.data_ram[63][24] ),
    .S(_13132_),
    .X(_13133_));
 sky130_fd_sc_hd__clkbuf_1 _29227_ (.A(_13133_),
    .X(_04383_));
 sky130_fd_sc_hd__mux2_1 _29228_ (.A0(_09305_),
    .A1(\datamem.data_ram[63][25] ),
    .S(_13132_),
    .X(_13134_));
 sky130_fd_sc_hd__clkbuf_1 _29229_ (.A(_13134_),
    .X(_04384_));
 sky130_fd_sc_hd__mux2_1 _29230_ (.A0(_09309_),
    .A1(\datamem.data_ram[63][26] ),
    .S(_13132_),
    .X(_13135_));
 sky130_fd_sc_hd__clkbuf_1 _29231_ (.A(_13135_),
    .X(_04385_));
 sky130_fd_sc_hd__mux2_1 _29232_ (.A0(_09313_),
    .A1(\datamem.data_ram[63][27] ),
    .S(_13132_),
    .X(_13136_));
 sky130_fd_sc_hd__clkbuf_1 _29233_ (.A(_13136_),
    .X(_04386_));
 sky130_fd_sc_hd__mux2_1 _29234_ (.A0(_09317_),
    .A1(\datamem.data_ram[63][28] ),
    .S(_13132_),
    .X(_13137_));
 sky130_fd_sc_hd__clkbuf_1 _29235_ (.A(_13137_),
    .X(_04387_));
 sky130_fd_sc_hd__mux2_1 _29236_ (.A0(_09321_),
    .A1(\datamem.data_ram[63][29] ),
    .S(_13132_),
    .X(_13138_));
 sky130_fd_sc_hd__clkbuf_1 _29237_ (.A(_13138_),
    .X(_04388_));
 sky130_fd_sc_hd__mux2_1 _29238_ (.A0(_09325_),
    .A1(\datamem.data_ram[63][30] ),
    .S(_13132_),
    .X(_13139_));
 sky130_fd_sc_hd__clkbuf_1 _29239_ (.A(_13139_),
    .X(_04389_));
 sky130_fd_sc_hd__mux2_1 _29240_ (.A0(_09329_),
    .A1(\datamem.data_ram[63][31] ),
    .S(_13132_),
    .X(_13140_));
 sky130_fd_sc_hd__clkbuf_1 _29241_ (.A(_13140_),
    .X(_04390_));
 sky130_fd_sc_hd__a21oi_4 _29242_ (.A1(_12601_),
    .A2(_09229_),
    .B1(_09230_),
    .Y(_13141_));
 sky130_fd_sc_hd__mux2_1 _29243_ (.A0(_09223_),
    .A1(\datamem.data_ram[63][16] ),
    .S(_13141_),
    .X(_13142_));
 sky130_fd_sc_hd__clkbuf_1 _29244_ (.A(_13142_),
    .X(_04391_));
 sky130_fd_sc_hd__mux2_1 _29245_ (.A0(_09235_),
    .A1(\datamem.data_ram[63][17] ),
    .S(_13141_),
    .X(_13143_));
 sky130_fd_sc_hd__clkbuf_1 _29246_ (.A(_13143_),
    .X(_04392_));
 sky130_fd_sc_hd__mux2_1 _29247_ (.A0(_09239_),
    .A1(\datamem.data_ram[63][18] ),
    .S(_13141_),
    .X(_13144_));
 sky130_fd_sc_hd__clkbuf_1 _29248_ (.A(_13144_),
    .X(_04393_));
 sky130_fd_sc_hd__mux2_1 _29249_ (.A0(_09243_),
    .A1(\datamem.data_ram[63][19] ),
    .S(_13141_),
    .X(_13145_));
 sky130_fd_sc_hd__clkbuf_1 _29250_ (.A(_13145_),
    .X(_04394_));
 sky130_fd_sc_hd__mux2_1 _29251_ (.A0(_09247_),
    .A1(\datamem.data_ram[63][20] ),
    .S(_13141_),
    .X(_13146_));
 sky130_fd_sc_hd__clkbuf_1 _29252_ (.A(_13146_),
    .X(_04395_));
 sky130_fd_sc_hd__mux2_1 _29253_ (.A0(_09251_),
    .A1(\datamem.data_ram[63][21] ),
    .S(_13141_),
    .X(_13147_));
 sky130_fd_sc_hd__clkbuf_1 _29254_ (.A(_13147_),
    .X(_04396_));
 sky130_fd_sc_hd__mux2_1 _29255_ (.A0(_09255_),
    .A1(\datamem.data_ram[63][22] ),
    .S(_13141_),
    .X(_13148_));
 sky130_fd_sc_hd__clkbuf_1 _29256_ (.A(_13148_),
    .X(_04397_));
 sky130_fd_sc_hd__mux2_1 _29257_ (.A0(_09259_),
    .A1(\datamem.data_ram[63][23] ),
    .S(_13141_),
    .X(_13149_));
 sky130_fd_sc_hd__clkbuf_1 _29258_ (.A(_13149_),
    .X(_04398_));
 sky130_fd_sc_hd__a21oi_4 _29259_ (.A1(_07125_),
    .A2(_09269_),
    .B1(_09230_),
    .Y(_13150_));
 sky130_fd_sc_hd__mux2_1 _29260_ (.A0(_09266_),
    .A1(\datamem.data_ram[63][8] ),
    .S(_13150_),
    .X(_13151_));
 sky130_fd_sc_hd__clkbuf_1 _29261_ (.A(_13151_),
    .X(_04399_));
 sky130_fd_sc_hd__mux2_1 _29262_ (.A0(_09272_),
    .A1(\datamem.data_ram[63][9] ),
    .S(_13150_),
    .X(_13152_));
 sky130_fd_sc_hd__clkbuf_1 _29263_ (.A(_13152_),
    .X(_04400_));
 sky130_fd_sc_hd__mux2_1 _29264_ (.A0(_09275_),
    .A1(\datamem.data_ram[63][10] ),
    .S(_13150_),
    .X(_13153_));
 sky130_fd_sc_hd__clkbuf_1 _29265_ (.A(_13153_),
    .X(_04401_));
 sky130_fd_sc_hd__mux2_1 _29266_ (.A0(_09278_),
    .A1(\datamem.data_ram[63][11] ),
    .S(_13150_),
    .X(_13154_));
 sky130_fd_sc_hd__clkbuf_1 _29267_ (.A(_13154_),
    .X(_04402_));
 sky130_fd_sc_hd__mux2_1 _29268_ (.A0(_09281_),
    .A1(\datamem.data_ram[63][12] ),
    .S(_13150_),
    .X(_13155_));
 sky130_fd_sc_hd__clkbuf_1 _29269_ (.A(_13155_),
    .X(_04403_));
 sky130_fd_sc_hd__mux2_1 _29270_ (.A0(_09284_),
    .A1(\datamem.data_ram[63][13] ),
    .S(_13150_),
    .X(_13156_));
 sky130_fd_sc_hd__clkbuf_1 _29271_ (.A(_13156_),
    .X(_04404_));
 sky130_fd_sc_hd__mux2_1 _29272_ (.A0(_09287_),
    .A1(\datamem.data_ram[63][14] ),
    .S(_13150_),
    .X(_13157_));
 sky130_fd_sc_hd__clkbuf_1 _29273_ (.A(_13157_),
    .X(_04405_));
 sky130_fd_sc_hd__mux2_1 _29274_ (.A0(_09290_),
    .A1(\datamem.data_ram[63][15] ),
    .S(_13150_),
    .X(_13158_));
 sky130_fd_sc_hd__clkbuf_1 _29275_ (.A(_13158_),
    .X(_04406_));
 sky130_fd_sc_hd__a21oi_4 _29276_ (.A1(_09225_),
    .A2(_09301_),
    .B1(_09230_),
    .Y(_13159_));
 sky130_fd_sc_hd__mux2_1 _29277_ (.A0(_09297_),
    .A1(\datamem.data_ram[62][24] ),
    .S(_13159_),
    .X(_13160_));
 sky130_fd_sc_hd__clkbuf_1 _29278_ (.A(_13160_),
    .X(_04407_));
 sky130_fd_sc_hd__mux2_1 _29279_ (.A0(_09305_),
    .A1(\datamem.data_ram[62][25] ),
    .S(_13159_),
    .X(_13161_));
 sky130_fd_sc_hd__clkbuf_1 _29280_ (.A(_13161_),
    .X(_04408_));
 sky130_fd_sc_hd__mux2_1 _29281_ (.A0(_09309_),
    .A1(\datamem.data_ram[62][26] ),
    .S(_13159_),
    .X(_13162_));
 sky130_fd_sc_hd__clkbuf_1 _29282_ (.A(_13162_),
    .X(_04409_));
 sky130_fd_sc_hd__mux2_1 _29283_ (.A0(_09313_),
    .A1(\datamem.data_ram[62][27] ),
    .S(_13159_),
    .X(_13163_));
 sky130_fd_sc_hd__clkbuf_1 _29284_ (.A(_13163_),
    .X(_04410_));
 sky130_fd_sc_hd__mux2_1 _29285_ (.A0(_09317_),
    .A1(\datamem.data_ram[62][28] ),
    .S(_13159_),
    .X(_13164_));
 sky130_fd_sc_hd__clkbuf_1 _29286_ (.A(_13164_),
    .X(_04411_));
 sky130_fd_sc_hd__mux2_1 _29287_ (.A0(_09321_),
    .A1(\datamem.data_ram[62][29] ),
    .S(_13159_),
    .X(_13165_));
 sky130_fd_sc_hd__clkbuf_1 _29288_ (.A(_13165_),
    .X(_04412_));
 sky130_fd_sc_hd__mux2_1 _29289_ (.A0(_09325_),
    .A1(\datamem.data_ram[62][30] ),
    .S(_13159_),
    .X(_13166_));
 sky130_fd_sc_hd__clkbuf_1 _29290_ (.A(_13166_),
    .X(_04413_));
 sky130_fd_sc_hd__mux2_1 _29291_ (.A0(_09329_),
    .A1(\datamem.data_ram[62][31] ),
    .S(_13159_),
    .X(_13167_));
 sky130_fd_sc_hd__clkbuf_1 _29292_ (.A(_13167_),
    .X(_04414_));
 sky130_fd_sc_hd__dfxtp_1 _29293_ (.CLK(clk),
    .D(_01028_),
    .Q(\rvcpu.dp.plde.RD1E[0] ));
 sky130_fd_sc_hd__dfxtp_1 _29294_ (.CLK(clk),
    .D(_01029_),
    .Q(\rvcpu.dp.plde.RD1E[1] ));
 sky130_fd_sc_hd__dfxtp_1 _29295_ (.CLK(clk),
    .D(_01030_),
    .Q(\rvcpu.dp.plde.RD1E[2] ));
 sky130_fd_sc_hd__dfxtp_1 _29296_ (.CLK(clk),
    .D(_01031_),
    .Q(\rvcpu.dp.plde.RD1E[3] ));
 sky130_fd_sc_hd__dfxtp_1 _29297_ (.CLK(clk),
    .D(_01032_),
    .Q(\rvcpu.dp.plde.RD1E[4] ));
 sky130_fd_sc_hd__dfxtp_1 _29298_ (.CLK(clk),
    .D(_01033_),
    .Q(\rvcpu.dp.plde.RD1E[5] ));
 sky130_fd_sc_hd__dfxtp_1 _29299_ (.CLK(clk),
    .D(_01034_),
    .Q(\rvcpu.dp.plde.RD1E[6] ));
 sky130_fd_sc_hd__dfxtp_1 _29300_ (.CLK(clk),
    .D(_01035_),
    .Q(\rvcpu.dp.plde.RD1E[7] ));
 sky130_fd_sc_hd__dfxtp_1 _29301_ (.CLK(clk),
    .D(_01036_),
    .Q(\rvcpu.dp.plde.RD1E[8] ));
 sky130_fd_sc_hd__dfxtp_1 _29302_ (.CLK(clk),
    .D(_01037_),
    .Q(\rvcpu.dp.plde.RD1E[9] ));
 sky130_fd_sc_hd__dfxtp_1 _29303_ (.CLK(clk),
    .D(_01038_),
    .Q(\rvcpu.dp.plde.RD1E[10] ));
 sky130_fd_sc_hd__dfxtp_1 _29304_ (.CLK(clk),
    .D(_01039_),
    .Q(\rvcpu.dp.plde.RD1E[11] ));
 sky130_fd_sc_hd__dfxtp_1 _29305_ (.CLK(clk),
    .D(_01040_),
    .Q(\rvcpu.dp.plde.RD1E[12] ));
 sky130_fd_sc_hd__dfxtp_1 _29306_ (.CLK(clk),
    .D(_01041_),
    .Q(\rvcpu.dp.plde.RD1E[13] ));
 sky130_fd_sc_hd__dfxtp_1 _29307_ (.CLK(clk),
    .D(_01042_),
    .Q(\rvcpu.dp.plde.RD1E[14] ));
 sky130_fd_sc_hd__dfxtp_1 _29308_ (.CLK(clk),
    .D(_01043_),
    .Q(\rvcpu.dp.plde.RD1E[15] ));
 sky130_fd_sc_hd__dfxtp_1 _29309_ (.CLK(clk),
    .D(_01044_),
    .Q(\rvcpu.dp.plde.RD1E[16] ));
 sky130_fd_sc_hd__dfxtp_1 _29310_ (.CLK(clk),
    .D(_01045_),
    .Q(\rvcpu.dp.plde.RD1E[17] ));
 sky130_fd_sc_hd__dfxtp_1 _29311_ (.CLK(clk),
    .D(_01046_),
    .Q(\rvcpu.dp.plde.RD1E[18] ));
 sky130_fd_sc_hd__dfxtp_1 _29312_ (.CLK(clk),
    .D(_01047_),
    .Q(\rvcpu.dp.plde.RD1E[19] ));
 sky130_fd_sc_hd__dfxtp_1 _29313_ (.CLK(clk),
    .D(_01048_),
    .Q(\rvcpu.dp.plde.RD1E[20] ));
 sky130_fd_sc_hd__dfxtp_1 _29314_ (.CLK(clk),
    .D(_01049_),
    .Q(\rvcpu.dp.plde.RD1E[21] ));
 sky130_fd_sc_hd__dfxtp_1 _29315_ (.CLK(clk),
    .D(_01050_),
    .Q(\rvcpu.dp.plde.RD1E[22] ));
 sky130_fd_sc_hd__dfxtp_1 _29316_ (.CLK(clk),
    .D(_01051_),
    .Q(\rvcpu.dp.plde.RD1E[23] ));
 sky130_fd_sc_hd__dfxtp_1 _29317_ (.CLK(clk),
    .D(_01052_),
    .Q(\rvcpu.dp.plde.RD1E[24] ));
 sky130_fd_sc_hd__dfxtp_1 _29318_ (.CLK(clk),
    .D(_01053_),
    .Q(\rvcpu.dp.plde.RD1E[25] ));
 sky130_fd_sc_hd__dfxtp_1 _29319_ (.CLK(clk),
    .D(_01054_),
    .Q(\rvcpu.dp.plde.RD1E[26] ));
 sky130_fd_sc_hd__dfxtp_1 _29320_ (.CLK(clk),
    .D(_01055_),
    .Q(\rvcpu.dp.plde.RD1E[27] ));
 sky130_fd_sc_hd__dfxtp_1 _29321_ (.CLK(clk),
    .D(_01056_),
    .Q(\rvcpu.dp.plde.RD1E[28] ));
 sky130_fd_sc_hd__dfxtp_1 _29322_ (.CLK(clk),
    .D(_01057_),
    .Q(\rvcpu.dp.plde.RD1E[29] ));
 sky130_fd_sc_hd__dfxtp_1 _29323_ (.CLK(clk),
    .D(_01058_),
    .Q(\rvcpu.dp.plde.RD1E[30] ));
 sky130_fd_sc_hd__dfxtp_1 _29324_ (.CLK(clk),
    .D(_01059_),
    .Q(\rvcpu.dp.plde.RD1E[31] ));
 sky130_fd_sc_hd__dfxtp_1 _29325_ (.CLK(clk),
    .D(_01060_),
    .Q(\datamem.data_ram[62][16] ));
 sky130_fd_sc_hd__dfxtp_1 _29326_ (.CLK(clk),
    .D(_01061_),
    .Q(\datamem.data_ram[62][17] ));
 sky130_fd_sc_hd__dfxtp_1 _29327_ (.CLK(clk),
    .D(_01062_),
    .Q(\datamem.data_ram[62][18] ));
 sky130_fd_sc_hd__dfxtp_1 _29328_ (.CLK(clk),
    .D(_01063_),
    .Q(\datamem.data_ram[62][19] ));
 sky130_fd_sc_hd__dfxtp_1 _29329_ (.CLK(clk),
    .D(_01064_),
    .Q(\datamem.data_ram[62][20] ));
 sky130_fd_sc_hd__dfxtp_1 _29330_ (.CLK(clk),
    .D(_01065_),
    .Q(\datamem.data_ram[62][21] ));
 sky130_fd_sc_hd__dfxtp_1 _29331_ (.CLK(clk),
    .D(_01066_),
    .Q(\datamem.data_ram[62][22] ));
 sky130_fd_sc_hd__dfxtp_1 _29332_ (.CLK(clk),
    .D(_01067_),
    .Q(\datamem.data_ram[62][23] ));
 sky130_fd_sc_hd__dfxtp_1 _29333_ (.CLK(clk),
    .D(_01068_),
    .Q(\datamem.data_ram[62][8] ));
 sky130_fd_sc_hd__dfxtp_1 _29334_ (.CLK(clk),
    .D(_01069_),
    .Q(\datamem.data_ram[62][9] ));
 sky130_fd_sc_hd__dfxtp_1 _29335_ (.CLK(clk),
    .D(_01070_),
    .Q(\datamem.data_ram[62][10] ));
 sky130_fd_sc_hd__dfxtp_1 _29336_ (.CLK(clk),
    .D(_01071_),
    .Q(\datamem.data_ram[62][11] ));
 sky130_fd_sc_hd__dfxtp_1 _29337_ (.CLK(clk),
    .D(_01072_),
    .Q(\datamem.data_ram[62][12] ));
 sky130_fd_sc_hd__dfxtp_1 _29338_ (.CLK(clk),
    .D(_01073_),
    .Q(\datamem.data_ram[62][13] ));
 sky130_fd_sc_hd__dfxtp_1 _29339_ (.CLK(clk),
    .D(_01074_),
    .Q(\datamem.data_ram[62][14] ));
 sky130_fd_sc_hd__dfxtp_1 _29340_ (.CLK(clk),
    .D(_01075_),
    .Q(\datamem.data_ram[62][15] ));
 sky130_fd_sc_hd__dfxtp_1 _29341_ (.CLK(clk),
    .D(_01076_),
    .Q(\datamem.data_ram[61][24] ));
 sky130_fd_sc_hd__dfxtp_1 _29342_ (.CLK(clk),
    .D(_01077_),
    .Q(\datamem.data_ram[61][25] ));
 sky130_fd_sc_hd__dfxtp_1 _29343_ (.CLK(clk),
    .D(_01078_),
    .Q(\datamem.data_ram[61][26] ));
 sky130_fd_sc_hd__dfxtp_1 _29344_ (.CLK(clk),
    .D(_01079_),
    .Q(\datamem.data_ram[61][27] ));
 sky130_fd_sc_hd__dfxtp_1 _29345_ (.CLK(clk),
    .D(_01080_),
    .Q(\datamem.data_ram[61][28] ));
 sky130_fd_sc_hd__dfxtp_1 _29346_ (.CLK(clk),
    .D(_01081_),
    .Q(\datamem.data_ram[61][29] ));
 sky130_fd_sc_hd__dfxtp_1 _29347_ (.CLK(clk),
    .D(_01082_),
    .Q(\datamem.data_ram[61][30] ));
 sky130_fd_sc_hd__dfxtp_1 _29348_ (.CLK(clk),
    .D(_01083_),
    .Q(\datamem.data_ram[61][31] ));
 sky130_fd_sc_hd__dfxtp_1 _29349_ (.CLK(clk),
    .D(_01084_),
    .Q(\datamem.data_ram[61][16] ));
 sky130_fd_sc_hd__dfxtp_1 _29350_ (.CLK(clk),
    .D(_01085_),
    .Q(\datamem.data_ram[61][17] ));
 sky130_fd_sc_hd__dfxtp_1 _29351_ (.CLK(clk),
    .D(_01086_),
    .Q(\datamem.data_ram[61][18] ));
 sky130_fd_sc_hd__dfxtp_1 _29352_ (.CLK(clk),
    .D(_01087_),
    .Q(\datamem.data_ram[61][19] ));
 sky130_fd_sc_hd__dfxtp_1 _29353_ (.CLK(clk),
    .D(_01088_),
    .Q(\datamem.data_ram[61][20] ));
 sky130_fd_sc_hd__dfxtp_1 _29354_ (.CLK(clk),
    .D(_01089_),
    .Q(\datamem.data_ram[61][21] ));
 sky130_fd_sc_hd__dfxtp_1 _29355_ (.CLK(clk),
    .D(_01090_),
    .Q(\datamem.data_ram[61][22] ));
 sky130_fd_sc_hd__dfxtp_1 _29356_ (.CLK(clk),
    .D(_01091_),
    .Q(\datamem.data_ram[61][23] ));
 sky130_fd_sc_hd__dfxtp_1 _29357_ (.CLK(clk),
    .D(_01092_),
    .Q(\datamem.data_ram[61][8] ));
 sky130_fd_sc_hd__dfxtp_1 _29358_ (.CLK(clk),
    .D(_01093_),
    .Q(\datamem.data_ram[61][9] ));
 sky130_fd_sc_hd__dfxtp_1 _29359_ (.CLK(clk),
    .D(_01094_),
    .Q(\datamem.data_ram[61][10] ));
 sky130_fd_sc_hd__dfxtp_1 _29360_ (.CLK(clk),
    .D(_01095_),
    .Q(\datamem.data_ram[61][11] ));
 sky130_fd_sc_hd__dfxtp_1 _29361_ (.CLK(clk),
    .D(_01096_),
    .Q(\datamem.data_ram[61][12] ));
 sky130_fd_sc_hd__dfxtp_1 _29362_ (.CLK(clk),
    .D(_01097_),
    .Q(\datamem.data_ram[61][13] ));
 sky130_fd_sc_hd__dfxtp_1 _29363_ (.CLK(clk),
    .D(_01098_),
    .Q(\datamem.data_ram[61][14] ));
 sky130_fd_sc_hd__dfxtp_1 _29364_ (.CLK(clk),
    .D(_01099_),
    .Q(\datamem.data_ram[61][15] ));
 sky130_fd_sc_hd__dfxtp_1 _29365_ (.CLK(clk),
    .D(_01100_),
    .Q(\datamem.data_ram[60][24] ));
 sky130_fd_sc_hd__dfxtp_1 _29366_ (.CLK(clk),
    .D(_01101_),
    .Q(\datamem.data_ram[60][25] ));
 sky130_fd_sc_hd__dfxtp_1 _29367_ (.CLK(clk),
    .D(_01102_),
    .Q(\datamem.data_ram[60][26] ));
 sky130_fd_sc_hd__dfxtp_1 _29368_ (.CLK(clk),
    .D(_01103_),
    .Q(\datamem.data_ram[60][27] ));
 sky130_fd_sc_hd__dfxtp_1 _29369_ (.CLK(clk),
    .D(_01104_),
    .Q(\datamem.data_ram[60][28] ));
 sky130_fd_sc_hd__dfxtp_1 _29370_ (.CLK(clk),
    .D(_01105_),
    .Q(\datamem.data_ram[60][29] ));
 sky130_fd_sc_hd__dfxtp_1 _29371_ (.CLK(clk),
    .D(_01106_),
    .Q(\datamem.data_ram[60][30] ));
 sky130_fd_sc_hd__dfxtp_1 _29372_ (.CLK(clk),
    .D(_01107_),
    .Q(\datamem.data_ram[60][31] ));
 sky130_fd_sc_hd__dfxtp_1 _29373_ (.CLK(clk),
    .D(_01108_),
    .Q(\datamem.data_ram[60][16] ));
 sky130_fd_sc_hd__dfxtp_1 _29374_ (.CLK(clk),
    .D(_01109_),
    .Q(\datamem.data_ram[60][17] ));
 sky130_fd_sc_hd__dfxtp_1 _29375_ (.CLK(clk),
    .D(_01110_),
    .Q(\datamem.data_ram[60][18] ));
 sky130_fd_sc_hd__dfxtp_1 _29376_ (.CLK(clk),
    .D(_01111_),
    .Q(\datamem.data_ram[60][19] ));
 sky130_fd_sc_hd__dfxtp_1 _29377_ (.CLK(clk),
    .D(_01112_),
    .Q(\datamem.data_ram[60][20] ));
 sky130_fd_sc_hd__dfxtp_1 _29378_ (.CLK(clk),
    .D(_01113_),
    .Q(\datamem.data_ram[60][21] ));
 sky130_fd_sc_hd__dfxtp_1 _29379_ (.CLK(clk),
    .D(_01114_),
    .Q(\datamem.data_ram[60][22] ));
 sky130_fd_sc_hd__dfxtp_1 _29380_ (.CLK(clk),
    .D(_01115_),
    .Q(\datamem.data_ram[60][23] ));
 sky130_fd_sc_hd__dfxtp_1 _29381_ (.CLK(clk),
    .D(_01116_),
    .Q(\datamem.data_ram[60][8] ));
 sky130_fd_sc_hd__dfxtp_1 _29382_ (.CLK(clk),
    .D(_01117_),
    .Q(\datamem.data_ram[60][9] ));
 sky130_fd_sc_hd__dfxtp_1 _29383_ (.CLK(clk),
    .D(_01118_),
    .Q(\datamem.data_ram[60][10] ));
 sky130_fd_sc_hd__dfxtp_1 _29384_ (.CLK(clk),
    .D(_01119_),
    .Q(\datamem.data_ram[60][11] ));
 sky130_fd_sc_hd__dfxtp_1 _29385_ (.CLK(clk),
    .D(_01120_),
    .Q(\datamem.data_ram[60][12] ));
 sky130_fd_sc_hd__dfxtp_1 _29386_ (.CLK(clk),
    .D(_01121_),
    .Q(\datamem.data_ram[60][13] ));
 sky130_fd_sc_hd__dfxtp_1 _29387_ (.CLK(clk),
    .D(_01122_),
    .Q(\datamem.data_ram[60][14] ));
 sky130_fd_sc_hd__dfxtp_1 _29388_ (.CLK(clk),
    .D(_01123_),
    .Q(\datamem.data_ram[60][15] ));
 sky130_fd_sc_hd__dfxtp_1 _29389_ (.CLK(clk),
    .D(_01124_),
    .Q(\rvcpu.dp.plde.RD2E[0] ));
 sky130_fd_sc_hd__dfxtp_1 _29390_ (.CLK(clk),
    .D(_01125_),
    .Q(\rvcpu.dp.plde.RD2E[1] ));
 sky130_fd_sc_hd__dfxtp_1 _29391_ (.CLK(clk),
    .D(_01126_),
    .Q(\rvcpu.dp.plde.RD2E[2] ));
 sky130_fd_sc_hd__dfxtp_1 _29392_ (.CLK(clk),
    .D(_01127_),
    .Q(\rvcpu.dp.plde.RD2E[3] ));
 sky130_fd_sc_hd__dfxtp_1 _29393_ (.CLK(clk),
    .D(_01128_),
    .Q(\rvcpu.dp.plde.RD2E[4] ));
 sky130_fd_sc_hd__dfxtp_1 _29394_ (.CLK(clk),
    .D(_01129_),
    .Q(\rvcpu.dp.plde.RD2E[5] ));
 sky130_fd_sc_hd__dfxtp_1 _29395_ (.CLK(clk),
    .D(_01130_),
    .Q(\rvcpu.dp.plde.RD2E[6] ));
 sky130_fd_sc_hd__dfxtp_1 _29396_ (.CLK(clk),
    .D(_01131_),
    .Q(\rvcpu.dp.plde.RD2E[7] ));
 sky130_fd_sc_hd__dfxtp_1 _29397_ (.CLK(clk),
    .D(_01132_),
    .Q(\rvcpu.dp.plde.RD2E[8] ));
 sky130_fd_sc_hd__dfxtp_1 _29398_ (.CLK(clk),
    .D(_01133_),
    .Q(\rvcpu.dp.plde.RD2E[9] ));
 sky130_fd_sc_hd__dfxtp_1 _29399_ (.CLK(clk),
    .D(_01134_),
    .Q(\rvcpu.dp.plde.RD2E[10] ));
 sky130_fd_sc_hd__dfxtp_1 _29400_ (.CLK(clk),
    .D(_01135_),
    .Q(\rvcpu.dp.plde.RD2E[11] ));
 sky130_fd_sc_hd__dfxtp_1 _29401_ (.CLK(clk),
    .D(_01136_),
    .Q(\rvcpu.dp.plde.RD2E[12] ));
 sky130_fd_sc_hd__dfxtp_1 _29402_ (.CLK(clk),
    .D(_01137_),
    .Q(\rvcpu.dp.plde.RD2E[13] ));
 sky130_fd_sc_hd__dfxtp_1 _29403_ (.CLK(clk),
    .D(_01138_),
    .Q(\rvcpu.dp.plde.RD2E[14] ));
 sky130_fd_sc_hd__dfxtp_1 _29404_ (.CLK(clk),
    .D(_01139_),
    .Q(\rvcpu.dp.plde.RD2E[15] ));
 sky130_fd_sc_hd__dfxtp_1 _29405_ (.CLK(clk),
    .D(_01140_),
    .Q(\rvcpu.dp.plde.RD2E[16] ));
 sky130_fd_sc_hd__dfxtp_1 _29406_ (.CLK(clk),
    .D(_01141_),
    .Q(\rvcpu.dp.plde.RD2E[17] ));
 sky130_fd_sc_hd__dfxtp_1 _29407_ (.CLK(clk),
    .D(_01142_),
    .Q(\rvcpu.dp.plde.RD2E[18] ));
 sky130_fd_sc_hd__dfxtp_1 _29408_ (.CLK(clk),
    .D(_01143_),
    .Q(\rvcpu.dp.plde.RD2E[19] ));
 sky130_fd_sc_hd__dfxtp_1 _29409_ (.CLK(clk),
    .D(_01144_),
    .Q(\rvcpu.dp.plde.RD2E[20] ));
 sky130_fd_sc_hd__dfxtp_1 _29410_ (.CLK(clk),
    .D(_01145_),
    .Q(\rvcpu.dp.plde.RD2E[21] ));
 sky130_fd_sc_hd__dfxtp_1 _29411_ (.CLK(clk),
    .D(_01146_),
    .Q(\rvcpu.dp.plde.RD2E[22] ));
 sky130_fd_sc_hd__dfxtp_1 _29412_ (.CLK(clk),
    .D(_01147_),
    .Q(\rvcpu.dp.plde.RD2E[23] ));
 sky130_fd_sc_hd__dfxtp_1 _29413_ (.CLK(clk),
    .D(_01148_),
    .Q(\rvcpu.dp.plde.RD2E[24] ));
 sky130_fd_sc_hd__dfxtp_1 _29414_ (.CLK(clk),
    .D(_01149_),
    .Q(\rvcpu.dp.plde.RD2E[25] ));
 sky130_fd_sc_hd__dfxtp_1 _29415_ (.CLK(clk),
    .D(_01150_),
    .Q(\rvcpu.dp.plde.RD2E[26] ));
 sky130_fd_sc_hd__dfxtp_1 _29416_ (.CLK(clk),
    .D(_01151_),
    .Q(\rvcpu.dp.plde.RD2E[27] ));
 sky130_fd_sc_hd__dfxtp_1 _29417_ (.CLK(clk),
    .D(_01152_),
    .Q(\rvcpu.dp.plde.RD2E[28] ));
 sky130_fd_sc_hd__dfxtp_1 _29418_ (.CLK(clk),
    .D(_01153_),
    .Q(\rvcpu.dp.plde.RD2E[29] ));
 sky130_fd_sc_hd__dfxtp_1 _29419_ (.CLK(clk),
    .D(_01154_),
    .Q(\rvcpu.dp.plde.RD2E[30] ));
 sky130_fd_sc_hd__dfxtp_1 _29420_ (.CLK(clk),
    .D(_01155_),
    .Q(\rvcpu.dp.plde.RD2E[31] ));
 sky130_fd_sc_hd__dfxtp_1 _29421_ (.CLK(clk),
    .D(_01156_),
    .Q(\datamem.data_ram[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _29422_ (.CLK(clk),
    .D(_01157_),
    .Q(\datamem.data_ram[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _29423_ (.CLK(clk),
    .D(_01158_),
    .Q(\datamem.data_ram[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _29424_ (.CLK(clk),
    .D(_01159_),
    .Q(\datamem.data_ram[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _29425_ (.CLK(clk),
    .D(_01160_),
    .Q(\datamem.data_ram[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _29426_ (.CLK(clk),
    .D(_01161_),
    .Q(\datamem.data_ram[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _29427_ (.CLK(clk),
    .D(_01162_),
    .Q(\datamem.data_ram[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _29428_ (.CLK(clk),
    .D(_01163_),
    .Q(\datamem.data_ram[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _29429_ (.CLK(_00004_),
    .D(_01164_),
    .Q(\rvcpu.dp.rf.reg_file_arr[30][0] ));
 sky130_fd_sc_hd__dfxtp_1 _29430_ (.CLK(_00005_),
    .D(_01165_),
    .Q(\rvcpu.dp.rf.reg_file_arr[30][1] ));
 sky130_fd_sc_hd__dfxtp_1 _29431_ (.CLK(_00006_),
    .D(_01166_),
    .Q(\rvcpu.dp.rf.reg_file_arr[30][2] ));
 sky130_fd_sc_hd__dfxtp_1 _29432_ (.CLK(_00007_),
    .D(_01167_),
    .Q(\rvcpu.dp.rf.reg_file_arr[30][3] ));
 sky130_fd_sc_hd__dfxtp_1 _29433_ (.CLK(_00008_),
    .D(_01168_),
    .Q(\rvcpu.dp.rf.reg_file_arr[30][4] ));
 sky130_fd_sc_hd__dfxtp_1 _29434_ (.CLK(_00009_),
    .D(_01169_),
    .Q(\rvcpu.dp.rf.reg_file_arr[30][5] ));
 sky130_fd_sc_hd__dfxtp_1 _29435_ (.CLK(_00010_),
    .D(_01170_),
    .Q(\rvcpu.dp.rf.reg_file_arr[30][6] ));
 sky130_fd_sc_hd__dfxtp_1 _29436_ (.CLK(_00011_),
    .D(_01171_),
    .Q(\rvcpu.dp.rf.reg_file_arr[30][7] ));
 sky130_fd_sc_hd__dfxtp_1 _29437_ (.CLK(_00012_),
    .D(_01172_),
    .Q(\rvcpu.dp.rf.reg_file_arr[30][8] ));
 sky130_fd_sc_hd__dfxtp_1 _29438_ (.CLK(_00013_),
    .D(_01173_),
    .Q(\rvcpu.dp.rf.reg_file_arr[30][9] ));
 sky130_fd_sc_hd__dfxtp_1 _29439_ (.CLK(_00014_),
    .D(_01174_),
    .Q(\rvcpu.dp.rf.reg_file_arr[30][10] ));
 sky130_fd_sc_hd__dfxtp_1 _29440_ (.CLK(_00015_),
    .D(_01175_),
    .Q(\rvcpu.dp.rf.reg_file_arr[30][11] ));
 sky130_fd_sc_hd__dfxtp_1 _29441_ (.CLK(_00016_),
    .D(_01176_),
    .Q(\rvcpu.dp.rf.reg_file_arr[30][12] ));
 sky130_fd_sc_hd__dfxtp_1 _29442_ (.CLK(_00017_),
    .D(_01177_),
    .Q(\rvcpu.dp.rf.reg_file_arr[30][13] ));
 sky130_fd_sc_hd__dfxtp_1 _29443_ (.CLK(_00018_),
    .D(_01178_),
    .Q(\rvcpu.dp.rf.reg_file_arr[30][14] ));
 sky130_fd_sc_hd__dfxtp_1 _29444_ (.CLK(_00019_),
    .D(_01179_),
    .Q(\rvcpu.dp.rf.reg_file_arr[30][15] ));
 sky130_fd_sc_hd__dfxtp_1 _29445_ (.CLK(_00020_),
    .D(_01180_),
    .Q(\rvcpu.dp.rf.reg_file_arr[30][16] ));
 sky130_fd_sc_hd__dfxtp_1 _29446_ (.CLK(_00021_),
    .D(_01181_),
    .Q(\rvcpu.dp.rf.reg_file_arr[30][17] ));
 sky130_fd_sc_hd__dfxtp_1 _29447_ (.CLK(_00022_),
    .D(_01182_),
    .Q(\rvcpu.dp.rf.reg_file_arr[30][18] ));
 sky130_fd_sc_hd__dfxtp_1 _29448_ (.CLK(_00023_),
    .D(_01183_),
    .Q(\rvcpu.dp.rf.reg_file_arr[30][19] ));
 sky130_fd_sc_hd__dfxtp_1 _29449_ (.CLK(_00024_),
    .D(_01184_),
    .Q(\rvcpu.dp.rf.reg_file_arr[30][20] ));
 sky130_fd_sc_hd__dfxtp_1 _29450_ (.CLK(_00025_),
    .D(_01185_),
    .Q(\rvcpu.dp.rf.reg_file_arr[30][21] ));
 sky130_fd_sc_hd__dfxtp_1 _29451_ (.CLK(_00026_),
    .D(_01186_),
    .Q(\rvcpu.dp.rf.reg_file_arr[30][22] ));
 sky130_fd_sc_hd__dfxtp_1 _29452_ (.CLK(_00027_),
    .D(_01187_),
    .Q(\rvcpu.dp.rf.reg_file_arr[30][23] ));
 sky130_fd_sc_hd__dfxtp_1 _29453_ (.CLK(_00028_),
    .D(_01188_),
    .Q(\rvcpu.dp.rf.reg_file_arr[30][24] ));
 sky130_fd_sc_hd__dfxtp_1 _29454_ (.CLK(_00029_),
    .D(_01189_),
    .Q(\rvcpu.dp.rf.reg_file_arr[30][25] ));
 sky130_fd_sc_hd__dfxtp_1 _29455_ (.CLK(_00030_),
    .D(_01190_),
    .Q(\rvcpu.dp.rf.reg_file_arr[30][26] ));
 sky130_fd_sc_hd__dfxtp_1 _29456_ (.CLK(_00031_),
    .D(_01191_),
    .Q(\rvcpu.dp.rf.reg_file_arr[30][27] ));
 sky130_fd_sc_hd__dfxtp_1 _29457_ (.CLK(_00032_),
    .D(_01192_),
    .Q(\rvcpu.dp.rf.reg_file_arr[30][28] ));
 sky130_fd_sc_hd__dfxtp_1 _29458_ (.CLK(_00033_),
    .D(_01193_),
    .Q(\rvcpu.dp.rf.reg_file_arr[30][29] ));
 sky130_fd_sc_hd__dfxtp_1 _29459_ (.CLK(_00034_),
    .D(_01194_),
    .Q(\rvcpu.dp.rf.reg_file_arr[30][30] ));
 sky130_fd_sc_hd__dfxtp_1 _29460_ (.CLK(_00035_),
    .D(_01195_),
    .Q(\rvcpu.dp.rf.reg_file_arr[30][31] ));
 sky130_fd_sc_hd__dfxtp_1 _29461_ (.CLK(_00036_),
    .D(_01196_),
    .Q(\rvcpu.dp.rf.reg_file_arr[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _29462_ (.CLK(_00037_),
    .D(_01197_),
    .Q(\rvcpu.dp.rf.reg_file_arr[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _29463_ (.CLK(_00038_),
    .D(_01198_),
    .Q(\rvcpu.dp.rf.reg_file_arr[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _29464_ (.CLK(_00039_),
    .D(_01199_),
    .Q(\rvcpu.dp.rf.reg_file_arr[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _29465_ (.CLK(_00040_),
    .D(_01200_),
    .Q(\rvcpu.dp.rf.reg_file_arr[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _29466_ (.CLK(_00041_),
    .D(_01201_),
    .Q(\rvcpu.dp.rf.reg_file_arr[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _29467_ (.CLK(_00042_),
    .D(_01202_),
    .Q(\rvcpu.dp.rf.reg_file_arr[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _29468_ (.CLK(_00043_),
    .D(_01203_),
    .Q(\rvcpu.dp.rf.reg_file_arr[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _29469_ (.CLK(_00044_),
    .D(_01204_),
    .Q(\rvcpu.dp.rf.reg_file_arr[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _29470_ (.CLK(_00045_),
    .D(_01205_),
    .Q(\rvcpu.dp.rf.reg_file_arr[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _29471_ (.CLK(_00046_),
    .D(_01206_),
    .Q(\rvcpu.dp.rf.reg_file_arr[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _29472_ (.CLK(_00047_),
    .D(_01207_),
    .Q(\rvcpu.dp.rf.reg_file_arr[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _29473_ (.CLK(_00048_),
    .D(_01208_),
    .Q(\rvcpu.dp.rf.reg_file_arr[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _29474_ (.CLK(_00049_),
    .D(_01209_),
    .Q(\rvcpu.dp.rf.reg_file_arr[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _29475_ (.CLK(_00050_),
    .D(_01210_),
    .Q(\rvcpu.dp.rf.reg_file_arr[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _29476_ (.CLK(_00051_),
    .D(_01211_),
    .Q(\rvcpu.dp.rf.reg_file_arr[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _29477_ (.CLK(_00052_),
    .D(_01212_),
    .Q(\rvcpu.dp.rf.reg_file_arr[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _29478_ (.CLK(_00053_),
    .D(_01213_),
    .Q(\rvcpu.dp.rf.reg_file_arr[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _29479_ (.CLK(_00054_),
    .D(_01214_),
    .Q(\rvcpu.dp.rf.reg_file_arr[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _29480_ (.CLK(_00055_),
    .D(_01215_),
    .Q(\rvcpu.dp.rf.reg_file_arr[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _29481_ (.CLK(_00056_),
    .D(_01216_),
    .Q(\rvcpu.dp.rf.reg_file_arr[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _29482_ (.CLK(_00057_),
    .D(_01217_),
    .Q(\rvcpu.dp.rf.reg_file_arr[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _29483_ (.CLK(_00058_),
    .D(_01218_),
    .Q(\rvcpu.dp.rf.reg_file_arr[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _29484_ (.CLK(_00059_),
    .D(_01219_),
    .Q(\rvcpu.dp.rf.reg_file_arr[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _29485_ (.CLK(_00060_),
    .D(_01220_),
    .Q(\rvcpu.dp.rf.reg_file_arr[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _29486_ (.CLK(_00061_),
    .D(_01221_),
    .Q(\rvcpu.dp.rf.reg_file_arr[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _29487_ (.CLK(_00062_),
    .D(_01222_),
    .Q(\rvcpu.dp.rf.reg_file_arr[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _29488_ (.CLK(_00063_),
    .D(_01223_),
    .Q(\rvcpu.dp.rf.reg_file_arr[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _29489_ (.CLK(_00064_),
    .D(_01224_),
    .Q(\rvcpu.dp.rf.reg_file_arr[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _29490_ (.CLK(_00065_),
    .D(_01225_),
    .Q(\rvcpu.dp.rf.reg_file_arr[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _29491_ (.CLK(_00066_),
    .D(_01226_),
    .Q(\rvcpu.dp.rf.reg_file_arr[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _29492_ (.CLK(_00067_),
    .D(_01227_),
    .Q(\rvcpu.dp.rf.reg_file_arr[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _29493_ (.CLK(_00068_),
    .D(_01228_),
    .Q(\rvcpu.dp.rf.reg_file_arr[28][0] ));
 sky130_fd_sc_hd__dfxtp_1 _29494_ (.CLK(_00069_),
    .D(_01229_),
    .Q(\rvcpu.dp.rf.reg_file_arr[28][1] ));
 sky130_fd_sc_hd__dfxtp_1 _29495_ (.CLK(_00070_),
    .D(_01230_),
    .Q(\rvcpu.dp.rf.reg_file_arr[28][2] ));
 sky130_fd_sc_hd__dfxtp_1 _29496_ (.CLK(_00071_),
    .D(_01231_),
    .Q(\rvcpu.dp.rf.reg_file_arr[28][3] ));
 sky130_fd_sc_hd__dfxtp_1 _29497_ (.CLK(_00072_),
    .D(_01232_),
    .Q(\rvcpu.dp.rf.reg_file_arr[28][4] ));
 sky130_fd_sc_hd__dfxtp_1 _29498_ (.CLK(_00073_),
    .D(_01233_),
    .Q(\rvcpu.dp.rf.reg_file_arr[28][5] ));
 sky130_fd_sc_hd__dfxtp_1 _29499_ (.CLK(_00074_),
    .D(_01234_),
    .Q(\rvcpu.dp.rf.reg_file_arr[28][6] ));
 sky130_fd_sc_hd__dfxtp_1 _29500_ (.CLK(_00075_),
    .D(_01235_),
    .Q(\rvcpu.dp.rf.reg_file_arr[28][7] ));
 sky130_fd_sc_hd__dfxtp_1 _29501_ (.CLK(_00076_),
    .D(_01236_),
    .Q(\rvcpu.dp.rf.reg_file_arr[28][8] ));
 sky130_fd_sc_hd__dfxtp_1 _29502_ (.CLK(_00077_),
    .D(_01237_),
    .Q(\rvcpu.dp.rf.reg_file_arr[28][9] ));
 sky130_fd_sc_hd__dfxtp_1 _29503_ (.CLK(_00078_),
    .D(_01238_),
    .Q(\rvcpu.dp.rf.reg_file_arr[28][10] ));
 sky130_fd_sc_hd__dfxtp_1 _29504_ (.CLK(_00079_),
    .D(_01239_),
    .Q(\rvcpu.dp.rf.reg_file_arr[28][11] ));
 sky130_fd_sc_hd__dfxtp_1 _29505_ (.CLK(_00080_),
    .D(_01240_),
    .Q(\rvcpu.dp.rf.reg_file_arr[28][12] ));
 sky130_fd_sc_hd__dfxtp_1 _29506_ (.CLK(_00081_),
    .D(_01241_),
    .Q(\rvcpu.dp.rf.reg_file_arr[28][13] ));
 sky130_fd_sc_hd__dfxtp_1 _29507_ (.CLK(_00082_),
    .D(_01242_),
    .Q(\rvcpu.dp.rf.reg_file_arr[28][14] ));
 sky130_fd_sc_hd__dfxtp_1 _29508_ (.CLK(_00083_),
    .D(_01243_),
    .Q(\rvcpu.dp.rf.reg_file_arr[28][15] ));
 sky130_fd_sc_hd__dfxtp_1 _29509_ (.CLK(_00084_),
    .D(_01244_),
    .Q(\rvcpu.dp.rf.reg_file_arr[28][16] ));
 sky130_fd_sc_hd__dfxtp_1 _29510_ (.CLK(_00085_),
    .D(_01245_),
    .Q(\rvcpu.dp.rf.reg_file_arr[28][17] ));
 sky130_fd_sc_hd__dfxtp_1 _29511_ (.CLK(_00086_),
    .D(_01246_),
    .Q(\rvcpu.dp.rf.reg_file_arr[28][18] ));
 sky130_fd_sc_hd__dfxtp_1 _29512_ (.CLK(_00087_),
    .D(_01247_),
    .Q(\rvcpu.dp.rf.reg_file_arr[28][19] ));
 sky130_fd_sc_hd__dfxtp_1 _29513_ (.CLK(_00088_),
    .D(_01248_),
    .Q(\rvcpu.dp.rf.reg_file_arr[28][20] ));
 sky130_fd_sc_hd__dfxtp_1 _29514_ (.CLK(_00089_),
    .D(_01249_),
    .Q(\rvcpu.dp.rf.reg_file_arr[28][21] ));
 sky130_fd_sc_hd__dfxtp_1 _29515_ (.CLK(_00090_),
    .D(_01250_),
    .Q(\rvcpu.dp.rf.reg_file_arr[28][22] ));
 sky130_fd_sc_hd__dfxtp_1 _29516_ (.CLK(_00091_),
    .D(_01251_),
    .Q(\rvcpu.dp.rf.reg_file_arr[28][23] ));
 sky130_fd_sc_hd__dfxtp_1 _29517_ (.CLK(_00092_),
    .D(_01252_),
    .Q(\rvcpu.dp.rf.reg_file_arr[28][24] ));
 sky130_fd_sc_hd__dfxtp_1 _29518_ (.CLK(_00093_),
    .D(_01253_),
    .Q(\rvcpu.dp.rf.reg_file_arr[28][25] ));
 sky130_fd_sc_hd__dfxtp_1 _29519_ (.CLK(_00094_),
    .D(_01254_),
    .Q(\rvcpu.dp.rf.reg_file_arr[28][26] ));
 sky130_fd_sc_hd__dfxtp_1 _29520_ (.CLK(_00095_),
    .D(_01255_),
    .Q(\rvcpu.dp.rf.reg_file_arr[28][27] ));
 sky130_fd_sc_hd__dfxtp_1 _29521_ (.CLK(_00096_),
    .D(_01256_),
    .Q(\rvcpu.dp.rf.reg_file_arr[28][28] ));
 sky130_fd_sc_hd__dfxtp_1 _29522_ (.CLK(_00097_),
    .D(_01257_),
    .Q(\rvcpu.dp.rf.reg_file_arr[28][29] ));
 sky130_fd_sc_hd__dfxtp_1 _29523_ (.CLK(_00098_),
    .D(_01258_),
    .Q(\rvcpu.dp.rf.reg_file_arr[28][30] ));
 sky130_fd_sc_hd__dfxtp_1 _29524_ (.CLK(_00099_),
    .D(_01259_),
    .Q(\rvcpu.dp.rf.reg_file_arr[28][31] ));
 sky130_fd_sc_hd__dfxtp_1 _29525_ (.CLK(clk),
    .D(_01260_),
    .Q(\datamem.data_ram[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _29526_ (.CLK(clk),
    .D(_01261_),
    .Q(\datamem.data_ram[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _29527_ (.CLK(clk),
    .D(_01262_),
    .Q(\datamem.data_ram[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _29528_ (.CLK(clk),
    .D(_01263_),
    .Q(\datamem.data_ram[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _29529_ (.CLK(clk),
    .D(_01264_),
    .Q(\datamem.data_ram[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _29530_ (.CLK(clk),
    .D(_01265_),
    .Q(\datamem.data_ram[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _29531_ (.CLK(clk),
    .D(_01266_),
    .Q(\datamem.data_ram[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _29532_ (.CLK(clk),
    .D(_01267_),
    .Q(\datamem.data_ram[5][15] ));
 sky130_fd_sc_hd__dfxtp_1 _29533_ (.CLK(_00100_),
    .D(_01268_),
    .Q(\rvcpu.dp.rf.reg_file_arr[27][0] ));
 sky130_fd_sc_hd__dfxtp_1 _29534_ (.CLK(_00101_),
    .D(_01269_),
    .Q(\rvcpu.dp.rf.reg_file_arr[27][1] ));
 sky130_fd_sc_hd__dfxtp_1 _29535_ (.CLK(_00102_),
    .D(_01270_),
    .Q(\rvcpu.dp.rf.reg_file_arr[27][2] ));
 sky130_fd_sc_hd__dfxtp_1 _29536_ (.CLK(_00103_),
    .D(_01271_),
    .Q(\rvcpu.dp.rf.reg_file_arr[27][3] ));
 sky130_fd_sc_hd__dfxtp_1 _29537_ (.CLK(_00104_),
    .D(_01272_),
    .Q(\rvcpu.dp.rf.reg_file_arr[27][4] ));
 sky130_fd_sc_hd__dfxtp_1 _29538_ (.CLK(_00105_),
    .D(_01273_),
    .Q(\rvcpu.dp.rf.reg_file_arr[27][5] ));
 sky130_fd_sc_hd__dfxtp_1 _29539_ (.CLK(_00106_),
    .D(_01274_),
    .Q(\rvcpu.dp.rf.reg_file_arr[27][6] ));
 sky130_fd_sc_hd__dfxtp_1 _29540_ (.CLK(_00107_),
    .D(_01275_),
    .Q(\rvcpu.dp.rf.reg_file_arr[27][7] ));
 sky130_fd_sc_hd__dfxtp_1 _29541_ (.CLK(_00108_),
    .D(_01276_),
    .Q(\rvcpu.dp.rf.reg_file_arr[27][8] ));
 sky130_fd_sc_hd__dfxtp_1 _29542_ (.CLK(_00109_),
    .D(_01277_),
    .Q(\rvcpu.dp.rf.reg_file_arr[27][9] ));
 sky130_fd_sc_hd__dfxtp_1 _29543_ (.CLK(_00110_),
    .D(_01278_),
    .Q(\rvcpu.dp.rf.reg_file_arr[27][10] ));
 sky130_fd_sc_hd__dfxtp_1 _29544_ (.CLK(_00111_),
    .D(_01279_),
    .Q(\rvcpu.dp.rf.reg_file_arr[27][11] ));
 sky130_fd_sc_hd__dfxtp_1 _29545_ (.CLK(_00112_),
    .D(_01280_),
    .Q(\rvcpu.dp.rf.reg_file_arr[27][12] ));
 sky130_fd_sc_hd__dfxtp_1 _29546_ (.CLK(_00113_),
    .D(_01281_),
    .Q(\rvcpu.dp.rf.reg_file_arr[27][13] ));
 sky130_fd_sc_hd__dfxtp_1 _29547_ (.CLK(_00114_),
    .D(_01282_),
    .Q(\rvcpu.dp.rf.reg_file_arr[27][14] ));
 sky130_fd_sc_hd__dfxtp_1 _29548_ (.CLK(_00115_),
    .D(_01283_),
    .Q(\rvcpu.dp.rf.reg_file_arr[27][15] ));
 sky130_fd_sc_hd__dfxtp_1 _29549_ (.CLK(_00116_),
    .D(_01284_),
    .Q(\rvcpu.dp.rf.reg_file_arr[27][16] ));
 sky130_fd_sc_hd__dfxtp_1 _29550_ (.CLK(_00117_),
    .D(_01285_),
    .Q(\rvcpu.dp.rf.reg_file_arr[27][17] ));
 sky130_fd_sc_hd__dfxtp_1 _29551_ (.CLK(_00118_),
    .D(_01286_),
    .Q(\rvcpu.dp.rf.reg_file_arr[27][18] ));
 sky130_fd_sc_hd__dfxtp_1 _29552_ (.CLK(_00119_),
    .D(_01287_),
    .Q(\rvcpu.dp.rf.reg_file_arr[27][19] ));
 sky130_fd_sc_hd__dfxtp_1 _29553_ (.CLK(_00120_),
    .D(_01288_),
    .Q(\rvcpu.dp.rf.reg_file_arr[27][20] ));
 sky130_fd_sc_hd__dfxtp_1 _29554_ (.CLK(_00121_),
    .D(_01289_),
    .Q(\rvcpu.dp.rf.reg_file_arr[27][21] ));
 sky130_fd_sc_hd__dfxtp_1 _29555_ (.CLK(_00122_),
    .D(_01290_),
    .Q(\rvcpu.dp.rf.reg_file_arr[27][22] ));
 sky130_fd_sc_hd__dfxtp_1 _29556_ (.CLK(_00123_),
    .D(_01291_),
    .Q(\rvcpu.dp.rf.reg_file_arr[27][23] ));
 sky130_fd_sc_hd__dfxtp_1 _29557_ (.CLK(_00124_),
    .D(_01292_),
    .Q(\rvcpu.dp.rf.reg_file_arr[27][24] ));
 sky130_fd_sc_hd__dfxtp_1 _29558_ (.CLK(_00125_),
    .D(_01293_),
    .Q(\rvcpu.dp.rf.reg_file_arr[27][25] ));
 sky130_fd_sc_hd__dfxtp_1 _29559_ (.CLK(_00126_),
    .D(_01294_),
    .Q(\rvcpu.dp.rf.reg_file_arr[27][26] ));
 sky130_fd_sc_hd__dfxtp_1 _29560_ (.CLK(_00127_),
    .D(_01295_),
    .Q(\rvcpu.dp.rf.reg_file_arr[27][27] ));
 sky130_fd_sc_hd__dfxtp_1 _29561_ (.CLK(_00128_),
    .D(_01296_),
    .Q(\rvcpu.dp.rf.reg_file_arr[27][28] ));
 sky130_fd_sc_hd__dfxtp_1 _29562_ (.CLK(_00129_),
    .D(_01297_),
    .Q(\rvcpu.dp.rf.reg_file_arr[27][29] ));
 sky130_fd_sc_hd__dfxtp_1 _29563_ (.CLK(_00130_),
    .D(_01298_),
    .Q(\rvcpu.dp.rf.reg_file_arr[27][30] ));
 sky130_fd_sc_hd__dfxtp_1 _29564_ (.CLK(_00131_),
    .D(_01299_),
    .Q(\rvcpu.dp.rf.reg_file_arr[27][31] ));
 sky130_fd_sc_hd__dfxtp_1 _29565_ (.CLK(_00132_),
    .D(_01300_),
    .Q(\rvcpu.dp.rf.reg_file_arr[26][0] ));
 sky130_fd_sc_hd__dfxtp_1 _29566_ (.CLK(_00133_),
    .D(_01301_),
    .Q(\rvcpu.dp.rf.reg_file_arr[26][1] ));
 sky130_fd_sc_hd__dfxtp_1 _29567_ (.CLK(_00134_),
    .D(_01302_),
    .Q(\rvcpu.dp.rf.reg_file_arr[26][2] ));
 sky130_fd_sc_hd__dfxtp_1 _29568_ (.CLK(_00135_),
    .D(_01303_),
    .Q(\rvcpu.dp.rf.reg_file_arr[26][3] ));
 sky130_fd_sc_hd__dfxtp_1 _29569_ (.CLK(_00136_),
    .D(_01304_),
    .Q(\rvcpu.dp.rf.reg_file_arr[26][4] ));
 sky130_fd_sc_hd__dfxtp_1 _29570_ (.CLK(_00137_),
    .D(_01305_),
    .Q(\rvcpu.dp.rf.reg_file_arr[26][5] ));
 sky130_fd_sc_hd__dfxtp_1 _29571_ (.CLK(_00138_),
    .D(_01306_),
    .Q(\rvcpu.dp.rf.reg_file_arr[26][6] ));
 sky130_fd_sc_hd__dfxtp_1 _29572_ (.CLK(_00139_),
    .D(_01307_),
    .Q(\rvcpu.dp.rf.reg_file_arr[26][7] ));
 sky130_fd_sc_hd__dfxtp_1 _29573_ (.CLK(_00140_),
    .D(_01308_),
    .Q(\rvcpu.dp.rf.reg_file_arr[26][8] ));
 sky130_fd_sc_hd__dfxtp_1 _29574_ (.CLK(_00141_),
    .D(_01309_),
    .Q(\rvcpu.dp.rf.reg_file_arr[26][9] ));
 sky130_fd_sc_hd__dfxtp_1 _29575_ (.CLK(_00142_),
    .D(_01310_),
    .Q(\rvcpu.dp.rf.reg_file_arr[26][10] ));
 sky130_fd_sc_hd__dfxtp_1 _29576_ (.CLK(_00143_),
    .D(_01311_),
    .Q(\rvcpu.dp.rf.reg_file_arr[26][11] ));
 sky130_fd_sc_hd__dfxtp_1 _29577_ (.CLK(_00144_),
    .D(_01312_),
    .Q(\rvcpu.dp.rf.reg_file_arr[26][12] ));
 sky130_fd_sc_hd__dfxtp_1 _29578_ (.CLK(_00145_),
    .D(_01313_),
    .Q(\rvcpu.dp.rf.reg_file_arr[26][13] ));
 sky130_fd_sc_hd__dfxtp_1 _29579_ (.CLK(_00146_),
    .D(_01314_),
    .Q(\rvcpu.dp.rf.reg_file_arr[26][14] ));
 sky130_fd_sc_hd__dfxtp_1 _29580_ (.CLK(_00147_),
    .D(_01315_),
    .Q(\rvcpu.dp.rf.reg_file_arr[26][15] ));
 sky130_fd_sc_hd__dfxtp_1 _29581_ (.CLK(_00148_),
    .D(_01316_),
    .Q(\rvcpu.dp.rf.reg_file_arr[26][16] ));
 sky130_fd_sc_hd__dfxtp_1 _29582_ (.CLK(_00149_),
    .D(_01317_),
    .Q(\rvcpu.dp.rf.reg_file_arr[26][17] ));
 sky130_fd_sc_hd__dfxtp_1 _29583_ (.CLK(_00150_),
    .D(_01318_),
    .Q(\rvcpu.dp.rf.reg_file_arr[26][18] ));
 sky130_fd_sc_hd__dfxtp_1 _29584_ (.CLK(_00151_),
    .D(_01319_),
    .Q(\rvcpu.dp.rf.reg_file_arr[26][19] ));
 sky130_fd_sc_hd__dfxtp_1 _29585_ (.CLK(_00152_),
    .D(_01320_),
    .Q(\rvcpu.dp.rf.reg_file_arr[26][20] ));
 sky130_fd_sc_hd__dfxtp_1 _29586_ (.CLK(_00153_),
    .D(_01321_),
    .Q(\rvcpu.dp.rf.reg_file_arr[26][21] ));
 sky130_fd_sc_hd__dfxtp_1 _29587_ (.CLK(_00154_),
    .D(_01322_),
    .Q(\rvcpu.dp.rf.reg_file_arr[26][22] ));
 sky130_fd_sc_hd__dfxtp_1 _29588_ (.CLK(_00155_),
    .D(_01323_),
    .Q(\rvcpu.dp.rf.reg_file_arr[26][23] ));
 sky130_fd_sc_hd__dfxtp_1 _29589_ (.CLK(_00156_),
    .D(_01324_),
    .Q(\rvcpu.dp.rf.reg_file_arr[26][24] ));
 sky130_fd_sc_hd__dfxtp_1 _29590_ (.CLK(_00157_),
    .D(_01325_),
    .Q(\rvcpu.dp.rf.reg_file_arr[26][25] ));
 sky130_fd_sc_hd__dfxtp_1 _29591_ (.CLK(_00158_),
    .D(_01326_),
    .Q(\rvcpu.dp.rf.reg_file_arr[26][26] ));
 sky130_fd_sc_hd__dfxtp_1 _29592_ (.CLK(_00159_),
    .D(_01327_),
    .Q(\rvcpu.dp.rf.reg_file_arr[26][27] ));
 sky130_fd_sc_hd__dfxtp_1 _29593_ (.CLK(_00160_),
    .D(_01328_),
    .Q(\rvcpu.dp.rf.reg_file_arr[26][28] ));
 sky130_fd_sc_hd__dfxtp_1 _29594_ (.CLK(_00161_),
    .D(_01329_),
    .Q(\rvcpu.dp.rf.reg_file_arr[26][29] ));
 sky130_fd_sc_hd__dfxtp_1 _29595_ (.CLK(_00162_),
    .D(_01330_),
    .Q(\rvcpu.dp.rf.reg_file_arr[26][30] ));
 sky130_fd_sc_hd__dfxtp_1 _29596_ (.CLK(_00163_),
    .D(_01331_),
    .Q(\rvcpu.dp.rf.reg_file_arr[26][31] ));
 sky130_fd_sc_hd__dfxtp_1 _29597_ (.CLK(_00164_),
    .D(_01332_),
    .Q(\rvcpu.dp.rf.reg_file_arr[25][0] ));
 sky130_fd_sc_hd__dfxtp_1 _29598_ (.CLK(_00165_),
    .D(_01333_),
    .Q(\rvcpu.dp.rf.reg_file_arr[25][1] ));
 sky130_fd_sc_hd__dfxtp_1 _29599_ (.CLK(_00166_),
    .D(_01334_),
    .Q(\rvcpu.dp.rf.reg_file_arr[25][2] ));
 sky130_fd_sc_hd__dfxtp_1 _29600_ (.CLK(_00167_),
    .D(_01335_),
    .Q(\rvcpu.dp.rf.reg_file_arr[25][3] ));
 sky130_fd_sc_hd__dfxtp_1 _29601_ (.CLK(_00168_),
    .D(_01336_),
    .Q(\rvcpu.dp.rf.reg_file_arr[25][4] ));
 sky130_fd_sc_hd__dfxtp_1 _29602_ (.CLK(_00169_),
    .D(_01337_),
    .Q(\rvcpu.dp.rf.reg_file_arr[25][5] ));
 sky130_fd_sc_hd__dfxtp_1 _29603_ (.CLK(_00170_),
    .D(_01338_),
    .Q(\rvcpu.dp.rf.reg_file_arr[25][6] ));
 sky130_fd_sc_hd__dfxtp_1 _29604_ (.CLK(_00171_),
    .D(_01339_),
    .Q(\rvcpu.dp.rf.reg_file_arr[25][7] ));
 sky130_fd_sc_hd__dfxtp_1 _29605_ (.CLK(_00172_),
    .D(_01340_),
    .Q(\rvcpu.dp.rf.reg_file_arr[25][8] ));
 sky130_fd_sc_hd__dfxtp_1 _29606_ (.CLK(_00173_),
    .D(_01341_),
    .Q(\rvcpu.dp.rf.reg_file_arr[25][9] ));
 sky130_fd_sc_hd__dfxtp_1 _29607_ (.CLK(_00174_),
    .D(_01342_),
    .Q(\rvcpu.dp.rf.reg_file_arr[25][10] ));
 sky130_fd_sc_hd__dfxtp_1 _29608_ (.CLK(_00175_),
    .D(_01343_),
    .Q(\rvcpu.dp.rf.reg_file_arr[25][11] ));
 sky130_fd_sc_hd__dfxtp_1 _29609_ (.CLK(_00176_),
    .D(_01344_),
    .Q(\rvcpu.dp.rf.reg_file_arr[25][12] ));
 sky130_fd_sc_hd__dfxtp_1 _29610_ (.CLK(_00177_),
    .D(_01345_),
    .Q(\rvcpu.dp.rf.reg_file_arr[25][13] ));
 sky130_fd_sc_hd__dfxtp_1 _29611_ (.CLK(_00178_),
    .D(_01346_),
    .Q(\rvcpu.dp.rf.reg_file_arr[25][14] ));
 sky130_fd_sc_hd__dfxtp_1 _29612_ (.CLK(_00179_),
    .D(_01347_),
    .Q(\rvcpu.dp.rf.reg_file_arr[25][15] ));
 sky130_fd_sc_hd__dfxtp_1 _29613_ (.CLK(_00180_),
    .D(_01348_),
    .Q(\rvcpu.dp.rf.reg_file_arr[25][16] ));
 sky130_fd_sc_hd__dfxtp_1 _29614_ (.CLK(_00181_),
    .D(_01349_),
    .Q(\rvcpu.dp.rf.reg_file_arr[25][17] ));
 sky130_fd_sc_hd__dfxtp_1 _29615_ (.CLK(_00182_),
    .D(_01350_),
    .Q(\rvcpu.dp.rf.reg_file_arr[25][18] ));
 sky130_fd_sc_hd__dfxtp_1 _29616_ (.CLK(_00183_),
    .D(_01351_),
    .Q(\rvcpu.dp.rf.reg_file_arr[25][19] ));
 sky130_fd_sc_hd__dfxtp_1 _29617_ (.CLK(_00184_),
    .D(_01352_),
    .Q(\rvcpu.dp.rf.reg_file_arr[25][20] ));
 sky130_fd_sc_hd__dfxtp_1 _29618_ (.CLK(_00185_),
    .D(_01353_),
    .Q(\rvcpu.dp.rf.reg_file_arr[25][21] ));
 sky130_fd_sc_hd__dfxtp_1 _29619_ (.CLK(_00186_),
    .D(_01354_),
    .Q(\rvcpu.dp.rf.reg_file_arr[25][22] ));
 sky130_fd_sc_hd__dfxtp_1 _29620_ (.CLK(_00187_),
    .D(_01355_),
    .Q(\rvcpu.dp.rf.reg_file_arr[25][23] ));
 sky130_fd_sc_hd__dfxtp_1 _29621_ (.CLK(_00188_),
    .D(_01356_),
    .Q(\rvcpu.dp.rf.reg_file_arr[25][24] ));
 sky130_fd_sc_hd__dfxtp_1 _29622_ (.CLK(_00189_),
    .D(_01357_),
    .Q(\rvcpu.dp.rf.reg_file_arr[25][25] ));
 sky130_fd_sc_hd__dfxtp_1 _29623_ (.CLK(_00190_),
    .D(_01358_),
    .Q(\rvcpu.dp.rf.reg_file_arr[25][26] ));
 sky130_fd_sc_hd__dfxtp_1 _29624_ (.CLK(_00191_),
    .D(_01359_),
    .Q(\rvcpu.dp.rf.reg_file_arr[25][27] ));
 sky130_fd_sc_hd__dfxtp_1 _29625_ (.CLK(_00192_),
    .D(_01360_),
    .Q(\rvcpu.dp.rf.reg_file_arr[25][28] ));
 sky130_fd_sc_hd__dfxtp_1 _29626_ (.CLK(_00193_),
    .D(_01361_),
    .Q(\rvcpu.dp.rf.reg_file_arr[25][29] ));
 sky130_fd_sc_hd__dfxtp_1 _29627_ (.CLK(_00194_),
    .D(_01362_),
    .Q(\rvcpu.dp.rf.reg_file_arr[25][30] ));
 sky130_fd_sc_hd__dfxtp_1 _29628_ (.CLK(_00195_),
    .D(_01363_),
    .Q(\rvcpu.dp.rf.reg_file_arr[25][31] ));
 sky130_fd_sc_hd__dfxtp_1 _29629_ (.CLK(clk),
    .D(_01364_),
    .Q(\datamem.data_ram[5][16] ));
 sky130_fd_sc_hd__dfxtp_1 _29630_ (.CLK(clk),
    .D(_01365_),
    .Q(\datamem.data_ram[5][17] ));
 sky130_fd_sc_hd__dfxtp_1 _29631_ (.CLK(clk),
    .D(_01366_),
    .Q(\datamem.data_ram[5][18] ));
 sky130_fd_sc_hd__dfxtp_1 _29632_ (.CLK(clk),
    .D(_01367_),
    .Q(\datamem.data_ram[5][19] ));
 sky130_fd_sc_hd__dfxtp_1 _29633_ (.CLK(clk),
    .D(_01368_),
    .Q(\datamem.data_ram[5][20] ));
 sky130_fd_sc_hd__dfxtp_1 _29634_ (.CLK(clk),
    .D(_01369_),
    .Q(\datamem.data_ram[5][21] ));
 sky130_fd_sc_hd__dfxtp_1 _29635_ (.CLK(clk),
    .D(_01370_),
    .Q(\datamem.data_ram[5][22] ));
 sky130_fd_sc_hd__dfxtp_1 _29636_ (.CLK(clk),
    .D(_01371_),
    .Q(\datamem.data_ram[5][23] ));
 sky130_fd_sc_hd__dfxtp_1 _29637_ (.CLK(_00196_),
    .D(_01372_),
    .Q(\rvcpu.dp.rf.reg_file_arr[24][0] ));
 sky130_fd_sc_hd__dfxtp_1 _29638_ (.CLK(_00197_),
    .D(_01373_),
    .Q(\rvcpu.dp.rf.reg_file_arr[24][1] ));
 sky130_fd_sc_hd__dfxtp_1 _29639_ (.CLK(_00198_),
    .D(_01374_),
    .Q(\rvcpu.dp.rf.reg_file_arr[24][2] ));
 sky130_fd_sc_hd__dfxtp_1 _29640_ (.CLK(_00199_),
    .D(_01375_),
    .Q(\rvcpu.dp.rf.reg_file_arr[24][3] ));
 sky130_fd_sc_hd__dfxtp_1 _29641_ (.CLK(_00200_),
    .D(_01376_),
    .Q(\rvcpu.dp.rf.reg_file_arr[24][4] ));
 sky130_fd_sc_hd__dfxtp_1 _29642_ (.CLK(_00201_),
    .D(_01377_),
    .Q(\rvcpu.dp.rf.reg_file_arr[24][5] ));
 sky130_fd_sc_hd__dfxtp_1 _29643_ (.CLK(_00202_),
    .D(_01378_),
    .Q(\rvcpu.dp.rf.reg_file_arr[24][6] ));
 sky130_fd_sc_hd__dfxtp_1 _29644_ (.CLK(_00203_),
    .D(_01379_),
    .Q(\rvcpu.dp.rf.reg_file_arr[24][7] ));
 sky130_fd_sc_hd__dfxtp_1 _29645_ (.CLK(_00204_),
    .D(_01380_),
    .Q(\rvcpu.dp.rf.reg_file_arr[24][8] ));
 sky130_fd_sc_hd__dfxtp_1 _29646_ (.CLK(_00205_),
    .D(_01381_),
    .Q(\rvcpu.dp.rf.reg_file_arr[24][9] ));
 sky130_fd_sc_hd__dfxtp_1 _29647_ (.CLK(_00206_),
    .D(_01382_),
    .Q(\rvcpu.dp.rf.reg_file_arr[24][10] ));
 sky130_fd_sc_hd__dfxtp_1 _29648_ (.CLK(_00207_),
    .D(_01383_),
    .Q(\rvcpu.dp.rf.reg_file_arr[24][11] ));
 sky130_fd_sc_hd__dfxtp_1 _29649_ (.CLK(_00208_),
    .D(_01384_),
    .Q(\rvcpu.dp.rf.reg_file_arr[24][12] ));
 sky130_fd_sc_hd__dfxtp_1 _29650_ (.CLK(_00209_),
    .D(_01385_),
    .Q(\rvcpu.dp.rf.reg_file_arr[24][13] ));
 sky130_fd_sc_hd__dfxtp_1 _29651_ (.CLK(_00210_),
    .D(_01386_),
    .Q(\rvcpu.dp.rf.reg_file_arr[24][14] ));
 sky130_fd_sc_hd__dfxtp_1 _29652_ (.CLK(_00211_),
    .D(_01387_),
    .Q(\rvcpu.dp.rf.reg_file_arr[24][15] ));
 sky130_fd_sc_hd__dfxtp_1 _29653_ (.CLK(_00212_),
    .D(_01388_),
    .Q(\rvcpu.dp.rf.reg_file_arr[24][16] ));
 sky130_fd_sc_hd__dfxtp_1 _29654_ (.CLK(_00213_),
    .D(_01389_),
    .Q(\rvcpu.dp.rf.reg_file_arr[24][17] ));
 sky130_fd_sc_hd__dfxtp_1 _29655_ (.CLK(_00214_),
    .D(_01390_),
    .Q(\rvcpu.dp.rf.reg_file_arr[24][18] ));
 sky130_fd_sc_hd__dfxtp_1 _29656_ (.CLK(_00215_),
    .D(_01391_),
    .Q(\rvcpu.dp.rf.reg_file_arr[24][19] ));
 sky130_fd_sc_hd__dfxtp_1 _29657_ (.CLK(_00216_),
    .D(_01392_),
    .Q(\rvcpu.dp.rf.reg_file_arr[24][20] ));
 sky130_fd_sc_hd__dfxtp_1 _29658_ (.CLK(_00217_),
    .D(_01393_),
    .Q(\rvcpu.dp.rf.reg_file_arr[24][21] ));
 sky130_fd_sc_hd__dfxtp_1 _29659_ (.CLK(_00218_),
    .D(_01394_),
    .Q(\rvcpu.dp.rf.reg_file_arr[24][22] ));
 sky130_fd_sc_hd__dfxtp_1 _29660_ (.CLK(_00219_),
    .D(_01395_),
    .Q(\rvcpu.dp.rf.reg_file_arr[24][23] ));
 sky130_fd_sc_hd__dfxtp_1 _29661_ (.CLK(_00220_),
    .D(_01396_),
    .Q(\rvcpu.dp.rf.reg_file_arr[24][24] ));
 sky130_fd_sc_hd__dfxtp_1 _29662_ (.CLK(_00221_),
    .D(_01397_),
    .Q(\rvcpu.dp.rf.reg_file_arr[24][25] ));
 sky130_fd_sc_hd__dfxtp_1 _29663_ (.CLK(_00222_),
    .D(_01398_),
    .Q(\rvcpu.dp.rf.reg_file_arr[24][26] ));
 sky130_fd_sc_hd__dfxtp_1 _29664_ (.CLK(_00223_),
    .D(_01399_),
    .Q(\rvcpu.dp.rf.reg_file_arr[24][27] ));
 sky130_fd_sc_hd__dfxtp_1 _29665_ (.CLK(_00224_),
    .D(_01400_),
    .Q(\rvcpu.dp.rf.reg_file_arr[24][28] ));
 sky130_fd_sc_hd__dfxtp_1 _29666_ (.CLK(_00225_),
    .D(_01401_),
    .Q(\rvcpu.dp.rf.reg_file_arr[24][29] ));
 sky130_fd_sc_hd__dfxtp_1 _29667_ (.CLK(_00226_),
    .D(_01402_),
    .Q(\rvcpu.dp.rf.reg_file_arr[24][30] ));
 sky130_fd_sc_hd__dfxtp_1 _29668_ (.CLK(_00227_),
    .D(_01403_),
    .Q(\rvcpu.dp.rf.reg_file_arr[24][31] ));
 sky130_fd_sc_hd__dfxtp_1 _29669_ (.CLK(_00228_),
    .D(_01404_),
    .Q(\rvcpu.dp.rf.reg_file_arr[23][0] ));
 sky130_fd_sc_hd__dfxtp_1 _29670_ (.CLK(_00229_),
    .D(_01405_),
    .Q(\rvcpu.dp.rf.reg_file_arr[23][1] ));
 sky130_fd_sc_hd__dfxtp_1 _29671_ (.CLK(_00230_),
    .D(_01406_),
    .Q(\rvcpu.dp.rf.reg_file_arr[23][2] ));
 sky130_fd_sc_hd__dfxtp_1 _29672_ (.CLK(_00231_),
    .D(_01407_),
    .Q(\rvcpu.dp.rf.reg_file_arr[23][3] ));
 sky130_fd_sc_hd__dfxtp_1 _29673_ (.CLK(_00232_),
    .D(_01408_),
    .Q(\rvcpu.dp.rf.reg_file_arr[23][4] ));
 sky130_fd_sc_hd__dfxtp_1 _29674_ (.CLK(_00233_),
    .D(_01409_),
    .Q(\rvcpu.dp.rf.reg_file_arr[23][5] ));
 sky130_fd_sc_hd__dfxtp_1 _29675_ (.CLK(_00234_),
    .D(_01410_),
    .Q(\rvcpu.dp.rf.reg_file_arr[23][6] ));
 sky130_fd_sc_hd__dfxtp_1 _29676_ (.CLK(_00235_),
    .D(_01411_),
    .Q(\rvcpu.dp.rf.reg_file_arr[23][7] ));
 sky130_fd_sc_hd__dfxtp_1 _29677_ (.CLK(_00236_),
    .D(_01412_),
    .Q(\rvcpu.dp.rf.reg_file_arr[23][8] ));
 sky130_fd_sc_hd__dfxtp_1 _29678_ (.CLK(_00237_),
    .D(_01413_),
    .Q(\rvcpu.dp.rf.reg_file_arr[23][9] ));
 sky130_fd_sc_hd__dfxtp_1 _29679_ (.CLK(_00238_),
    .D(_01414_),
    .Q(\rvcpu.dp.rf.reg_file_arr[23][10] ));
 sky130_fd_sc_hd__dfxtp_1 _29680_ (.CLK(_00239_),
    .D(_01415_),
    .Q(\rvcpu.dp.rf.reg_file_arr[23][11] ));
 sky130_fd_sc_hd__dfxtp_1 _29681_ (.CLK(_00240_),
    .D(_01416_),
    .Q(\rvcpu.dp.rf.reg_file_arr[23][12] ));
 sky130_fd_sc_hd__dfxtp_1 _29682_ (.CLK(_00241_),
    .D(_01417_),
    .Q(\rvcpu.dp.rf.reg_file_arr[23][13] ));
 sky130_fd_sc_hd__dfxtp_1 _29683_ (.CLK(_00242_),
    .D(_01418_),
    .Q(\rvcpu.dp.rf.reg_file_arr[23][14] ));
 sky130_fd_sc_hd__dfxtp_1 _29684_ (.CLK(_00243_),
    .D(_01419_),
    .Q(\rvcpu.dp.rf.reg_file_arr[23][15] ));
 sky130_fd_sc_hd__dfxtp_1 _29685_ (.CLK(_00244_),
    .D(_01420_),
    .Q(\rvcpu.dp.rf.reg_file_arr[23][16] ));
 sky130_fd_sc_hd__dfxtp_1 _29686_ (.CLK(_00245_),
    .D(_01421_),
    .Q(\rvcpu.dp.rf.reg_file_arr[23][17] ));
 sky130_fd_sc_hd__dfxtp_1 _29687_ (.CLK(_00246_),
    .D(_01422_),
    .Q(\rvcpu.dp.rf.reg_file_arr[23][18] ));
 sky130_fd_sc_hd__dfxtp_1 _29688_ (.CLK(_00247_),
    .D(_01423_),
    .Q(\rvcpu.dp.rf.reg_file_arr[23][19] ));
 sky130_fd_sc_hd__dfxtp_1 _29689_ (.CLK(_00248_),
    .D(_01424_),
    .Q(\rvcpu.dp.rf.reg_file_arr[23][20] ));
 sky130_fd_sc_hd__dfxtp_1 _29690_ (.CLK(_00249_),
    .D(_01425_),
    .Q(\rvcpu.dp.rf.reg_file_arr[23][21] ));
 sky130_fd_sc_hd__dfxtp_1 _29691_ (.CLK(_00250_),
    .D(_01426_),
    .Q(\rvcpu.dp.rf.reg_file_arr[23][22] ));
 sky130_fd_sc_hd__dfxtp_1 _29692_ (.CLK(_00251_),
    .D(_01427_),
    .Q(\rvcpu.dp.rf.reg_file_arr[23][23] ));
 sky130_fd_sc_hd__dfxtp_1 _29693_ (.CLK(_00252_),
    .D(_01428_),
    .Q(\rvcpu.dp.rf.reg_file_arr[23][24] ));
 sky130_fd_sc_hd__dfxtp_1 _29694_ (.CLK(_00253_),
    .D(_01429_),
    .Q(\rvcpu.dp.rf.reg_file_arr[23][25] ));
 sky130_fd_sc_hd__dfxtp_1 _29695_ (.CLK(_00254_),
    .D(_01430_),
    .Q(\rvcpu.dp.rf.reg_file_arr[23][26] ));
 sky130_fd_sc_hd__dfxtp_1 _29696_ (.CLK(_00255_),
    .D(_01431_),
    .Q(\rvcpu.dp.rf.reg_file_arr[23][27] ));
 sky130_fd_sc_hd__dfxtp_1 _29697_ (.CLK(_00256_),
    .D(_01432_),
    .Q(\rvcpu.dp.rf.reg_file_arr[23][28] ));
 sky130_fd_sc_hd__dfxtp_1 _29698_ (.CLK(_00257_),
    .D(_01433_),
    .Q(\rvcpu.dp.rf.reg_file_arr[23][29] ));
 sky130_fd_sc_hd__dfxtp_1 _29699_ (.CLK(_00258_),
    .D(_01434_),
    .Q(\rvcpu.dp.rf.reg_file_arr[23][30] ));
 sky130_fd_sc_hd__dfxtp_1 _29700_ (.CLK(_00259_),
    .D(_01435_),
    .Q(\rvcpu.dp.rf.reg_file_arr[23][31] ));
 sky130_fd_sc_hd__dfxtp_1 _29701_ (.CLK(_00260_),
    .D(_01436_),
    .Q(\rvcpu.dp.rf.reg_file_arr[22][0] ));
 sky130_fd_sc_hd__dfxtp_1 _29702_ (.CLK(_00261_),
    .D(_01437_),
    .Q(\rvcpu.dp.rf.reg_file_arr[22][1] ));
 sky130_fd_sc_hd__dfxtp_1 _29703_ (.CLK(_00262_),
    .D(_01438_),
    .Q(\rvcpu.dp.rf.reg_file_arr[22][2] ));
 sky130_fd_sc_hd__dfxtp_1 _29704_ (.CLK(_00263_),
    .D(_01439_),
    .Q(\rvcpu.dp.rf.reg_file_arr[22][3] ));
 sky130_fd_sc_hd__dfxtp_1 _29705_ (.CLK(_00264_),
    .D(_01440_),
    .Q(\rvcpu.dp.rf.reg_file_arr[22][4] ));
 sky130_fd_sc_hd__dfxtp_1 _29706_ (.CLK(_00265_),
    .D(_01441_),
    .Q(\rvcpu.dp.rf.reg_file_arr[22][5] ));
 sky130_fd_sc_hd__dfxtp_1 _29707_ (.CLK(_00266_),
    .D(_01442_),
    .Q(\rvcpu.dp.rf.reg_file_arr[22][6] ));
 sky130_fd_sc_hd__dfxtp_1 _29708_ (.CLK(_00267_),
    .D(_01443_),
    .Q(\rvcpu.dp.rf.reg_file_arr[22][7] ));
 sky130_fd_sc_hd__dfxtp_1 _29709_ (.CLK(_00268_),
    .D(_01444_),
    .Q(\rvcpu.dp.rf.reg_file_arr[22][8] ));
 sky130_fd_sc_hd__dfxtp_1 _29710_ (.CLK(_00269_),
    .D(_01445_),
    .Q(\rvcpu.dp.rf.reg_file_arr[22][9] ));
 sky130_fd_sc_hd__dfxtp_1 _29711_ (.CLK(_00270_),
    .D(_01446_),
    .Q(\rvcpu.dp.rf.reg_file_arr[22][10] ));
 sky130_fd_sc_hd__dfxtp_1 _29712_ (.CLK(_00271_),
    .D(_01447_),
    .Q(\rvcpu.dp.rf.reg_file_arr[22][11] ));
 sky130_fd_sc_hd__dfxtp_1 _29713_ (.CLK(_00272_),
    .D(_01448_),
    .Q(\rvcpu.dp.rf.reg_file_arr[22][12] ));
 sky130_fd_sc_hd__dfxtp_1 _29714_ (.CLK(_00273_),
    .D(_01449_),
    .Q(\rvcpu.dp.rf.reg_file_arr[22][13] ));
 sky130_fd_sc_hd__dfxtp_1 _29715_ (.CLK(_00274_),
    .D(_01450_),
    .Q(\rvcpu.dp.rf.reg_file_arr[22][14] ));
 sky130_fd_sc_hd__dfxtp_1 _29716_ (.CLK(_00275_),
    .D(_01451_),
    .Q(\rvcpu.dp.rf.reg_file_arr[22][15] ));
 sky130_fd_sc_hd__dfxtp_1 _29717_ (.CLK(_00276_),
    .D(_01452_),
    .Q(\rvcpu.dp.rf.reg_file_arr[22][16] ));
 sky130_fd_sc_hd__dfxtp_1 _29718_ (.CLK(_00277_),
    .D(_01453_),
    .Q(\rvcpu.dp.rf.reg_file_arr[22][17] ));
 sky130_fd_sc_hd__dfxtp_1 _29719_ (.CLK(_00278_),
    .D(_01454_),
    .Q(\rvcpu.dp.rf.reg_file_arr[22][18] ));
 sky130_fd_sc_hd__dfxtp_1 _29720_ (.CLK(_00279_),
    .D(_01455_),
    .Q(\rvcpu.dp.rf.reg_file_arr[22][19] ));
 sky130_fd_sc_hd__dfxtp_1 _29721_ (.CLK(_00280_),
    .D(_01456_),
    .Q(\rvcpu.dp.rf.reg_file_arr[22][20] ));
 sky130_fd_sc_hd__dfxtp_1 _29722_ (.CLK(_00281_),
    .D(_01457_),
    .Q(\rvcpu.dp.rf.reg_file_arr[22][21] ));
 sky130_fd_sc_hd__dfxtp_1 _29723_ (.CLK(_00282_),
    .D(_01458_),
    .Q(\rvcpu.dp.rf.reg_file_arr[22][22] ));
 sky130_fd_sc_hd__dfxtp_1 _29724_ (.CLK(_00283_),
    .D(_01459_),
    .Q(\rvcpu.dp.rf.reg_file_arr[22][23] ));
 sky130_fd_sc_hd__dfxtp_1 _29725_ (.CLK(_00284_),
    .D(_01460_),
    .Q(\rvcpu.dp.rf.reg_file_arr[22][24] ));
 sky130_fd_sc_hd__dfxtp_1 _29726_ (.CLK(_00285_),
    .D(_01461_),
    .Q(\rvcpu.dp.rf.reg_file_arr[22][25] ));
 sky130_fd_sc_hd__dfxtp_1 _29727_ (.CLK(_00286_),
    .D(_01462_),
    .Q(\rvcpu.dp.rf.reg_file_arr[22][26] ));
 sky130_fd_sc_hd__dfxtp_1 _29728_ (.CLK(_00287_),
    .D(_01463_),
    .Q(\rvcpu.dp.rf.reg_file_arr[22][27] ));
 sky130_fd_sc_hd__dfxtp_1 _29729_ (.CLK(_00288_),
    .D(_01464_),
    .Q(\rvcpu.dp.rf.reg_file_arr[22][28] ));
 sky130_fd_sc_hd__dfxtp_1 _29730_ (.CLK(_00289_),
    .D(_01465_),
    .Q(\rvcpu.dp.rf.reg_file_arr[22][29] ));
 sky130_fd_sc_hd__dfxtp_1 _29731_ (.CLK(_00290_),
    .D(_01466_),
    .Q(\rvcpu.dp.rf.reg_file_arr[22][30] ));
 sky130_fd_sc_hd__dfxtp_1 _29732_ (.CLK(_00291_),
    .D(_01467_),
    .Q(\rvcpu.dp.rf.reg_file_arr[22][31] ));
 sky130_fd_sc_hd__dfxtp_1 _29733_ (.CLK(_00292_),
    .D(_01468_),
    .Q(\rvcpu.dp.rf.reg_file_arr[21][0] ));
 sky130_fd_sc_hd__dfxtp_1 _29734_ (.CLK(_00293_),
    .D(_01469_),
    .Q(\rvcpu.dp.rf.reg_file_arr[21][1] ));
 sky130_fd_sc_hd__dfxtp_1 _29735_ (.CLK(_00294_),
    .D(_01470_),
    .Q(\rvcpu.dp.rf.reg_file_arr[21][2] ));
 sky130_fd_sc_hd__dfxtp_1 _29736_ (.CLK(_00295_),
    .D(_01471_),
    .Q(\rvcpu.dp.rf.reg_file_arr[21][3] ));
 sky130_fd_sc_hd__dfxtp_1 _29737_ (.CLK(_00296_),
    .D(_01472_),
    .Q(\rvcpu.dp.rf.reg_file_arr[21][4] ));
 sky130_fd_sc_hd__dfxtp_1 _29738_ (.CLK(_00297_),
    .D(_01473_),
    .Q(\rvcpu.dp.rf.reg_file_arr[21][5] ));
 sky130_fd_sc_hd__dfxtp_1 _29739_ (.CLK(_00298_),
    .D(_01474_),
    .Q(\rvcpu.dp.rf.reg_file_arr[21][6] ));
 sky130_fd_sc_hd__dfxtp_1 _29740_ (.CLK(_00299_),
    .D(_01475_),
    .Q(\rvcpu.dp.rf.reg_file_arr[21][7] ));
 sky130_fd_sc_hd__dfxtp_1 _29741_ (.CLK(_00300_),
    .D(_01476_),
    .Q(\rvcpu.dp.rf.reg_file_arr[21][8] ));
 sky130_fd_sc_hd__dfxtp_1 _29742_ (.CLK(_00301_),
    .D(_01477_),
    .Q(\rvcpu.dp.rf.reg_file_arr[21][9] ));
 sky130_fd_sc_hd__dfxtp_1 _29743_ (.CLK(_00302_),
    .D(_01478_),
    .Q(\rvcpu.dp.rf.reg_file_arr[21][10] ));
 sky130_fd_sc_hd__dfxtp_1 _29744_ (.CLK(_00303_),
    .D(_01479_),
    .Q(\rvcpu.dp.rf.reg_file_arr[21][11] ));
 sky130_fd_sc_hd__dfxtp_1 _29745_ (.CLK(_00304_),
    .D(_01480_),
    .Q(\rvcpu.dp.rf.reg_file_arr[21][12] ));
 sky130_fd_sc_hd__dfxtp_1 _29746_ (.CLK(_00305_),
    .D(_01481_),
    .Q(\rvcpu.dp.rf.reg_file_arr[21][13] ));
 sky130_fd_sc_hd__dfxtp_1 _29747_ (.CLK(_00306_),
    .D(_01482_),
    .Q(\rvcpu.dp.rf.reg_file_arr[21][14] ));
 sky130_fd_sc_hd__dfxtp_1 _29748_ (.CLK(_00307_),
    .D(_01483_),
    .Q(\rvcpu.dp.rf.reg_file_arr[21][15] ));
 sky130_fd_sc_hd__dfxtp_1 _29749_ (.CLK(_00308_),
    .D(_01484_),
    .Q(\rvcpu.dp.rf.reg_file_arr[21][16] ));
 sky130_fd_sc_hd__dfxtp_1 _29750_ (.CLK(_00309_),
    .D(_01485_),
    .Q(\rvcpu.dp.rf.reg_file_arr[21][17] ));
 sky130_fd_sc_hd__dfxtp_1 _29751_ (.CLK(_00310_),
    .D(_01486_),
    .Q(\rvcpu.dp.rf.reg_file_arr[21][18] ));
 sky130_fd_sc_hd__dfxtp_1 _29752_ (.CLK(_00311_),
    .D(_01487_),
    .Q(\rvcpu.dp.rf.reg_file_arr[21][19] ));
 sky130_fd_sc_hd__dfxtp_1 _29753_ (.CLK(_00312_),
    .D(_01488_),
    .Q(\rvcpu.dp.rf.reg_file_arr[21][20] ));
 sky130_fd_sc_hd__dfxtp_1 _29754_ (.CLK(_00313_),
    .D(_01489_),
    .Q(\rvcpu.dp.rf.reg_file_arr[21][21] ));
 sky130_fd_sc_hd__dfxtp_1 _29755_ (.CLK(_00314_),
    .D(_01490_),
    .Q(\rvcpu.dp.rf.reg_file_arr[21][22] ));
 sky130_fd_sc_hd__dfxtp_1 _29756_ (.CLK(_00315_),
    .D(_01491_),
    .Q(\rvcpu.dp.rf.reg_file_arr[21][23] ));
 sky130_fd_sc_hd__dfxtp_1 _29757_ (.CLK(_00316_),
    .D(_01492_),
    .Q(\rvcpu.dp.rf.reg_file_arr[21][24] ));
 sky130_fd_sc_hd__dfxtp_1 _29758_ (.CLK(_00317_),
    .D(_01493_),
    .Q(\rvcpu.dp.rf.reg_file_arr[21][25] ));
 sky130_fd_sc_hd__dfxtp_1 _29759_ (.CLK(_00318_),
    .D(_01494_),
    .Q(\rvcpu.dp.rf.reg_file_arr[21][26] ));
 sky130_fd_sc_hd__dfxtp_1 _29760_ (.CLK(_00319_),
    .D(_01495_),
    .Q(\rvcpu.dp.rf.reg_file_arr[21][27] ));
 sky130_fd_sc_hd__dfxtp_1 _29761_ (.CLK(_00320_),
    .D(_01496_),
    .Q(\rvcpu.dp.rf.reg_file_arr[21][28] ));
 sky130_fd_sc_hd__dfxtp_1 _29762_ (.CLK(_00321_),
    .D(_01497_),
    .Q(\rvcpu.dp.rf.reg_file_arr[21][29] ));
 sky130_fd_sc_hd__dfxtp_1 _29763_ (.CLK(_00322_),
    .D(_01498_),
    .Q(\rvcpu.dp.rf.reg_file_arr[21][30] ));
 sky130_fd_sc_hd__dfxtp_1 _29764_ (.CLK(_00323_),
    .D(_01499_),
    .Q(\rvcpu.dp.rf.reg_file_arr[21][31] ));
 sky130_fd_sc_hd__dfxtp_1 _29765_ (.CLK(_00324_),
    .D(_01500_),
    .Q(\rvcpu.dp.rf.reg_file_arr[20][0] ));
 sky130_fd_sc_hd__dfxtp_1 _29766_ (.CLK(_00325_),
    .D(_01501_),
    .Q(\rvcpu.dp.rf.reg_file_arr[20][1] ));
 sky130_fd_sc_hd__dfxtp_1 _29767_ (.CLK(_00326_),
    .D(_01502_),
    .Q(\rvcpu.dp.rf.reg_file_arr[20][2] ));
 sky130_fd_sc_hd__dfxtp_1 _29768_ (.CLK(_00327_),
    .D(_01503_),
    .Q(\rvcpu.dp.rf.reg_file_arr[20][3] ));
 sky130_fd_sc_hd__dfxtp_1 _29769_ (.CLK(_00328_),
    .D(_01504_),
    .Q(\rvcpu.dp.rf.reg_file_arr[20][4] ));
 sky130_fd_sc_hd__dfxtp_1 _29770_ (.CLK(_00329_),
    .D(_01505_),
    .Q(\rvcpu.dp.rf.reg_file_arr[20][5] ));
 sky130_fd_sc_hd__dfxtp_1 _29771_ (.CLK(_00330_),
    .D(_01506_),
    .Q(\rvcpu.dp.rf.reg_file_arr[20][6] ));
 sky130_fd_sc_hd__dfxtp_1 _29772_ (.CLK(_00331_),
    .D(_01507_),
    .Q(\rvcpu.dp.rf.reg_file_arr[20][7] ));
 sky130_fd_sc_hd__dfxtp_1 _29773_ (.CLK(_00332_),
    .D(_01508_),
    .Q(\rvcpu.dp.rf.reg_file_arr[20][8] ));
 sky130_fd_sc_hd__dfxtp_1 _29774_ (.CLK(_00333_),
    .D(_01509_),
    .Q(\rvcpu.dp.rf.reg_file_arr[20][9] ));
 sky130_fd_sc_hd__dfxtp_1 _29775_ (.CLK(_00334_),
    .D(_01510_),
    .Q(\rvcpu.dp.rf.reg_file_arr[20][10] ));
 sky130_fd_sc_hd__dfxtp_1 _29776_ (.CLK(_00335_),
    .D(_01511_),
    .Q(\rvcpu.dp.rf.reg_file_arr[20][11] ));
 sky130_fd_sc_hd__dfxtp_1 _29777_ (.CLK(_00336_),
    .D(_01512_),
    .Q(\rvcpu.dp.rf.reg_file_arr[20][12] ));
 sky130_fd_sc_hd__dfxtp_1 _29778_ (.CLK(_00337_),
    .D(_01513_),
    .Q(\rvcpu.dp.rf.reg_file_arr[20][13] ));
 sky130_fd_sc_hd__dfxtp_1 _29779_ (.CLK(_00338_),
    .D(_01514_),
    .Q(\rvcpu.dp.rf.reg_file_arr[20][14] ));
 sky130_fd_sc_hd__dfxtp_1 _29780_ (.CLK(_00339_),
    .D(_01515_),
    .Q(\rvcpu.dp.rf.reg_file_arr[20][15] ));
 sky130_fd_sc_hd__dfxtp_1 _29781_ (.CLK(_00340_),
    .D(_01516_),
    .Q(\rvcpu.dp.rf.reg_file_arr[20][16] ));
 sky130_fd_sc_hd__dfxtp_1 _29782_ (.CLK(_00341_),
    .D(_01517_),
    .Q(\rvcpu.dp.rf.reg_file_arr[20][17] ));
 sky130_fd_sc_hd__dfxtp_1 _29783_ (.CLK(_00342_),
    .D(_01518_),
    .Q(\rvcpu.dp.rf.reg_file_arr[20][18] ));
 sky130_fd_sc_hd__dfxtp_1 _29784_ (.CLK(_00343_),
    .D(_01519_),
    .Q(\rvcpu.dp.rf.reg_file_arr[20][19] ));
 sky130_fd_sc_hd__dfxtp_1 _29785_ (.CLK(_00344_),
    .D(_01520_),
    .Q(\rvcpu.dp.rf.reg_file_arr[20][20] ));
 sky130_fd_sc_hd__dfxtp_1 _29786_ (.CLK(_00345_),
    .D(_01521_),
    .Q(\rvcpu.dp.rf.reg_file_arr[20][21] ));
 sky130_fd_sc_hd__dfxtp_1 _29787_ (.CLK(_00346_),
    .D(_01522_),
    .Q(\rvcpu.dp.rf.reg_file_arr[20][22] ));
 sky130_fd_sc_hd__dfxtp_1 _29788_ (.CLK(_00347_),
    .D(_01523_),
    .Q(\rvcpu.dp.rf.reg_file_arr[20][23] ));
 sky130_fd_sc_hd__dfxtp_1 _29789_ (.CLK(_00348_),
    .D(_01524_),
    .Q(\rvcpu.dp.rf.reg_file_arr[20][24] ));
 sky130_fd_sc_hd__dfxtp_1 _29790_ (.CLK(_00349_),
    .D(_01525_),
    .Q(\rvcpu.dp.rf.reg_file_arr[20][25] ));
 sky130_fd_sc_hd__dfxtp_1 _29791_ (.CLK(_00350_),
    .D(_01526_),
    .Q(\rvcpu.dp.rf.reg_file_arr[20][26] ));
 sky130_fd_sc_hd__dfxtp_1 _29792_ (.CLK(_00351_),
    .D(_01527_),
    .Q(\rvcpu.dp.rf.reg_file_arr[20][27] ));
 sky130_fd_sc_hd__dfxtp_1 _29793_ (.CLK(_00352_),
    .D(_01528_),
    .Q(\rvcpu.dp.rf.reg_file_arr[20][28] ));
 sky130_fd_sc_hd__dfxtp_1 _29794_ (.CLK(_00353_),
    .D(_01529_),
    .Q(\rvcpu.dp.rf.reg_file_arr[20][29] ));
 sky130_fd_sc_hd__dfxtp_1 _29795_ (.CLK(_00354_),
    .D(_01530_),
    .Q(\rvcpu.dp.rf.reg_file_arr[20][30] ));
 sky130_fd_sc_hd__dfxtp_1 _29796_ (.CLK(_00355_),
    .D(_01531_),
    .Q(\rvcpu.dp.rf.reg_file_arr[20][31] ));
 sky130_fd_sc_hd__dfxtp_1 _29797_ (.CLK(clk),
    .D(_01532_),
    .Q(\datamem.data_ram[59][24] ));
 sky130_fd_sc_hd__dfxtp_1 _29798_ (.CLK(clk),
    .D(_01533_),
    .Q(\datamem.data_ram[59][25] ));
 sky130_fd_sc_hd__dfxtp_1 _29799_ (.CLK(clk),
    .D(_01534_),
    .Q(\datamem.data_ram[59][26] ));
 sky130_fd_sc_hd__dfxtp_1 _29800_ (.CLK(clk),
    .D(_01535_),
    .Q(\datamem.data_ram[59][27] ));
 sky130_fd_sc_hd__dfxtp_1 _29801_ (.CLK(clk),
    .D(_01536_),
    .Q(\datamem.data_ram[59][28] ));
 sky130_fd_sc_hd__dfxtp_1 _29802_ (.CLK(clk),
    .D(_01537_),
    .Q(\datamem.data_ram[59][29] ));
 sky130_fd_sc_hd__dfxtp_1 _29803_ (.CLK(clk),
    .D(_01538_),
    .Q(\datamem.data_ram[59][30] ));
 sky130_fd_sc_hd__dfxtp_1 _29804_ (.CLK(clk),
    .D(_01539_),
    .Q(\datamem.data_ram[59][31] ));
 sky130_fd_sc_hd__dfxtp_1 _29805_ (.CLK(_00356_),
    .D(_01540_),
    .Q(\rvcpu.dp.rf.reg_file_arr[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _29806_ (.CLK(_00357_),
    .D(_01541_),
    .Q(\rvcpu.dp.rf.reg_file_arr[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _29807_ (.CLK(_00358_),
    .D(_01542_),
    .Q(\rvcpu.dp.rf.reg_file_arr[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _29808_ (.CLK(_00359_),
    .D(_01543_),
    .Q(\rvcpu.dp.rf.reg_file_arr[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _29809_ (.CLK(_00360_),
    .D(_01544_),
    .Q(\rvcpu.dp.rf.reg_file_arr[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _29810_ (.CLK(_00361_),
    .D(_01545_),
    .Q(\rvcpu.dp.rf.reg_file_arr[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _29811_ (.CLK(_00362_),
    .D(_01546_),
    .Q(\rvcpu.dp.rf.reg_file_arr[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _29812_ (.CLK(_00363_),
    .D(_01547_),
    .Q(\rvcpu.dp.rf.reg_file_arr[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _29813_ (.CLK(_00364_),
    .D(_01548_),
    .Q(\rvcpu.dp.rf.reg_file_arr[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _29814_ (.CLK(_00365_),
    .D(_01549_),
    .Q(\rvcpu.dp.rf.reg_file_arr[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _29815_ (.CLK(_00366_),
    .D(_01550_),
    .Q(\rvcpu.dp.rf.reg_file_arr[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _29816_ (.CLK(_00367_),
    .D(_01551_),
    .Q(\rvcpu.dp.rf.reg_file_arr[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _29817_ (.CLK(_00368_),
    .D(_01552_),
    .Q(\rvcpu.dp.rf.reg_file_arr[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _29818_ (.CLK(_00369_),
    .D(_01553_),
    .Q(\rvcpu.dp.rf.reg_file_arr[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _29819_ (.CLK(_00370_),
    .D(_01554_),
    .Q(\rvcpu.dp.rf.reg_file_arr[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _29820_ (.CLK(_00371_),
    .D(_01555_),
    .Q(\rvcpu.dp.rf.reg_file_arr[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _29821_ (.CLK(_00372_),
    .D(_01556_),
    .Q(\rvcpu.dp.rf.reg_file_arr[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _29822_ (.CLK(_00373_),
    .D(_01557_),
    .Q(\rvcpu.dp.rf.reg_file_arr[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _29823_ (.CLK(_00374_),
    .D(_01558_),
    .Q(\rvcpu.dp.rf.reg_file_arr[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _29824_ (.CLK(_00375_),
    .D(_01559_),
    .Q(\rvcpu.dp.rf.reg_file_arr[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _29825_ (.CLK(_00376_),
    .D(_01560_),
    .Q(\rvcpu.dp.rf.reg_file_arr[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _29826_ (.CLK(_00377_),
    .D(_01561_),
    .Q(\rvcpu.dp.rf.reg_file_arr[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _29827_ (.CLK(_00378_),
    .D(_01562_),
    .Q(\rvcpu.dp.rf.reg_file_arr[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _29828_ (.CLK(_00379_),
    .D(_01563_),
    .Q(\rvcpu.dp.rf.reg_file_arr[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _29829_ (.CLK(_00380_),
    .D(_01564_),
    .Q(\rvcpu.dp.rf.reg_file_arr[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _29830_ (.CLK(_00381_),
    .D(_01565_),
    .Q(\rvcpu.dp.rf.reg_file_arr[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _29831_ (.CLK(_00382_),
    .D(_01566_),
    .Q(\rvcpu.dp.rf.reg_file_arr[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _29832_ (.CLK(_00383_),
    .D(_01567_),
    .Q(\rvcpu.dp.rf.reg_file_arr[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _29833_ (.CLK(_00384_),
    .D(_01568_),
    .Q(\rvcpu.dp.rf.reg_file_arr[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _29834_ (.CLK(_00385_),
    .D(_01569_),
    .Q(\rvcpu.dp.rf.reg_file_arr[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _29835_ (.CLK(_00386_),
    .D(_01570_),
    .Q(\rvcpu.dp.rf.reg_file_arr[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _29836_ (.CLK(_00387_),
    .D(_01571_),
    .Q(\rvcpu.dp.rf.reg_file_arr[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _29837_ (.CLK(_00388_),
    .D(_01572_),
    .Q(\rvcpu.dp.rf.reg_file_arr[18][0] ));
 sky130_fd_sc_hd__dfxtp_1 _29838_ (.CLK(_00389_),
    .D(_01573_),
    .Q(\rvcpu.dp.rf.reg_file_arr[18][1] ));
 sky130_fd_sc_hd__dfxtp_1 _29839_ (.CLK(_00390_),
    .D(_01574_),
    .Q(\rvcpu.dp.rf.reg_file_arr[18][2] ));
 sky130_fd_sc_hd__dfxtp_1 _29840_ (.CLK(_00391_),
    .D(_01575_),
    .Q(\rvcpu.dp.rf.reg_file_arr[18][3] ));
 sky130_fd_sc_hd__dfxtp_1 _29841_ (.CLK(_00392_),
    .D(_01576_),
    .Q(\rvcpu.dp.rf.reg_file_arr[18][4] ));
 sky130_fd_sc_hd__dfxtp_1 _29842_ (.CLK(_00393_),
    .D(_01577_),
    .Q(\rvcpu.dp.rf.reg_file_arr[18][5] ));
 sky130_fd_sc_hd__dfxtp_1 _29843_ (.CLK(_00394_),
    .D(_01578_),
    .Q(\rvcpu.dp.rf.reg_file_arr[18][6] ));
 sky130_fd_sc_hd__dfxtp_1 _29844_ (.CLK(_00395_),
    .D(_01579_),
    .Q(\rvcpu.dp.rf.reg_file_arr[18][7] ));
 sky130_fd_sc_hd__dfxtp_1 _29845_ (.CLK(_00396_),
    .D(_01580_),
    .Q(\rvcpu.dp.rf.reg_file_arr[18][8] ));
 sky130_fd_sc_hd__dfxtp_1 _29846_ (.CLK(_00397_),
    .D(_01581_),
    .Q(\rvcpu.dp.rf.reg_file_arr[18][9] ));
 sky130_fd_sc_hd__dfxtp_1 _29847_ (.CLK(_00398_),
    .D(_01582_),
    .Q(\rvcpu.dp.rf.reg_file_arr[18][10] ));
 sky130_fd_sc_hd__dfxtp_1 _29848_ (.CLK(_00399_),
    .D(_01583_),
    .Q(\rvcpu.dp.rf.reg_file_arr[18][11] ));
 sky130_fd_sc_hd__dfxtp_1 _29849_ (.CLK(_00400_),
    .D(_01584_),
    .Q(\rvcpu.dp.rf.reg_file_arr[18][12] ));
 sky130_fd_sc_hd__dfxtp_1 _29850_ (.CLK(_00401_),
    .D(_01585_),
    .Q(\rvcpu.dp.rf.reg_file_arr[18][13] ));
 sky130_fd_sc_hd__dfxtp_1 _29851_ (.CLK(_00402_),
    .D(_01586_),
    .Q(\rvcpu.dp.rf.reg_file_arr[18][14] ));
 sky130_fd_sc_hd__dfxtp_1 _29852_ (.CLK(_00403_),
    .D(_01587_),
    .Q(\rvcpu.dp.rf.reg_file_arr[18][15] ));
 sky130_fd_sc_hd__dfxtp_1 _29853_ (.CLK(_00404_),
    .D(_01588_),
    .Q(\rvcpu.dp.rf.reg_file_arr[18][16] ));
 sky130_fd_sc_hd__dfxtp_1 _29854_ (.CLK(_00405_),
    .D(_01589_),
    .Q(\rvcpu.dp.rf.reg_file_arr[18][17] ));
 sky130_fd_sc_hd__dfxtp_1 _29855_ (.CLK(_00406_),
    .D(_01590_),
    .Q(\rvcpu.dp.rf.reg_file_arr[18][18] ));
 sky130_fd_sc_hd__dfxtp_1 _29856_ (.CLK(_00407_),
    .D(_01591_),
    .Q(\rvcpu.dp.rf.reg_file_arr[18][19] ));
 sky130_fd_sc_hd__dfxtp_1 _29857_ (.CLK(_00408_),
    .D(_01592_),
    .Q(\rvcpu.dp.rf.reg_file_arr[18][20] ));
 sky130_fd_sc_hd__dfxtp_1 _29858_ (.CLK(_00409_),
    .D(_01593_),
    .Q(\rvcpu.dp.rf.reg_file_arr[18][21] ));
 sky130_fd_sc_hd__dfxtp_1 _29859_ (.CLK(_00410_),
    .D(_01594_),
    .Q(\rvcpu.dp.rf.reg_file_arr[18][22] ));
 sky130_fd_sc_hd__dfxtp_1 _29860_ (.CLK(_00411_),
    .D(_01595_),
    .Q(\rvcpu.dp.rf.reg_file_arr[18][23] ));
 sky130_fd_sc_hd__dfxtp_1 _29861_ (.CLK(_00412_),
    .D(_01596_),
    .Q(\rvcpu.dp.rf.reg_file_arr[18][24] ));
 sky130_fd_sc_hd__dfxtp_1 _29862_ (.CLK(_00413_),
    .D(_01597_),
    .Q(\rvcpu.dp.rf.reg_file_arr[18][25] ));
 sky130_fd_sc_hd__dfxtp_1 _29863_ (.CLK(_00414_),
    .D(_01598_),
    .Q(\rvcpu.dp.rf.reg_file_arr[18][26] ));
 sky130_fd_sc_hd__dfxtp_1 _29864_ (.CLK(_00415_),
    .D(_01599_),
    .Q(\rvcpu.dp.rf.reg_file_arr[18][27] ));
 sky130_fd_sc_hd__dfxtp_1 _29865_ (.CLK(_00416_),
    .D(_01600_),
    .Q(\rvcpu.dp.rf.reg_file_arr[18][28] ));
 sky130_fd_sc_hd__dfxtp_1 _29866_ (.CLK(_00417_),
    .D(_01601_),
    .Q(\rvcpu.dp.rf.reg_file_arr[18][29] ));
 sky130_fd_sc_hd__dfxtp_1 _29867_ (.CLK(_00418_),
    .D(_01602_),
    .Q(\rvcpu.dp.rf.reg_file_arr[18][30] ));
 sky130_fd_sc_hd__dfxtp_1 _29868_ (.CLK(_00419_),
    .D(_01603_),
    .Q(\rvcpu.dp.rf.reg_file_arr[18][31] ));
 sky130_fd_sc_hd__dfxtp_1 _29869_ (.CLK(_00420_),
    .D(_01604_),
    .Q(\rvcpu.dp.rf.reg_file_arr[17][0] ));
 sky130_fd_sc_hd__dfxtp_1 _29870_ (.CLK(_00421_),
    .D(_01605_),
    .Q(\rvcpu.dp.rf.reg_file_arr[17][1] ));
 sky130_fd_sc_hd__dfxtp_1 _29871_ (.CLK(_00422_),
    .D(_01606_),
    .Q(\rvcpu.dp.rf.reg_file_arr[17][2] ));
 sky130_fd_sc_hd__dfxtp_1 _29872_ (.CLK(_00423_),
    .D(_01607_),
    .Q(\rvcpu.dp.rf.reg_file_arr[17][3] ));
 sky130_fd_sc_hd__dfxtp_1 _29873_ (.CLK(_00424_),
    .D(_01608_),
    .Q(\rvcpu.dp.rf.reg_file_arr[17][4] ));
 sky130_fd_sc_hd__dfxtp_1 _29874_ (.CLK(_00425_),
    .D(_01609_),
    .Q(\rvcpu.dp.rf.reg_file_arr[17][5] ));
 sky130_fd_sc_hd__dfxtp_1 _29875_ (.CLK(_00426_),
    .D(_01610_),
    .Q(\rvcpu.dp.rf.reg_file_arr[17][6] ));
 sky130_fd_sc_hd__dfxtp_1 _29876_ (.CLK(_00427_),
    .D(_01611_),
    .Q(\rvcpu.dp.rf.reg_file_arr[17][7] ));
 sky130_fd_sc_hd__dfxtp_1 _29877_ (.CLK(_00428_),
    .D(_01612_),
    .Q(\rvcpu.dp.rf.reg_file_arr[17][8] ));
 sky130_fd_sc_hd__dfxtp_1 _29878_ (.CLK(_00429_),
    .D(_01613_),
    .Q(\rvcpu.dp.rf.reg_file_arr[17][9] ));
 sky130_fd_sc_hd__dfxtp_1 _29879_ (.CLK(_00430_),
    .D(_01614_),
    .Q(\rvcpu.dp.rf.reg_file_arr[17][10] ));
 sky130_fd_sc_hd__dfxtp_1 _29880_ (.CLK(_00431_),
    .D(_01615_),
    .Q(\rvcpu.dp.rf.reg_file_arr[17][11] ));
 sky130_fd_sc_hd__dfxtp_1 _29881_ (.CLK(_00432_),
    .D(_01616_),
    .Q(\rvcpu.dp.rf.reg_file_arr[17][12] ));
 sky130_fd_sc_hd__dfxtp_1 _29882_ (.CLK(_00433_),
    .D(_01617_),
    .Q(\rvcpu.dp.rf.reg_file_arr[17][13] ));
 sky130_fd_sc_hd__dfxtp_1 _29883_ (.CLK(_00434_),
    .D(_01618_),
    .Q(\rvcpu.dp.rf.reg_file_arr[17][14] ));
 sky130_fd_sc_hd__dfxtp_1 _29884_ (.CLK(_00435_),
    .D(_01619_),
    .Q(\rvcpu.dp.rf.reg_file_arr[17][15] ));
 sky130_fd_sc_hd__dfxtp_1 _29885_ (.CLK(_00436_),
    .D(_01620_),
    .Q(\rvcpu.dp.rf.reg_file_arr[17][16] ));
 sky130_fd_sc_hd__dfxtp_1 _29886_ (.CLK(_00437_),
    .D(_01621_),
    .Q(\rvcpu.dp.rf.reg_file_arr[17][17] ));
 sky130_fd_sc_hd__dfxtp_1 _29887_ (.CLK(_00438_),
    .D(_01622_),
    .Q(\rvcpu.dp.rf.reg_file_arr[17][18] ));
 sky130_fd_sc_hd__dfxtp_1 _29888_ (.CLK(_00439_),
    .D(_01623_),
    .Q(\rvcpu.dp.rf.reg_file_arr[17][19] ));
 sky130_fd_sc_hd__dfxtp_1 _29889_ (.CLK(_00440_),
    .D(_01624_),
    .Q(\rvcpu.dp.rf.reg_file_arr[17][20] ));
 sky130_fd_sc_hd__dfxtp_1 _29890_ (.CLK(_00441_),
    .D(_01625_),
    .Q(\rvcpu.dp.rf.reg_file_arr[17][21] ));
 sky130_fd_sc_hd__dfxtp_1 _29891_ (.CLK(_00442_),
    .D(_01626_),
    .Q(\rvcpu.dp.rf.reg_file_arr[17][22] ));
 sky130_fd_sc_hd__dfxtp_1 _29892_ (.CLK(_00443_),
    .D(_01627_),
    .Q(\rvcpu.dp.rf.reg_file_arr[17][23] ));
 sky130_fd_sc_hd__dfxtp_1 _29893_ (.CLK(_00444_),
    .D(_01628_),
    .Q(\rvcpu.dp.rf.reg_file_arr[17][24] ));
 sky130_fd_sc_hd__dfxtp_1 _29894_ (.CLK(_00445_),
    .D(_01629_),
    .Q(\rvcpu.dp.rf.reg_file_arr[17][25] ));
 sky130_fd_sc_hd__dfxtp_1 _29895_ (.CLK(_00446_),
    .D(_01630_),
    .Q(\rvcpu.dp.rf.reg_file_arr[17][26] ));
 sky130_fd_sc_hd__dfxtp_1 _29896_ (.CLK(_00447_),
    .D(_01631_),
    .Q(\rvcpu.dp.rf.reg_file_arr[17][27] ));
 sky130_fd_sc_hd__dfxtp_1 _29897_ (.CLK(_00448_),
    .D(_01632_),
    .Q(\rvcpu.dp.rf.reg_file_arr[17][28] ));
 sky130_fd_sc_hd__dfxtp_1 _29898_ (.CLK(_00449_),
    .D(_01633_),
    .Q(\rvcpu.dp.rf.reg_file_arr[17][29] ));
 sky130_fd_sc_hd__dfxtp_1 _29899_ (.CLK(_00450_),
    .D(_01634_),
    .Q(\rvcpu.dp.rf.reg_file_arr[17][30] ));
 sky130_fd_sc_hd__dfxtp_1 _29900_ (.CLK(_00451_),
    .D(_01635_),
    .Q(\rvcpu.dp.rf.reg_file_arr[17][31] ));
 sky130_fd_sc_hd__dfxtp_1 _29901_ (.CLK(clk),
    .D(_01636_),
    .Q(\datamem.data_ram[59][16] ));
 sky130_fd_sc_hd__dfxtp_1 _29902_ (.CLK(clk),
    .D(_01637_),
    .Q(\datamem.data_ram[59][17] ));
 sky130_fd_sc_hd__dfxtp_1 _29903_ (.CLK(clk),
    .D(_01638_),
    .Q(\datamem.data_ram[59][18] ));
 sky130_fd_sc_hd__dfxtp_1 _29904_ (.CLK(clk),
    .D(_01639_),
    .Q(\datamem.data_ram[59][19] ));
 sky130_fd_sc_hd__dfxtp_1 _29905_ (.CLK(clk),
    .D(_01640_),
    .Q(\datamem.data_ram[59][20] ));
 sky130_fd_sc_hd__dfxtp_1 _29906_ (.CLK(clk),
    .D(_01641_),
    .Q(\datamem.data_ram[59][21] ));
 sky130_fd_sc_hd__dfxtp_1 _29907_ (.CLK(clk),
    .D(_01642_),
    .Q(\datamem.data_ram[59][22] ));
 sky130_fd_sc_hd__dfxtp_1 _29908_ (.CLK(clk),
    .D(_01643_),
    .Q(\datamem.data_ram[59][23] ));
 sky130_fd_sc_hd__dfxtp_1 _29909_ (.CLK(_00452_),
    .D(_01644_),
    .Q(\rvcpu.dp.rf.reg_file_arr[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 _29910_ (.CLK(_00453_),
    .D(_01645_),
    .Q(\rvcpu.dp.rf.reg_file_arr[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 _29911_ (.CLK(_00454_),
    .D(_01646_),
    .Q(\rvcpu.dp.rf.reg_file_arr[16][2] ));
 sky130_fd_sc_hd__dfxtp_1 _29912_ (.CLK(_00455_),
    .D(_01647_),
    .Q(\rvcpu.dp.rf.reg_file_arr[16][3] ));
 sky130_fd_sc_hd__dfxtp_1 _29913_ (.CLK(_00456_),
    .D(_01648_),
    .Q(\rvcpu.dp.rf.reg_file_arr[16][4] ));
 sky130_fd_sc_hd__dfxtp_1 _29914_ (.CLK(_00457_),
    .D(_01649_),
    .Q(\rvcpu.dp.rf.reg_file_arr[16][5] ));
 sky130_fd_sc_hd__dfxtp_1 _29915_ (.CLK(_00458_),
    .D(_01650_),
    .Q(\rvcpu.dp.rf.reg_file_arr[16][6] ));
 sky130_fd_sc_hd__dfxtp_1 _29916_ (.CLK(_00459_),
    .D(_01651_),
    .Q(\rvcpu.dp.rf.reg_file_arr[16][7] ));
 sky130_fd_sc_hd__dfxtp_1 _29917_ (.CLK(_00460_),
    .D(_01652_),
    .Q(\rvcpu.dp.rf.reg_file_arr[16][8] ));
 sky130_fd_sc_hd__dfxtp_1 _29918_ (.CLK(_00461_),
    .D(_01653_),
    .Q(\rvcpu.dp.rf.reg_file_arr[16][9] ));
 sky130_fd_sc_hd__dfxtp_1 _29919_ (.CLK(_00462_),
    .D(_01654_),
    .Q(\rvcpu.dp.rf.reg_file_arr[16][10] ));
 sky130_fd_sc_hd__dfxtp_1 _29920_ (.CLK(_00463_),
    .D(_01655_),
    .Q(\rvcpu.dp.rf.reg_file_arr[16][11] ));
 sky130_fd_sc_hd__dfxtp_1 _29921_ (.CLK(_00464_),
    .D(_01656_),
    .Q(\rvcpu.dp.rf.reg_file_arr[16][12] ));
 sky130_fd_sc_hd__dfxtp_1 _29922_ (.CLK(_00465_),
    .D(_01657_),
    .Q(\rvcpu.dp.rf.reg_file_arr[16][13] ));
 sky130_fd_sc_hd__dfxtp_1 _29923_ (.CLK(_00466_),
    .D(_01658_),
    .Q(\rvcpu.dp.rf.reg_file_arr[16][14] ));
 sky130_fd_sc_hd__dfxtp_1 _29924_ (.CLK(_00467_),
    .D(_01659_),
    .Q(\rvcpu.dp.rf.reg_file_arr[16][15] ));
 sky130_fd_sc_hd__dfxtp_1 _29925_ (.CLK(_00468_),
    .D(_01660_),
    .Q(\rvcpu.dp.rf.reg_file_arr[16][16] ));
 sky130_fd_sc_hd__dfxtp_1 _29926_ (.CLK(_00469_),
    .D(_01661_),
    .Q(\rvcpu.dp.rf.reg_file_arr[16][17] ));
 sky130_fd_sc_hd__dfxtp_1 _29927_ (.CLK(_00470_),
    .D(_01662_),
    .Q(\rvcpu.dp.rf.reg_file_arr[16][18] ));
 sky130_fd_sc_hd__dfxtp_1 _29928_ (.CLK(_00471_),
    .D(_01663_),
    .Q(\rvcpu.dp.rf.reg_file_arr[16][19] ));
 sky130_fd_sc_hd__dfxtp_1 _29929_ (.CLK(_00472_),
    .D(_01664_),
    .Q(\rvcpu.dp.rf.reg_file_arr[16][20] ));
 sky130_fd_sc_hd__dfxtp_1 _29930_ (.CLK(_00473_),
    .D(_01665_),
    .Q(\rvcpu.dp.rf.reg_file_arr[16][21] ));
 sky130_fd_sc_hd__dfxtp_1 _29931_ (.CLK(_00474_),
    .D(_01666_),
    .Q(\rvcpu.dp.rf.reg_file_arr[16][22] ));
 sky130_fd_sc_hd__dfxtp_1 _29932_ (.CLK(_00475_),
    .D(_01667_),
    .Q(\rvcpu.dp.rf.reg_file_arr[16][23] ));
 sky130_fd_sc_hd__dfxtp_1 _29933_ (.CLK(_00476_),
    .D(_01668_),
    .Q(\rvcpu.dp.rf.reg_file_arr[16][24] ));
 sky130_fd_sc_hd__dfxtp_1 _29934_ (.CLK(_00477_),
    .D(_01669_),
    .Q(\rvcpu.dp.rf.reg_file_arr[16][25] ));
 sky130_fd_sc_hd__dfxtp_1 _29935_ (.CLK(_00478_),
    .D(_01670_),
    .Q(\rvcpu.dp.rf.reg_file_arr[16][26] ));
 sky130_fd_sc_hd__dfxtp_1 _29936_ (.CLK(_00479_),
    .D(_01671_),
    .Q(\rvcpu.dp.rf.reg_file_arr[16][27] ));
 sky130_fd_sc_hd__dfxtp_1 _29937_ (.CLK(_00480_),
    .D(_01672_),
    .Q(\rvcpu.dp.rf.reg_file_arr[16][28] ));
 sky130_fd_sc_hd__dfxtp_1 _29938_ (.CLK(_00481_),
    .D(_01673_),
    .Q(\rvcpu.dp.rf.reg_file_arr[16][29] ));
 sky130_fd_sc_hd__dfxtp_1 _29939_ (.CLK(_00482_),
    .D(_01674_),
    .Q(\rvcpu.dp.rf.reg_file_arr[16][30] ));
 sky130_fd_sc_hd__dfxtp_1 _29940_ (.CLK(_00483_),
    .D(_01675_),
    .Q(\rvcpu.dp.rf.reg_file_arr[16][31] ));
 sky130_fd_sc_hd__dfxtp_1 _29941_ (.CLK(_00484_),
    .D(_01676_),
    .Q(\rvcpu.dp.rf.reg_file_arr[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _29942_ (.CLK(_00485_),
    .D(_01677_),
    .Q(\rvcpu.dp.rf.reg_file_arr[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _29943_ (.CLK(_00486_),
    .D(_01678_),
    .Q(\rvcpu.dp.rf.reg_file_arr[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _29944_ (.CLK(_00487_),
    .D(_01679_),
    .Q(\rvcpu.dp.rf.reg_file_arr[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _29945_ (.CLK(_00488_),
    .D(_01680_),
    .Q(\rvcpu.dp.rf.reg_file_arr[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _29946_ (.CLK(_00489_),
    .D(_01681_),
    .Q(\rvcpu.dp.rf.reg_file_arr[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _29947_ (.CLK(_00490_),
    .D(_01682_),
    .Q(\rvcpu.dp.rf.reg_file_arr[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _29948_ (.CLK(_00491_),
    .D(_01683_),
    .Q(\rvcpu.dp.rf.reg_file_arr[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _29949_ (.CLK(_00492_),
    .D(_01684_),
    .Q(\rvcpu.dp.rf.reg_file_arr[15][8] ));
 sky130_fd_sc_hd__dfxtp_1 _29950_ (.CLK(_00493_),
    .D(_01685_),
    .Q(\rvcpu.dp.rf.reg_file_arr[15][9] ));
 sky130_fd_sc_hd__dfxtp_1 _29951_ (.CLK(_00494_),
    .D(_01686_),
    .Q(\rvcpu.dp.rf.reg_file_arr[15][10] ));
 sky130_fd_sc_hd__dfxtp_1 _29952_ (.CLK(_00495_),
    .D(_01687_),
    .Q(\rvcpu.dp.rf.reg_file_arr[15][11] ));
 sky130_fd_sc_hd__dfxtp_1 _29953_ (.CLK(_00496_),
    .D(_01688_),
    .Q(\rvcpu.dp.rf.reg_file_arr[15][12] ));
 sky130_fd_sc_hd__dfxtp_1 _29954_ (.CLK(_00497_),
    .D(_01689_),
    .Q(\rvcpu.dp.rf.reg_file_arr[15][13] ));
 sky130_fd_sc_hd__dfxtp_1 _29955_ (.CLK(_00498_),
    .D(_01690_),
    .Q(\rvcpu.dp.rf.reg_file_arr[15][14] ));
 sky130_fd_sc_hd__dfxtp_1 _29956_ (.CLK(_00499_),
    .D(_01691_),
    .Q(\rvcpu.dp.rf.reg_file_arr[15][15] ));
 sky130_fd_sc_hd__dfxtp_1 _29957_ (.CLK(_00500_),
    .D(_01692_),
    .Q(\rvcpu.dp.rf.reg_file_arr[15][16] ));
 sky130_fd_sc_hd__dfxtp_1 _29958_ (.CLK(_00501_),
    .D(_01693_),
    .Q(\rvcpu.dp.rf.reg_file_arr[15][17] ));
 sky130_fd_sc_hd__dfxtp_1 _29959_ (.CLK(_00502_),
    .D(_01694_),
    .Q(\rvcpu.dp.rf.reg_file_arr[15][18] ));
 sky130_fd_sc_hd__dfxtp_1 _29960_ (.CLK(_00503_),
    .D(_01695_),
    .Q(\rvcpu.dp.rf.reg_file_arr[15][19] ));
 sky130_fd_sc_hd__dfxtp_1 _29961_ (.CLK(_00504_),
    .D(_01696_),
    .Q(\rvcpu.dp.rf.reg_file_arr[15][20] ));
 sky130_fd_sc_hd__dfxtp_1 _29962_ (.CLK(_00505_),
    .D(_01697_),
    .Q(\rvcpu.dp.rf.reg_file_arr[15][21] ));
 sky130_fd_sc_hd__dfxtp_1 _29963_ (.CLK(_00506_),
    .D(_01698_),
    .Q(\rvcpu.dp.rf.reg_file_arr[15][22] ));
 sky130_fd_sc_hd__dfxtp_1 _29964_ (.CLK(_00507_),
    .D(_01699_),
    .Q(\rvcpu.dp.rf.reg_file_arr[15][23] ));
 sky130_fd_sc_hd__dfxtp_1 _29965_ (.CLK(_00508_),
    .D(_01700_),
    .Q(\rvcpu.dp.rf.reg_file_arr[15][24] ));
 sky130_fd_sc_hd__dfxtp_1 _29966_ (.CLK(_00509_),
    .D(_01701_),
    .Q(\rvcpu.dp.rf.reg_file_arr[15][25] ));
 sky130_fd_sc_hd__dfxtp_1 _29967_ (.CLK(_00510_),
    .D(_01702_),
    .Q(\rvcpu.dp.rf.reg_file_arr[15][26] ));
 sky130_fd_sc_hd__dfxtp_1 _29968_ (.CLK(_00511_),
    .D(_01703_),
    .Q(\rvcpu.dp.rf.reg_file_arr[15][27] ));
 sky130_fd_sc_hd__dfxtp_1 _29969_ (.CLK(_00512_),
    .D(_01704_),
    .Q(\rvcpu.dp.rf.reg_file_arr[15][28] ));
 sky130_fd_sc_hd__dfxtp_1 _29970_ (.CLK(_00513_),
    .D(_01705_),
    .Q(\rvcpu.dp.rf.reg_file_arr[15][29] ));
 sky130_fd_sc_hd__dfxtp_1 _29971_ (.CLK(_00514_),
    .D(_01706_),
    .Q(\rvcpu.dp.rf.reg_file_arr[15][30] ));
 sky130_fd_sc_hd__dfxtp_1 _29972_ (.CLK(_00515_),
    .D(_01707_),
    .Q(\rvcpu.dp.rf.reg_file_arr[15][31] ));
 sky130_fd_sc_hd__dfxtp_1 _29973_ (.CLK(_00516_),
    .D(_01708_),
    .Q(\rvcpu.dp.rf.reg_file_arr[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _29974_ (.CLK(_00517_),
    .D(_01709_),
    .Q(\rvcpu.dp.rf.reg_file_arr[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _29975_ (.CLK(_00518_),
    .D(_01710_),
    .Q(\rvcpu.dp.rf.reg_file_arr[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _29976_ (.CLK(_00519_),
    .D(_01711_),
    .Q(\rvcpu.dp.rf.reg_file_arr[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _29977_ (.CLK(_00520_),
    .D(_01712_),
    .Q(\rvcpu.dp.rf.reg_file_arr[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _29978_ (.CLK(_00521_),
    .D(_01713_),
    .Q(\rvcpu.dp.rf.reg_file_arr[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _29979_ (.CLK(_00522_),
    .D(_01714_),
    .Q(\rvcpu.dp.rf.reg_file_arr[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _29980_ (.CLK(_00523_),
    .D(_01715_),
    .Q(\rvcpu.dp.rf.reg_file_arr[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _29981_ (.CLK(_00524_),
    .D(_01716_),
    .Q(\rvcpu.dp.rf.reg_file_arr[14][8] ));
 sky130_fd_sc_hd__dfxtp_1 _29982_ (.CLK(_00525_),
    .D(_01717_),
    .Q(\rvcpu.dp.rf.reg_file_arr[14][9] ));
 sky130_fd_sc_hd__dfxtp_1 _29983_ (.CLK(_00526_),
    .D(_01718_),
    .Q(\rvcpu.dp.rf.reg_file_arr[14][10] ));
 sky130_fd_sc_hd__dfxtp_1 _29984_ (.CLK(_00527_),
    .D(_01719_),
    .Q(\rvcpu.dp.rf.reg_file_arr[14][11] ));
 sky130_fd_sc_hd__dfxtp_1 _29985_ (.CLK(_00528_),
    .D(_01720_),
    .Q(\rvcpu.dp.rf.reg_file_arr[14][12] ));
 sky130_fd_sc_hd__dfxtp_1 _29986_ (.CLK(_00529_),
    .D(_01721_),
    .Q(\rvcpu.dp.rf.reg_file_arr[14][13] ));
 sky130_fd_sc_hd__dfxtp_1 _29987_ (.CLK(_00530_),
    .D(_01722_),
    .Q(\rvcpu.dp.rf.reg_file_arr[14][14] ));
 sky130_fd_sc_hd__dfxtp_1 _29988_ (.CLK(_00531_),
    .D(_01723_),
    .Q(\rvcpu.dp.rf.reg_file_arr[14][15] ));
 sky130_fd_sc_hd__dfxtp_1 _29989_ (.CLK(_00532_),
    .D(_01724_),
    .Q(\rvcpu.dp.rf.reg_file_arr[14][16] ));
 sky130_fd_sc_hd__dfxtp_1 _29990_ (.CLK(_00533_),
    .D(_01725_),
    .Q(\rvcpu.dp.rf.reg_file_arr[14][17] ));
 sky130_fd_sc_hd__dfxtp_1 _29991_ (.CLK(_00534_),
    .D(_01726_),
    .Q(\rvcpu.dp.rf.reg_file_arr[14][18] ));
 sky130_fd_sc_hd__dfxtp_1 _29992_ (.CLK(_00535_),
    .D(_01727_),
    .Q(\rvcpu.dp.rf.reg_file_arr[14][19] ));
 sky130_fd_sc_hd__dfxtp_1 _29993_ (.CLK(_00536_),
    .D(_01728_),
    .Q(\rvcpu.dp.rf.reg_file_arr[14][20] ));
 sky130_fd_sc_hd__dfxtp_1 _29994_ (.CLK(_00537_),
    .D(_01729_),
    .Q(\rvcpu.dp.rf.reg_file_arr[14][21] ));
 sky130_fd_sc_hd__dfxtp_1 _29995_ (.CLK(_00538_),
    .D(_01730_),
    .Q(\rvcpu.dp.rf.reg_file_arr[14][22] ));
 sky130_fd_sc_hd__dfxtp_1 _29996_ (.CLK(_00539_),
    .D(_01731_),
    .Q(\rvcpu.dp.rf.reg_file_arr[14][23] ));
 sky130_fd_sc_hd__dfxtp_1 _29997_ (.CLK(_00540_),
    .D(_01732_),
    .Q(\rvcpu.dp.rf.reg_file_arr[14][24] ));
 sky130_fd_sc_hd__dfxtp_1 _29998_ (.CLK(_00541_),
    .D(_01733_),
    .Q(\rvcpu.dp.rf.reg_file_arr[14][25] ));
 sky130_fd_sc_hd__dfxtp_1 _29999_ (.CLK(_00542_),
    .D(_01734_),
    .Q(\rvcpu.dp.rf.reg_file_arr[14][26] ));
 sky130_fd_sc_hd__dfxtp_1 _30000_ (.CLK(_00543_),
    .D(_01735_),
    .Q(\rvcpu.dp.rf.reg_file_arr[14][27] ));
 sky130_fd_sc_hd__dfxtp_1 _30001_ (.CLK(_00544_),
    .D(_01736_),
    .Q(\rvcpu.dp.rf.reg_file_arr[14][28] ));
 sky130_fd_sc_hd__dfxtp_1 _30002_ (.CLK(_00545_),
    .D(_01737_),
    .Q(\rvcpu.dp.rf.reg_file_arr[14][29] ));
 sky130_fd_sc_hd__dfxtp_1 _30003_ (.CLK(_00546_),
    .D(_01738_),
    .Q(\rvcpu.dp.rf.reg_file_arr[14][30] ));
 sky130_fd_sc_hd__dfxtp_1 _30004_ (.CLK(_00547_),
    .D(_01739_),
    .Q(\rvcpu.dp.rf.reg_file_arr[14][31] ));
 sky130_fd_sc_hd__dfxtp_1 _30005_ (.CLK(clk),
    .D(_01740_),
    .Q(\datamem.data_ram[59][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30006_ (.CLK(clk),
    .D(_01741_),
    .Q(\datamem.data_ram[59][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30007_ (.CLK(clk),
    .D(_01742_),
    .Q(\datamem.data_ram[59][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30008_ (.CLK(clk),
    .D(_01743_),
    .Q(\datamem.data_ram[59][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30009_ (.CLK(clk),
    .D(_01744_),
    .Q(\datamem.data_ram[59][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30010_ (.CLK(clk),
    .D(_01745_),
    .Q(\datamem.data_ram[59][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30011_ (.CLK(clk),
    .D(_01746_),
    .Q(\datamem.data_ram[59][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30012_ (.CLK(clk),
    .D(_01747_),
    .Q(\datamem.data_ram[59][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30013_ (.CLK(_00548_),
    .D(_01748_),
    .Q(\rvcpu.dp.rf.reg_file_arr[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _30014_ (.CLK(_00549_),
    .D(_01749_),
    .Q(\rvcpu.dp.rf.reg_file_arr[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _30015_ (.CLK(_00550_),
    .D(_01750_),
    .Q(\rvcpu.dp.rf.reg_file_arr[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _30016_ (.CLK(_00551_),
    .D(_01751_),
    .Q(\rvcpu.dp.rf.reg_file_arr[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _30017_ (.CLK(_00552_),
    .D(_01752_),
    .Q(\rvcpu.dp.rf.reg_file_arr[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _30018_ (.CLK(_00553_),
    .D(_01753_),
    .Q(\rvcpu.dp.rf.reg_file_arr[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _30019_ (.CLK(_00554_),
    .D(_01754_),
    .Q(\rvcpu.dp.rf.reg_file_arr[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _30020_ (.CLK(_00555_),
    .D(_01755_),
    .Q(\rvcpu.dp.rf.reg_file_arr[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _30021_ (.CLK(_00556_),
    .D(_01756_),
    .Q(\rvcpu.dp.rf.reg_file_arr[13][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30022_ (.CLK(_00557_),
    .D(_01757_),
    .Q(\rvcpu.dp.rf.reg_file_arr[13][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30023_ (.CLK(_00558_),
    .D(_01758_),
    .Q(\rvcpu.dp.rf.reg_file_arr[13][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30024_ (.CLK(_00559_),
    .D(_01759_),
    .Q(\rvcpu.dp.rf.reg_file_arr[13][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30025_ (.CLK(_00560_),
    .D(_01760_),
    .Q(\rvcpu.dp.rf.reg_file_arr[13][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30026_ (.CLK(_00561_),
    .D(_01761_),
    .Q(\rvcpu.dp.rf.reg_file_arr[13][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30027_ (.CLK(_00562_),
    .D(_01762_),
    .Q(\rvcpu.dp.rf.reg_file_arr[13][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30028_ (.CLK(_00563_),
    .D(_01763_),
    .Q(\rvcpu.dp.rf.reg_file_arr[13][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30029_ (.CLK(_00564_),
    .D(_01764_),
    .Q(\rvcpu.dp.rf.reg_file_arr[13][16] ));
 sky130_fd_sc_hd__dfxtp_1 _30030_ (.CLK(_00565_),
    .D(_01765_),
    .Q(\rvcpu.dp.rf.reg_file_arr[13][17] ));
 sky130_fd_sc_hd__dfxtp_1 _30031_ (.CLK(_00566_),
    .D(_01766_),
    .Q(\rvcpu.dp.rf.reg_file_arr[13][18] ));
 sky130_fd_sc_hd__dfxtp_1 _30032_ (.CLK(_00567_),
    .D(_01767_),
    .Q(\rvcpu.dp.rf.reg_file_arr[13][19] ));
 sky130_fd_sc_hd__dfxtp_1 _30033_ (.CLK(_00568_),
    .D(_01768_),
    .Q(\rvcpu.dp.rf.reg_file_arr[13][20] ));
 sky130_fd_sc_hd__dfxtp_1 _30034_ (.CLK(_00569_),
    .D(_01769_),
    .Q(\rvcpu.dp.rf.reg_file_arr[13][21] ));
 sky130_fd_sc_hd__dfxtp_1 _30035_ (.CLK(_00570_),
    .D(_01770_),
    .Q(\rvcpu.dp.rf.reg_file_arr[13][22] ));
 sky130_fd_sc_hd__dfxtp_1 _30036_ (.CLK(_00571_),
    .D(_01771_),
    .Q(\rvcpu.dp.rf.reg_file_arr[13][23] ));
 sky130_fd_sc_hd__dfxtp_1 _30037_ (.CLK(_00572_),
    .D(_01772_),
    .Q(\rvcpu.dp.rf.reg_file_arr[13][24] ));
 sky130_fd_sc_hd__dfxtp_1 _30038_ (.CLK(_00573_),
    .D(_01773_),
    .Q(\rvcpu.dp.rf.reg_file_arr[13][25] ));
 sky130_fd_sc_hd__dfxtp_1 _30039_ (.CLK(_00574_),
    .D(_01774_),
    .Q(\rvcpu.dp.rf.reg_file_arr[13][26] ));
 sky130_fd_sc_hd__dfxtp_1 _30040_ (.CLK(_00575_),
    .D(_01775_),
    .Q(\rvcpu.dp.rf.reg_file_arr[13][27] ));
 sky130_fd_sc_hd__dfxtp_1 _30041_ (.CLK(_00576_),
    .D(_01776_),
    .Q(\rvcpu.dp.rf.reg_file_arr[13][28] ));
 sky130_fd_sc_hd__dfxtp_1 _30042_ (.CLK(_00577_),
    .D(_01777_),
    .Q(\rvcpu.dp.rf.reg_file_arr[13][29] ));
 sky130_fd_sc_hd__dfxtp_1 _30043_ (.CLK(_00578_),
    .D(_01778_),
    .Q(\rvcpu.dp.rf.reg_file_arr[13][30] ));
 sky130_fd_sc_hd__dfxtp_1 _30044_ (.CLK(_00579_),
    .D(_01779_),
    .Q(\rvcpu.dp.rf.reg_file_arr[13][31] ));
 sky130_fd_sc_hd__dfxtp_1 _30045_ (.CLK(_00580_),
    .D(_01780_),
    .Q(\rvcpu.dp.rf.reg_file_arr[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _30046_ (.CLK(_00581_),
    .D(_01781_),
    .Q(\rvcpu.dp.rf.reg_file_arr[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _30047_ (.CLK(_00582_),
    .D(_01782_),
    .Q(\rvcpu.dp.rf.reg_file_arr[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _30048_ (.CLK(_00583_),
    .D(_01783_),
    .Q(\rvcpu.dp.rf.reg_file_arr[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _30049_ (.CLK(_00584_),
    .D(_01784_),
    .Q(\rvcpu.dp.rf.reg_file_arr[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _30050_ (.CLK(_00585_),
    .D(_01785_),
    .Q(\rvcpu.dp.rf.reg_file_arr[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _30051_ (.CLK(_00586_),
    .D(_01786_),
    .Q(\rvcpu.dp.rf.reg_file_arr[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _30052_ (.CLK(_00587_),
    .D(_01787_),
    .Q(\rvcpu.dp.rf.reg_file_arr[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _30053_ (.CLK(_00588_),
    .D(_01788_),
    .Q(\rvcpu.dp.rf.reg_file_arr[12][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30054_ (.CLK(_00589_),
    .D(_01789_),
    .Q(\rvcpu.dp.rf.reg_file_arr[12][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30055_ (.CLK(_00590_),
    .D(_01790_),
    .Q(\rvcpu.dp.rf.reg_file_arr[12][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30056_ (.CLK(_00591_),
    .D(_01791_),
    .Q(\rvcpu.dp.rf.reg_file_arr[12][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30057_ (.CLK(_00592_),
    .D(_01792_),
    .Q(\rvcpu.dp.rf.reg_file_arr[12][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30058_ (.CLK(_00593_),
    .D(_01793_),
    .Q(\rvcpu.dp.rf.reg_file_arr[12][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30059_ (.CLK(_00594_),
    .D(_01794_),
    .Q(\rvcpu.dp.rf.reg_file_arr[12][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30060_ (.CLK(_00595_),
    .D(_01795_),
    .Q(\rvcpu.dp.rf.reg_file_arr[12][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30061_ (.CLK(_00596_),
    .D(_01796_),
    .Q(\rvcpu.dp.rf.reg_file_arr[12][16] ));
 sky130_fd_sc_hd__dfxtp_1 _30062_ (.CLK(_00597_),
    .D(_01797_),
    .Q(\rvcpu.dp.rf.reg_file_arr[12][17] ));
 sky130_fd_sc_hd__dfxtp_1 _30063_ (.CLK(_00598_),
    .D(_01798_),
    .Q(\rvcpu.dp.rf.reg_file_arr[12][18] ));
 sky130_fd_sc_hd__dfxtp_1 _30064_ (.CLK(_00599_),
    .D(_01799_),
    .Q(\rvcpu.dp.rf.reg_file_arr[12][19] ));
 sky130_fd_sc_hd__dfxtp_1 _30065_ (.CLK(_00600_),
    .D(_01800_),
    .Q(\rvcpu.dp.rf.reg_file_arr[12][20] ));
 sky130_fd_sc_hd__dfxtp_1 _30066_ (.CLK(_00601_),
    .D(_01801_),
    .Q(\rvcpu.dp.rf.reg_file_arr[12][21] ));
 sky130_fd_sc_hd__dfxtp_1 _30067_ (.CLK(_00602_),
    .D(_01802_),
    .Q(\rvcpu.dp.rf.reg_file_arr[12][22] ));
 sky130_fd_sc_hd__dfxtp_1 _30068_ (.CLK(_00603_),
    .D(_01803_),
    .Q(\rvcpu.dp.rf.reg_file_arr[12][23] ));
 sky130_fd_sc_hd__dfxtp_1 _30069_ (.CLK(_00604_),
    .D(_01804_),
    .Q(\rvcpu.dp.rf.reg_file_arr[12][24] ));
 sky130_fd_sc_hd__dfxtp_1 _30070_ (.CLK(_00605_),
    .D(_01805_),
    .Q(\rvcpu.dp.rf.reg_file_arr[12][25] ));
 sky130_fd_sc_hd__dfxtp_1 _30071_ (.CLK(_00606_),
    .D(_01806_),
    .Q(\rvcpu.dp.rf.reg_file_arr[12][26] ));
 sky130_fd_sc_hd__dfxtp_1 _30072_ (.CLK(_00607_),
    .D(_01807_),
    .Q(\rvcpu.dp.rf.reg_file_arr[12][27] ));
 sky130_fd_sc_hd__dfxtp_1 _30073_ (.CLK(_00608_),
    .D(_01808_),
    .Q(\rvcpu.dp.rf.reg_file_arr[12][28] ));
 sky130_fd_sc_hd__dfxtp_1 _30074_ (.CLK(_00609_),
    .D(_01809_),
    .Q(\rvcpu.dp.rf.reg_file_arr[12][29] ));
 sky130_fd_sc_hd__dfxtp_1 _30075_ (.CLK(_00610_),
    .D(_01810_),
    .Q(\rvcpu.dp.rf.reg_file_arr[12][30] ));
 sky130_fd_sc_hd__dfxtp_1 _30076_ (.CLK(_00611_),
    .D(_01811_),
    .Q(\rvcpu.dp.rf.reg_file_arr[12][31] ));
 sky130_fd_sc_hd__dfxtp_1 _30077_ (.CLK(_00612_),
    .D(_01812_),
    .Q(\rvcpu.dp.rf.reg_file_arr[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _30078_ (.CLK(_00613_),
    .D(_01813_),
    .Q(\rvcpu.dp.rf.reg_file_arr[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _30079_ (.CLK(_00614_),
    .D(_01814_),
    .Q(\rvcpu.dp.rf.reg_file_arr[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _30080_ (.CLK(_00615_),
    .D(_01815_),
    .Q(\rvcpu.dp.rf.reg_file_arr[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _30081_ (.CLK(_00616_),
    .D(_01816_),
    .Q(\rvcpu.dp.rf.reg_file_arr[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _30082_ (.CLK(_00617_),
    .D(_01817_),
    .Q(\rvcpu.dp.rf.reg_file_arr[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _30083_ (.CLK(_00618_),
    .D(_01818_),
    .Q(\rvcpu.dp.rf.reg_file_arr[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _30084_ (.CLK(_00619_),
    .D(_01819_),
    .Q(\rvcpu.dp.rf.reg_file_arr[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _30085_ (.CLK(_00620_),
    .D(_01820_),
    .Q(\rvcpu.dp.rf.reg_file_arr[11][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30086_ (.CLK(_00621_),
    .D(_01821_),
    .Q(\rvcpu.dp.rf.reg_file_arr[11][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30087_ (.CLK(_00622_),
    .D(_01822_),
    .Q(\rvcpu.dp.rf.reg_file_arr[11][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30088_ (.CLK(_00623_),
    .D(_01823_),
    .Q(\rvcpu.dp.rf.reg_file_arr[11][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30089_ (.CLK(_00624_),
    .D(_01824_),
    .Q(\rvcpu.dp.rf.reg_file_arr[11][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30090_ (.CLK(_00625_),
    .D(_01825_),
    .Q(\rvcpu.dp.rf.reg_file_arr[11][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30091_ (.CLK(_00626_),
    .D(_01826_),
    .Q(\rvcpu.dp.rf.reg_file_arr[11][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30092_ (.CLK(_00627_),
    .D(_01827_),
    .Q(\rvcpu.dp.rf.reg_file_arr[11][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30093_ (.CLK(_00628_),
    .D(_01828_),
    .Q(\rvcpu.dp.rf.reg_file_arr[11][16] ));
 sky130_fd_sc_hd__dfxtp_1 _30094_ (.CLK(_00629_),
    .D(_01829_),
    .Q(\rvcpu.dp.rf.reg_file_arr[11][17] ));
 sky130_fd_sc_hd__dfxtp_1 _30095_ (.CLK(_00630_),
    .D(_01830_),
    .Q(\rvcpu.dp.rf.reg_file_arr[11][18] ));
 sky130_fd_sc_hd__dfxtp_1 _30096_ (.CLK(_00631_),
    .D(_01831_),
    .Q(\rvcpu.dp.rf.reg_file_arr[11][19] ));
 sky130_fd_sc_hd__dfxtp_1 _30097_ (.CLK(_00632_),
    .D(_01832_),
    .Q(\rvcpu.dp.rf.reg_file_arr[11][20] ));
 sky130_fd_sc_hd__dfxtp_1 _30098_ (.CLK(_00633_),
    .D(_01833_),
    .Q(\rvcpu.dp.rf.reg_file_arr[11][21] ));
 sky130_fd_sc_hd__dfxtp_1 _30099_ (.CLK(_00634_),
    .D(_01834_),
    .Q(\rvcpu.dp.rf.reg_file_arr[11][22] ));
 sky130_fd_sc_hd__dfxtp_1 _30100_ (.CLK(_00635_),
    .D(_01835_),
    .Q(\rvcpu.dp.rf.reg_file_arr[11][23] ));
 sky130_fd_sc_hd__dfxtp_1 _30101_ (.CLK(_00636_),
    .D(_01836_),
    .Q(\rvcpu.dp.rf.reg_file_arr[11][24] ));
 sky130_fd_sc_hd__dfxtp_1 _30102_ (.CLK(_00637_),
    .D(_01837_),
    .Q(\rvcpu.dp.rf.reg_file_arr[11][25] ));
 sky130_fd_sc_hd__dfxtp_1 _30103_ (.CLK(_00638_),
    .D(_01838_),
    .Q(\rvcpu.dp.rf.reg_file_arr[11][26] ));
 sky130_fd_sc_hd__dfxtp_1 _30104_ (.CLK(_00639_),
    .D(_01839_),
    .Q(\rvcpu.dp.rf.reg_file_arr[11][27] ));
 sky130_fd_sc_hd__dfxtp_1 _30105_ (.CLK(_00640_),
    .D(_01840_),
    .Q(\rvcpu.dp.rf.reg_file_arr[11][28] ));
 sky130_fd_sc_hd__dfxtp_1 _30106_ (.CLK(_00641_),
    .D(_01841_),
    .Q(\rvcpu.dp.rf.reg_file_arr[11][29] ));
 sky130_fd_sc_hd__dfxtp_1 _30107_ (.CLK(_00642_),
    .D(_01842_),
    .Q(\rvcpu.dp.rf.reg_file_arr[11][30] ));
 sky130_fd_sc_hd__dfxtp_1 _30108_ (.CLK(_00643_),
    .D(_01843_),
    .Q(\rvcpu.dp.rf.reg_file_arr[11][31] ));
 sky130_fd_sc_hd__dfxtp_1 _30109_ (.CLK(_00644_),
    .D(_01844_),
    .Q(\rvcpu.dp.rf.reg_file_arr[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _30110_ (.CLK(_00645_),
    .D(_01845_),
    .Q(\rvcpu.dp.rf.reg_file_arr[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _30111_ (.CLK(_00646_),
    .D(_01846_),
    .Q(\rvcpu.dp.rf.reg_file_arr[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _30112_ (.CLK(_00647_),
    .D(_01847_),
    .Q(\rvcpu.dp.rf.reg_file_arr[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _30113_ (.CLK(_00648_),
    .D(_01848_),
    .Q(\rvcpu.dp.rf.reg_file_arr[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _30114_ (.CLK(_00649_),
    .D(_01849_),
    .Q(\rvcpu.dp.rf.reg_file_arr[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _30115_ (.CLK(_00650_),
    .D(_01850_),
    .Q(\rvcpu.dp.rf.reg_file_arr[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _30116_ (.CLK(_00651_),
    .D(_01851_),
    .Q(\rvcpu.dp.rf.reg_file_arr[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _30117_ (.CLK(_00652_),
    .D(_01852_),
    .Q(\rvcpu.dp.rf.reg_file_arr[10][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30118_ (.CLK(_00653_),
    .D(_01853_),
    .Q(\rvcpu.dp.rf.reg_file_arr[10][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30119_ (.CLK(_00654_),
    .D(_01854_),
    .Q(\rvcpu.dp.rf.reg_file_arr[10][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30120_ (.CLK(_00655_),
    .D(_01855_),
    .Q(\rvcpu.dp.rf.reg_file_arr[10][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30121_ (.CLK(_00656_),
    .D(_01856_),
    .Q(\rvcpu.dp.rf.reg_file_arr[10][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30122_ (.CLK(_00657_),
    .D(_01857_),
    .Q(\rvcpu.dp.rf.reg_file_arr[10][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30123_ (.CLK(_00658_),
    .D(_01858_),
    .Q(\rvcpu.dp.rf.reg_file_arr[10][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30124_ (.CLK(_00659_),
    .D(_01859_),
    .Q(\rvcpu.dp.rf.reg_file_arr[10][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30125_ (.CLK(_00660_),
    .D(_01860_),
    .Q(\rvcpu.dp.rf.reg_file_arr[10][16] ));
 sky130_fd_sc_hd__dfxtp_1 _30126_ (.CLK(_00661_),
    .D(_01861_),
    .Q(\rvcpu.dp.rf.reg_file_arr[10][17] ));
 sky130_fd_sc_hd__dfxtp_1 _30127_ (.CLK(_00662_),
    .D(_01862_),
    .Q(\rvcpu.dp.rf.reg_file_arr[10][18] ));
 sky130_fd_sc_hd__dfxtp_1 _30128_ (.CLK(_00663_),
    .D(_01863_),
    .Q(\rvcpu.dp.rf.reg_file_arr[10][19] ));
 sky130_fd_sc_hd__dfxtp_1 _30129_ (.CLK(_00664_),
    .D(_01864_),
    .Q(\rvcpu.dp.rf.reg_file_arr[10][20] ));
 sky130_fd_sc_hd__dfxtp_1 _30130_ (.CLK(_00665_),
    .D(_01865_),
    .Q(\rvcpu.dp.rf.reg_file_arr[10][21] ));
 sky130_fd_sc_hd__dfxtp_1 _30131_ (.CLK(_00666_),
    .D(_01866_),
    .Q(\rvcpu.dp.rf.reg_file_arr[10][22] ));
 sky130_fd_sc_hd__dfxtp_1 _30132_ (.CLK(_00667_),
    .D(_01867_),
    .Q(\rvcpu.dp.rf.reg_file_arr[10][23] ));
 sky130_fd_sc_hd__dfxtp_1 _30133_ (.CLK(_00668_),
    .D(_01868_),
    .Q(\rvcpu.dp.rf.reg_file_arr[10][24] ));
 sky130_fd_sc_hd__dfxtp_1 _30134_ (.CLK(_00669_),
    .D(_01869_),
    .Q(\rvcpu.dp.rf.reg_file_arr[10][25] ));
 sky130_fd_sc_hd__dfxtp_1 _30135_ (.CLK(_00670_),
    .D(_01870_),
    .Q(\rvcpu.dp.rf.reg_file_arr[10][26] ));
 sky130_fd_sc_hd__dfxtp_1 _30136_ (.CLK(_00671_),
    .D(_01871_),
    .Q(\rvcpu.dp.rf.reg_file_arr[10][27] ));
 sky130_fd_sc_hd__dfxtp_1 _30137_ (.CLK(_00672_),
    .D(_01872_),
    .Q(\rvcpu.dp.rf.reg_file_arr[10][28] ));
 sky130_fd_sc_hd__dfxtp_1 _30138_ (.CLK(_00673_),
    .D(_01873_),
    .Q(\rvcpu.dp.rf.reg_file_arr[10][29] ));
 sky130_fd_sc_hd__dfxtp_1 _30139_ (.CLK(_00674_),
    .D(_01874_),
    .Q(\rvcpu.dp.rf.reg_file_arr[10][30] ));
 sky130_fd_sc_hd__dfxtp_1 _30140_ (.CLK(_00675_),
    .D(_01875_),
    .Q(\rvcpu.dp.rf.reg_file_arr[10][31] ));
 sky130_fd_sc_hd__dfxtp_1 _30141_ (.CLK(_00676_),
    .D(_01876_),
    .Q(\rvcpu.dp.rf.reg_file_arr[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _30142_ (.CLK(_00677_),
    .D(_01877_),
    .Q(\rvcpu.dp.rf.reg_file_arr[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _30143_ (.CLK(_00678_),
    .D(_01878_),
    .Q(\rvcpu.dp.rf.reg_file_arr[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _30144_ (.CLK(_00679_),
    .D(_01879_),
    .Q(\rvcpu.dp.rf.reg_file_arr[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _30145_ (.CLK(_00680_),
    .D(_01880_),
    .Q(\rvcpu.dp.rf.reg_file_arr[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _30146_ (.CLK(_00681_),
    .D(_01881_),
    .Q(\rvcpu.dp.rf.reg_file_arr[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _30147_ (.CLK(_00682_),
    .D(_01882_),
    .Q(\rvcpu.dp.rf.reg_file_arr[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _30148_ (.CLK(_00683_),
    .D(_01883_),
    .Q(\rvcpu.dp.rf.reg_file_arr[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _30149_ (.CLK(_00684_),
    .D(_01884_),
    .Q(\rvcpu.dp.rf.reg_file_arr[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30150_ (.CLK(_00685_),
    .D(_01885_),
    .Q(\rvcpu.dp.rf.reg_file_arr[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30151_ (.CLK(_00686_),
    .D(_01886_),
    .Q(\rvcpu.dp.rf.reg_file_arr[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30152_ (.CLK(_00687_),
    .D(_01887_),
    .Q(\rvcpu.dp.rf.reg_file_arr[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30153_ (.CLK(_00688_),
    .D(_01888_),
    .Q(\rvcpu.dp.rf.reg_file_arr[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30154_ (.CLK(_00689_),
    .D(_01889_),
    .Q(\rvcpu.dp.rf.reg_file_arr[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30155_ (.CLK(_00690_),
    .D(_01890_),
    .Q(\rvcpu.dp.rf.reg_file_arr[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30156_ (.CLK(_00691_),
    .D(_01891_),
    .Q(\rvcpu.dp.rf.reg_file_arr[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30157_ (.CLK(_00692_),
    .D(_01892_),
    .Q(\rvcpu.dp.rf.reg_file_arr[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _30158_ (.CLK(_00693_),
    .D(_01893_),
    .Q(\rvcpu.dp.rf.reg_file_arr[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _30159_ (.CLK(_00694_),
    .D(_01894_),
    .Q(\rvcpu.dp.rf.reg_file_arr[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _30160_ (.CLK(_00695_),
    .D(_01895_),
    .Q(\rvcpu.dp.rf.reg_file_arr[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _30161_ (.CLK(_00696_),
    .D(_01896_),
    .Q(\rvcpu.dp.rf.reg_file_arr[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _30162_ (.CLK(_00697_),
    .D(_01897_),
    .Q(\rvcpu.dp.rf.reg_file_arr[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _30163_ (.CLK(_00698_),
    .D(_01898_),
    .Q(\rvcpu.dp.rf.reg_file_arr[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _30164_ (.CLK(_00699_),
    .D(_01899_),
    .Q(\rvcpu.dp.rf.reg_file_arr[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _30165_ (.CLK(_00700_),
    .D(_01900_),
    .Q(\rvcpu.dp.rf.reg_file_arr[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _30166_ (.CLK(_00701_),
    .D(_01901_),
    .Q(\rvcpu.dp.rf.reg_file_arr[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _30167_ (.CLK(_00702_),
    .D(_01902_),
    .Q(\rvcpu.dp.rf.reg_file_arr[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _30168_ (.CLK(_00703_),
    .D(_01903_),
    .Q(\rvcpu.dp.rf.reg_file_arr[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _30169_ (.CLK(_00704_),
    .D(_01904_),
    .Q(\rvcpu.dp.rf.reg_file_arr[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _30170_ (.CLK(_00705_),
    .D(_01905_),
    .Q(\rvcpu.dp.rf.reg_file_arr[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _30171_ (.CLK(_00706_),
    .D(_01906_),
    .Q(\rvcpu.dp.rf.reg_file_arr[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _30172_ (.CLK(_00707_),
    .D(_01907_),
    .Q(\rvcpu.dp.rf.reg_file_arr[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _30173_ (.CLK(clk),
    .D(_01908_),
    .Q(\datamem.data_ram[58][24] ));
 sky130_fd_sc_hd__dfxtp_1 _30174_ (.CLK(clk),
    .D(_01909_),
    .Q(\datamem.data_ram[58][25] ));
 sky130_fd_sc_hd__dfxtp_1 _30175_ (.CLK(clk),
    .D(_01910_),
    .Q(\datamem.data_ram[58][26] ));
 sky130_fd_sc_hd__dfxtp_1 _30176_ (.CLK(clk),
    .D(_01911_),
    .Q(\datamem.data_ram[58][27] ));
 sky130_fd_sc_hd__dfxtp_1 _30177_ (.CLK(clk),
    .D(_01912_),
    .Q(\datamem.data_ram[58][28] ));
 sky130_fd_sc_hd__dfxtp_1 _30178_ (.CLK(clk),
    .D(_01913_),
    .Q(\datamem.data_ram[58][29] ));
 sky130_fd_sc_hd__dfxtp_1 _30179_ (.CLK(clk),
    .D(_01914_),
    .Q(\datamem.data_ram[58][30] ));
 sky130_fd_sc_hd__dfxtp_1 _30180_ (.CLK(clk),
    .D(_01915_),
    .Q(\datamem.data_ram[58][31] ));
 sky130_fd_sc_hd__dfxtp_1 _30181_ (.CLK(_00708_),
    .D(_01916_),
    .Q(\rvcpu.dp.rf.reg_file_arr[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _30182_ (.CLK(_00709_),
    .D(_01917_),
    .Q(\rvcpu.dp.rf.reg_file_arr[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _30183_ (.CLK(_00710_),
    .D(_01918_),
    .Q(\rvcpu.dp.rf.reg_file_arr[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _30184_ (.CLK(_00711_),
    .D(_01919_),
    .Q(\rvcpu.dp.rf.reg_file_arr[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _30185_ (.CLK(_00712_),
    .D(_01920_),
    .Q(\rvcpu.dp.rf.reg_file_arr[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _30186_ (.CLK(_00713_),
    .D(_01921_),
    .Q(\rvcpu.dp.rf.reg_file_arr[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _30187_ (.CLK(_00714_),
    .D(_01922_),
    .Q(\rvcpu.dp.rf.reg_file_arr[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _30188_ (.CLK(_00715_),
    .D(_01923_),
    .Q(\rvcpu.dp.rf.reg_file_arr[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _30189_ (.CLK(_00716_),
    .D(_01924_),
    .Q(\rvcpu.dp.rf.reg_file_arr[8][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30190_ (.CLK(_00717_),
    .D(_01925_),
    .Q(\rvcpu.dp.rf.reg_file_arr[8][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30191_ (.CLK(_00718_),
    .D(_01926_),
    .Q(\rvcpu.dp.rf.reg_file_arr[8][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30192_ (.CLK(_00719_),
    .D(_01927_),
    .Q(\rvcpu.dp.rf.reg_file_arr[8][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30193_ (.CLK(_00720_),
    .D(_01928_),
    .Q(\rvcpu.dp.rf.reg_file_arr[8][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30194_ (.CLK(_00721_),
    .D(_01929_),
    .Q(\rvcpu.dp.rf.reg_file_arr[8][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30195_ (.CLK(_00722_),
    .D(_01930_),
    .Q(\rvcpu.dp.rf.reg_file_arr[8][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30196_ (.CLK(_00723_),
    .D(_01931_),
    .Q(\rvcpu.dp.rf.reg_file_arr[8][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30197_ (.CLK(_00724_),
    .D(_01932_),
    .Q(\rvcpu.dp.rf.reg_file_arr[8][16] ));
 sky130_fd_sc_hd__dfxtp_1 _30198_ (.CLK(_00725_),
    .D(_01933_),
    .Q(\rvcpu.dp.rf.reg_file_arr[8][17] ));
 sky130_fd_sc_hd__dfxtp_1 _30199_ (.CLK(_00726_),
    .D(_01934_),
    .Q(\rvcpu.dp.rf.reg_file_arr[8][18] ));
 sky130_fd_sc_hd__dfxtp_1 _30200_ (.CLK(_00727_),
    .D(_01935_),
    .Q(\rvcpu.dp.rf.reg_file_arr[8][19] ));
 sky130_fd_sc_hd__dfxtp_1 _30201_ (.CLK(_00728_),
    .D(_01936_),
    .Q(\rvcpu.dp.rf.reg_file_arr[8][20] ));
 sky130_fd_sc_hd__dfxtp_1 _30202_ (.CLK(_00729_),
    .D(_01937_),
    .Q(\rvcpu.dp.rf.reg_file_arr[8][21] ));
 sky130_fd_sc_hd__dfxtp_1 _30203_ (.CLK(_00730_),
    .D(_01938_),
    .Q(\rvcpu.dp.rf.reg_file_arr[8][22] ));
 sky130_fd_sc_hd__dfxtp_1 _30204_ (.CLK(_00731_),
    .D(_01939_),
    .Q(\rvcpu.dp.rf.reg_file_arr[8][23] ));
 sky130_fd_sc_hd__dfxtp_1 _30205_ (.CLK(_00732_),
    .D(_01940_),
    .Q(\rvcpu.dp.rf.reg_file_arr[8][24] ));
 sky130_fd_sc_hd__dfxtp_1 _30206_ (.CLK(_00733_),
    .D(_01941_),
    .Q(\rvcpu.dp.rf.reg_file_arr[8][25] ));
 sky130_fd_sc_hd__dfxtp_1 _30207_ (.CLK(_00734_),
    .D(_01942_),
    .Q(\rvcpu.dp.rf.reg_file_arr[8][26] ));
 sky130_fd_sc_hd__dfxtp_1 _30208_ (.CLK(_00735_),
    .D(_01943_),
    .Q(\rvcpu.dp.rf.reg_file_arr[8][27] ));
 sky130_fd_sc_hd__dfxtp_1 _30209_ (.CLK(_00736_),
    .D(_01944_),
    .Q(\rvcpu.dp.rf.reg_file_arr[8][28] ));
 sky130_fd_sc_hd__dfxtp_1 _30210_ (.CLK(_00737_),
    .D(_01945_),
    .Q(\rvcpu.dp.rf.reg_file_arr[8][29] ));
 sky130_fd_sc_hd__dfxtp_1 _30211_ (.CLK(_00738_),
    .D(_01946_),
    .Q(\rvcpu.dp.rf.reg_file_arr[8][30] ));
 sky130_fd_sc_hd__dfxtp_1 _30212_ (.CLK(_00739_),
    .D(_01947_),
    .Q(\rvcpu.dp.rf.reg_file_arr[8][31] ));
 sky130_fd_sc_hd__dfxtp_1 _30213_ (.CLK(_00740_),
    .D(_01948_),
    .Q(\rvcpu.dp.rf.reg_file_arr[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _30214_ (.CLK(_00741_),
    .D(_01949_),
    .Q(\rvcpu.dp.rf.reg_file_arr[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _30215_ (.CLK(_00742_),
    .D(_01950_),
    .Q(\rvcpu.dp.rf.reg_file_arr[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _30216_ (.CLK(_00743_),
    .D(_01951_),
    .Q(\rvcpu.dp.rf.reg_file_arr[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _30217_ (.CLK(_00744_),
    .D(_01952_),
    .Q(\rvcpu.dp.rf.reg_file_arr[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _30218_ (.CLK(_00745_),
    .D(_01953_),
    .Q(\rvcpu.dp.rf.reg_file_arr[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _30219_ (.CLK(_00746_),
    .D(_01954_),
    .Q(\rvcpu.dp.rf.reg_file_arr[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _30220_ (.CLK(_00747_),
    .D(_01955_),
    .Q(\rvcpu.dp.rf.reg_file_arr[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _30221_ (.CLK(_00748_),
    .D(_01956_),
    .Q(\rvcpu.dp.rf.reg_file_arr[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30222_ (.CLK(_00749_),
    .D(_01957_),
    .Q(\rvcpu.dp.rf.reg_file_arr[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30223_ (.CLK(_00750_),
    .D(_01958_),
    .Q(\rvcpu.dp.rf.reg_file_arr[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30224_ (.CLK(_00751_),
    .D(_01959_),
    .Q(\rvcpu.dp.rf.reg_file_arr[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30225_ (.CLK(_00752_),
    .D(_01960_),
    .Q(\rvcpu.dp.rf.reg_file_arr[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30226_ (.CLK(_00753_),
    .D(_01961_),
    .Q(\rvcpu.dp.rf.reg_file_arr[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30227_ (.CLK(_00754_),
    .D(_01962_),
    .Q(\rvcpu.dp.rf.reg_file_arr[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30228_ (.CLK(_00755_),
    .D(_01963_),
    .Q(\rvcpu.dp.rf.reg_file_arr[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30229_ (.CLK(_00756_),
    .D(_01964_),
    .Q(\rvcpu.dp.rf.reg_file_arr[7][16] ));
 sky130_fd_sc_hd__dfxtp_1 _30230_ (.CLK(_00757_),
    .D(_01965_),
    .Q(\rvcpu.dp.rf.reg_file_arr[7][17] ));
 sky130_fd_sc_hd__dfxtp_1 _30231_ (.CLK(_00758_),
    .D(_01966_),
    .Q(\rvcpu.dp.rf.reg_file_arr[7][18] ));
 sky130_fd_sc_hd__dfxtp_1 _30232_ (.CLK(_00759_),
    .D(_01967_),
    .Q(\rvcpu.dp.rf.reg_file_arr[7][19] ));
 sky130_fd_sc_hd__dfxtp_1 _30233_ (.CLK(_00760_),
    .D(_01968_),
    .Q(\rvcpu.dp.rf.reg_file_arr[7][20] ));
 sky130_fd_sc_hd__dfxtp_1 _30234_ (.CLK(_00761_),
    .D(_01969_),
    .Q(\rvcpu.dp.rf.reg_file_arr[7][21] ));
 sky130_fd_sc_hd__dfxtp_1 _30235_ (.CLK(_00762_),
    .D(_01970_),
    .Q(\rvcpu.dp.rf.reg_file_arr[7][22] ));
 sky130_fd_sc_hd__dfxtp_1 _30236_ (.CLK(_00763_),
    .D(_01971_),
    .Q(\rvcpu.dp.rf.reg_file_arr[7][23] ));
 sky130_fd_sc_hd__dfxtp_1 _30237_ (.CLK(_00764_),
    .D(_01972_),
    .Q(\rvcpu.dp.rf.reg_file_arr[7][24] ));
 sky130_fd_sc_hd__dfxtp_1 _30238_ (.CLK(_00765_),
    .D(_01973_),
    .Q(\rvcpu.dp.rf.reg_file_arr[7][25] ));
 sky130_fd_sc_hd__dfxtp_1 _30239_ (.CLK(_00766_),
    .D(_01974_),
    .Q(\rvcpu.dp.rf.reg_file_arr[7][26] ));
 sky130_fd_sc_hd__dfxtp_1 _30240_ (.CLK(_00767_),
    .D(_01975_),
    .Q(\rvcpu.dp.rf.reg_file_arr[7][27] ));
 sky130_fd_sc_hd__dfxtp_1 _30241_ (.CLK(_00768_),
    .D(_01976_),
    .Q(\rvcpu.dp.rf.reg_file_arr[7][28] ));
 sky130_fd_sc_hd__dfxtp_1 _30242_ (.CLK(_00769_),
    .D(_01977_),
    .Q(\rvcpu.dp.rf.reg_file_arr[7][29] ));
 sky130_fd_sc_hd__dfxtp_1 _30243_ (.CLK(_00770_),
    .D(_01978_),
    .Q(\rvcpu.dp.rf.reg_file_arr[7][30] ));
 sky130_fd_sc_hd__dfxtp_1 _30244_ (.CLK(_00771_),
    .D(_01979_),
    .Q(\rvcpu.dp.rf.reg_file_arr[7][31] ));
 sky130_fd_sc_hd__dfxtp_1 _30245_ (.CLK(_00772_),
    .D(_01980_),
    .Q(\rvcpu.dp.rf.reg_file_arr[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _30246_ (.CLK(_00773_),
    .D(_01981_),
    .Q(\rvcpu.dp.rf.reg_file_arr[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _30247_ (.CLK(_00774_),
    .D(_01982_),
    .Q(\rvcpu.dp.rf.reg_file_arr[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _30248_ (.CLK(_00775_),
    .D(_01983_),
    .Q(\rvcpu.dp.rf.reg_file_arr[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _30249_ (.CLK(_00776_),
    .D(_01984_),
    .Q(\rvcpu.dp.rf.reg_file_arr[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _30250_ (.CLK(_00777_),
    .D(_01985_),
    .Q(\rvcpu.dp.rf.reg_file_arr[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _30251_ (.CLK(_00778_),
    .D(_01986_),
    .Q(\rvcpu.dp.rf.reg_file_arr[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _30252_ (.CLK(_00779_),
    .D(_01987_),
    .Q(\rvcpu.dp.rf.reg_file_arr[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _30253_ (.CLK(_00780_),
    .D(_01988_),
    .Q(\rvcpu.dp.rf.reg_file_arr[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30254_ (.CLK(_00781_),
    .D(_01989_),
    .Q(\rvcpu.dp.rf.reg_file_arr[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30255_ (.CLK(_00782_),
    .D(_01990_),
    .Q(\rvcpu.dp.rf.reg_file_arr[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30256_ (.CLK(_00783_),
    .D(_01991_),
    .Q(\rvcpu.dp.rf.reg_file_arr[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30257_ (.CLK(_00784_),
    .D(_01992_),
    .Q(\rvcpu.dp.rf.reg_file_arr[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30258_ (.CLK(_00785_),
    .D(_01993_),
    .Q(\rvcpu.dp.rf.reg_file_arr[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30259_ (.CLK(_00786_),
    .D(_01994_),
    .Q(\rvcpu.dp.rf.reg_file_arr[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30260_ (.CLK(_00787_),
    .D(_01995_),
    .Q(\rvcpu.dp.rf.reg_file_arr[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30261_ (.CLK(_00788_),
    .D(_01996_),
    .Q(\rvcpu.dp.rf.reg_file_arr[6][16] ));
 sky130_fd_sc_hd__dfxtp_1 _30262_ (.CLK(_00789_),
    .D(_01997_),
    .Q(\rvcpu.dp.rf.reg_file_arr[6][17] ));
 sky130_fd_sc_hd__dfxtp_1 _30263_ (.CLK(_00790_),
    .D(_01998_),
    .Q(\rvcpu.dp.rf.reg_file_arr[6][18] ));
 sky130_fd_sc_hd__dfxtp_1 _30264_ (.CLK(_00791_),
    .D(_01999_),
    .Q(\rvcpu.dp.rf.reg_file_arr[6][19] ));
 sky130_fd_sc_hd__dfxtp_1 _30265_ (.CLK(_00792_),
    .D(_02000_),
    .Q(\rvcpu.dp.rf.reg_file_arr[6][20] ));
 sky130_fd_sc_hd__dfxtp_1 _30266_ (.CLK(_00793_),
    .D(_02001_),
    .Q(\rvcpu.dp.rf.reg_file_arr[6][21] ));
 sky130_fd_sc_hd__dfxtp_1 _30267_ (.CLK(_00794_),
    .D(_02002_),
    .Q(\rvcpu.dp.rf.reg_file_arr[6][22] ));
 sky130_fd_sc_hd__dfxtp_1 _30268_ (.CLK(_00795_),
    .D(_02003_),
    .Q(\rvcpu.dp.rf.reg_file_arr[6][23] ));
 sky130_fd_sc_hd__dfxtp_1 _30269_ (.CLK(_00796_),
    .D(_02004_),
    .Q(\rvcpu.dp.rf.reg_file_arr[6][24] ));
 sky130_fd_sc_hd__dfxtp_1 _30270_ (.CLK(_00797_),
    .D(_02005_),
    .Q(\rvcpu.dp.rf.reg_file_arr[6][25] ));
 sky130_fd_sc_hd__dfxtp_1 _30271_ (.CLK(_00798_),
    .D(_02006_),
    .Q(\rvcpu.dp.rf.reg_file_arr[6][26] ));
 sky130_fd_sc_hd__dfxtp_1 _30272_ (.CLK(_00799_),
    .D(_02007_),
    .Q(\rvcpu.dp.rf.reg_file_arr[6][27] ));
 sky130_fd_sc_hd__dfxtp_1 _30273_ (.CLK(_00800_),
    .D(_02008_),
    .Q(\rvcpu.dp.rf.reg_file_arr[6][28] ));
 sky130_fd_sc_hd__dfxtp_1 _30274_ (.CLK(_00801_),
    .D(_02009_),
    .Q(\rvcpu.dp.rf.reg_file_arr[6][29] ));
 sky130_fd_sc_hd__dfxtp_1 _30275_ (.CLK(_00802_),
    .D(_02010_),
    .Q(\rvcpu.dp.rf.reg_file_arr[6][30] ));
 sky130_fd_sc_hd__dfxtp_1 _30276_ (.CLK(_00803_),
    .D(_02011_),
    .Q(\rvcpu.dp.rf.reg_file_arr[6][31] ));
 sky130_fd_sc_hd__dfxtp_1 _30277_ (.CLK(clk),
    .D(_02012_),
    .Q(\datamem.data_ram[58][16] ));
 sky130_fd_sc_hd__dfxtp_1 _30278_ (.CLK(clk),
    .D(_02013_),
    .Q(\datamem.data_ram[58][17] ));
 sky130_fd_sc_hd__dfxtp_1 _30279_ (.CLK(clk),
    .D(_02014_),
    .Q(\datamem.data_ram[58][18] ));
 sky130_fd_sc_hd__dfxtp_1 _30280_ (.CLK(clk),
    .D(_02015_),
    .Q(\datamem.data_ram[58][19] ));
 sky130_fd_sc_hd__dfxtp_1 _30281_ (.CLK(clk),
    .D(_02016_),
    .Q(\datamem.data_ram[58][20] ));
 sky130_fd_sc_hd__dfxtp_1 _30282_ (.CLK(clk),
    .D(_02017_),
    .Q(\datamem.data_ram[58][21] ));
 sky130_fd_sc_hd__dfxtp_1 _30283_ (.CLK(clk),
    .D(_02018_),
    .Q(\datamem.data_ram[58][22] ));
 sky130_fd_sc_hd__dfxtp_1 _30284_ (.CLK(clk),
    .D(_02019_),
    .Q(\datamem.data_ram[58][23] ));
 sky130_fd_sc_hd__dfxtp_1 _30285_ (.CLK(_00804_),
    .D(_02020_),
    .Q(\rvcpu.dp.rf.reg_file_arr[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _30286_ (.CLK(_00805_),
    .D(_02021_),
    .Q(\rvcpu.dp.rf.reg_file_arr[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _30287_ (.CLK(_00806_),
    .D(_02022_),
    .Q(\rvcpu.dp.rf.reg_file_arr[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _30288_ (.CLK(_00807_),
    .D(_02023_),
    .Q(\rvcpu.dp.rf.reg_file_arr[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _30289_ (.CLK(_00808_),
    .D(_02024_),
    .Q(\rvcpu.dp.rf.reg_file_arr[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _30290_ (.CLK(_00809_),
    .D(_02025_),
    .Q(\rvcpu.dp.rf.reg_file_arr[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _30291_ (.CLK(_00810_),
    .D(_02026_),
    .Q(\rvcpu.dp.rf.reg_file_arr[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _30292_ (.CLK(_00811_),
    .D(_02027_),
    .Q(\rvcpu.dp.rf.reg_file_arr[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _30293_ (.CLK(_00812_),
    .D(_02028_),
    .Q(\rvcpu.dp.rf.reg_file_arr[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30294_ (.CLK(_00813_),
    .D(_02029_),
    .Q(\rvcpu.dp.rf.reg_file_arr[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30295_ (.CLK(_00814_),
    .D(_02030_),
    .Q(\rvcpu.dp.rf.reg_file_arr[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30296_ (.CLK(_00815_),
    .D(_02031_),
    .Q(\rvcpu.dp.rf.reg_file_arr[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30297_ (.CLK(_00816_),
    .D(_02032_),
    .Q(\rvcpu.dp.rf.reg_file_arr[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30298_ (.CLK(_00817_),
    .D(_02033_),
    .Q(\rvcpu.dp.rf.reg_file_arr[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30299_ (.CLK(_00818_),
    .D(_02034_),
    .Q(\rvcpu.dp.rf.reg_file_arr[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30300_ (.CLK(_00819_),
    .D(_02035_),
    .Q(\rvcpu.dp.rf.reg_file_arr[5][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30301_ (.CLK(_00820_),
    .D(_02036_),
    .Q(\rvcpu.dp.rf.reg_file_arr[5][16] ));
 sky130_fd_sc_hd__dfxtp_1 _30302_ (.CLK(_00821_),
    .D(_02037_),
    .Q(\rvcpu.dp.rf.reg_file_arr[5][17] ));
 sky130_fd_sc_hd__dfxtp_1 _30303_ (.CLK(_00822_),
    .D(_02038_),
    .Q(\rvcpu.dp.rf.reg_file_arr[5][18] ));
 sky130_fd_sc_hd__dfxtp_1 _30304_ (.CLK(_00823_),
    .D(_02039_),
    .Q(\rvcpu.dp.rf.reg_file_arr[5][19] ));
 sky130_fd_sc_hd__dfxtp_1 _30305_ (.CLK(_00824_),
    .D(_02040_),
    .Q(\rvcpu.dp.rf.reg_file_arr[5][20] ));
 sky130_fd_sc_hd__dfxtp_1 _30306_ (.CLK(_00825_),
    .D(_02041_),
    .Q(\rvcpu.dp.rf.reg_file_arr[5][21] ));
 sky130_fd_sc_hd__dfxtp_1 _30307_ (.CLK(_00826_),
    .D(_02042_),
    .Q(\rvcpu.dp.rf.reg_file_arr[5][22] ));
 sky130_fd_sc_hd__dfxtp_1 _30308_ (.CLK(_00827_),
    .D(_02043_),
    .Q(\rvcpu.dp.rf.reg_file_arr[5][23] ));
 sky130_fd_sc_hd__dfxtp_1 _30309_ (.CLK(_00828_),
    .D(_02044_),
    .Q(\rvcpu.dp.rf.reg_file_arr[5][24] ));
 sky130_fd_sc_hd__dfxtp_1 _30310_ (.CLK(_00829_),
    .D(_02045_),
    .Q(\rvcpu.dp.rf.reg_file_arr[5][25] ));
 sky130_fd_sc_hd__dfxtp_1 _30311_ (.CLK(_00830_),
    .D(_02046_),
    .Q(\rvcpu.dp.rf.reg_file_arr[5][26] ));
 sky130_fd_sc_hd__dfxtp_1 _30312_ (.CLK(_00831_),
    .D(_02047_),
    .Q(\rvcpu.dp.rf.reg_file_arr[5][27] ));
 sky130_fd_sc_hd__dfxtp_1 _30313_ (.CLK(_00832_),
    .D(_02048_),
    .Q(\rvcpu.dp.rf.reg_file_arr[5][28] ));
 sky130_fd_sc_hd__dfxtp_1 _30314_ (.CLK(_00833_),
    .D(_02049_),
    .Q(\rvcpu.dp.rf.reg_file_arr[5][29] ));
 sky130_fd_sc_hd__dfxtp_1 _30315_ (.CLK(_00834_),
    .D(_02050_),
    .Q(\rvcpu.dp.rf.reg_file_arr[5][30] ));
 sky130_fd_sc_hd__dfxtp_1 _30316_ (.CLK(_00835_),
    .D(_02051_),
    .Q(\rvcpu.dp.rf.reg_file_arr[5][31] ));
 sky130_fd_sc_hd__dfxtp_1 _30317_ (.CLK(_00836_),
    .D(_02052_),
    .Q(\rvcpu.dp.rf.reg_file_arr[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _30318_ (.CLK(_00837_),
    .D(_02053_),
    .Q(\rvcpu.dp.rf.reg_file_arr[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _30319_ (.CLK(_00838_),
    .D(_02054_),
    .Q(\rvcpu.dp.rf.reg_file_arr[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _30320_ (.CLK(_00839_),
    .D(_02055_),
    .Q(\rvcpu.dp.rf.reg_file_arr[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _30321_ (.CLK(_00840_),
    .D(_02056_),
    .Q(\rvcpu.dp.rf.reg_file_arr[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _30322_ (.CLK(_00841_),
    .D(_02057_),
    .Q(\rvcpu.dp.rf.reg_file_arr[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _30323_ (.CLK(_00842_),
    .D(_02058_),
    .Q(\rvcpu.dp.rf.reg_file_arr[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _30324_ (.CLK(_00843_),
    .D(_02059_),
    .Q(\rvcpu.dp.rf.reg_file_arr[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _30325_ (.CLK(_00844_),
    .D(_02060_),
    .Q(\rvcpu.dp.rf.reg_file_arr[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30326_ (.CLK(_00845_),
    .D(_02061_),
    .Q(\rvcpu.dp.rf.reg_file_arr[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30327_ (.CLK(_00846_),
    .D(_02062_),
    .Q(\rvcpu.dp.rf.reg_file_arr[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30328_ (.CLK(_00847_),
    .D(_02063_),
    .Q(\rvcpu.dp.rf.reg_file_arr[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30329_ (.CLK(_00848_),
    .D(_02064_),
    .Q(\rvcpu.dp.rf.reg_file_arr[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30330_ (.CLK(_00849_),
    .D(_02065_),
    .Q(\rvcpu.dp.rf.reg_file_arr[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30331_ (.CLK(_00850_),
    .D(_02066_),
    .Q(\rvcpu.dp.rf.reg_file_arr[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30332_ (.CLK(_00851_),
    .D(_02067_),
    .Q(\rvcpu.dp.rf.reg_file_arr[4][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30333_ (.CLK(_00852_),
    .D(_02068_),
    .Q(\rvcpu.dp.rf.reg_file_arr[4][16] ));
 sky130_fd_sc_hd__dfxtp_1 _30334_ (.CLK(_00853_),
    .D(_02069_),
    .Q(\rvcpu.dp.rf.reg_file_arr[4][17] ));
 sky130_fd_sc_hd__dfxtp_1 _30335_ (.CLK(_00854_),
    .D(_02070_),
    .Q(\rvcpu.dp.rf.reg_file_arr[4][18] ));
 sky130_fd_sc_hd__dfxtp_1 _30336_ (.CLK(_00855_),
    .D(_02071_),
    .Q(\rvcpu.dp.rf.reg_file_arr[4][19] ));
 sky130_fd_sc_hd__dfxtp_1 _30337_ (.CLK(_00856_),
    .D(_02072_),
    .Q(\rvcpu.dp.rf.reg_file_arr[4][20] ));
 sky130_fd_sc_hd__dfxtp_1 _30338_ (.CLK(_00857_),
    .D(_02073_),
    .Q(\rvcpu.dp.rf.reg_file_arr[4][21] ));
 sky130_fd_sc_hd__dfxtp_1 _30339_ (.CLK(_00858_),
    .D(_02074_),
    .Q(\rvcpu.dp.rf.reg_file_arr[4][22] ));
 sky130_fd_sc_hd__dfxtp_1 _30340_ (.CLK(_00859_),
    .D(_02075_),
    .Q(\rvcpu.dp.rf.reg_file_arr[4][23] ));
 sky130_fd_sc_hd__dfxtp_1 _30341_ (.CLK(_00860_),
    .D(_02076_),
    .Q(\rvcpu.dp.rf.reg_file_arr[4][24] ));
 sky130_fd_sc_hd__dfxtp_1 _30342_ (.CLK(_00861_),
    .D(_02077_),
    .Q(\rvcpu.dp.rf.reg_file_arr[4][25] ));
 sky130_fd_sc_hd__dfxtp_1 _30343_ (.CLK(_00862_),
    .D(_02078_),
    .Q(\rvcpu.dp.rf.reg_file_arr[4][26] ));
 sky130_fd_sc_hd__dfxtp_1 _30344_ (.CLK(_00863_),
    .D(_02079_),
    .Q(\rvcpu.dp.rf.reg_file_arr[4][27] ));
 sky130_fd_sc_hd__dfxtp_1 _30345_ (.CLK(_00864_),
    .D(_02080_),
    .Q(\rvcpu.dp.rf.reg_file_arr[4][28] ));
 sky130_fd_sc_hd__dfxtp_1 _30346_ (.CLK(_00865_),
    .D(_02081_),
    .Q(\rvcpu.dp.rf.reg_file_arr[4][29] ));
 sky130_fd_sc_hd__dfxtp_1 _30347_ (.CLK(_00866_),
    .D(_02082_),
    .Q(\rvcpu.dp.rf.reg_file_arr[4][30] ));
 sky130_fd_sc_hd__dfxtp_1 _30348_ (.CLK(_00867_),
    .D(_02083_),
    .Q(\rvcpu.dp.rf.reg_file_arr[4][31] ));
 sky130_fd_sc_hd__dfxtp_1 _30349_ (.CLK(_00868_),
    .D(_02084_),
    .Q(\rvcpu.dp.rf.reg_file_arr[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _30350_ (.CLK(_00869_),
    .D(_02085_),
    .Q(\rvcpu.dp.rf.reg_file_arr[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _30351_ (.CLK(_00870_),
    .D(_02086_),
    .Q(\rvcpu.dp.rf.reg_file_arr[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _30352_ (.CLK(_00871_),
    .D(_02087_),
    .Q(\rvcpu.dp.rf.reg_file_arr[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _30353_ (.CLK(_00872_),
    .D(_02088_),
    .Q(\rvcpu.dp.rf.reg_file_arr[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _30354_ (.CLK(_00873_),
    .D(_02089_),
    .Q(\rvcpu.dp.rf.reg_file_arr[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _30355_ (.CLK(_00874_),
    .D(_02090_),
    .Q(\rvcpu.dp.rf.reg_file_arr[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _30356_ (.CLK(_00875_),
    .D(_02091_),
    .Q(\rvcpu.dp.rf.reg_file_arr[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _30357_ (.CLK(_00876_),
    .D(_02092_),
    .Q(\rvcpu.dp.rf.reg_file_arr[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30358_ (.CLK(_00877_),
    .D(_02093_),
    .Q(\rvcpu.dp.rf.reg_file_arr[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30359_ (.CLK(_00878_),
    .D(_02094_),
    .Q(\rvcpu.dp.rf.reg_file_arr[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30360_ (.CLK(_00879_),
    .D(_02095_),
    .Q(\rvcpu.dp.rf.reg_file_arr[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30361_ (.CLK(_00880_),
    .D(_02096_),
    .Q(\rvcpu.dp.rf.reg_file_arr[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30362_ (.CLK(_00881_),
    .D(_02097_),
    .Q(\rvcpu.dp.rf.reg_file_arr[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30363_ (.CLK(_00882_),
    .D(_02098_),
    .Q(\rvcpu.dp.rf.reg_file_arr[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30364_ (.CLK(_00883_),
    .D(_02099_),
    .Q(\rvcpu.dp.rf.reg_file_arr[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30365_ (.CLK(_00884_),
    .D(_02100_),
    .Q(\rvcpu.dp.rf.reg_file_arr[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 _30366_ (.CLK(_00885_),
    .D(_02101_),
    .Q(\rvcpu.dp.rf.reg_file_arr[3][17] ));
 sky130_fd_sc_hd__dfxtp_1 _30367_ (.CLK(_00886_),
    .D(_02102_),
    .Q(\rvcpu.dp.rf.reg_file_arr[3][18] ));
 sky130_fd_sc_hd__dfxtp_1 _30368_ (.CLK(_00887_),
    .D(_02103_),
    .Q(\rvcpu.dp.rf.reg_file_arr[3][19] ));
 sky130_fd_sc_hd__dfxtp_1 _30369_ (.CLK(_00888_),
    .D(_02104_),
    .Q(\rvcpu.dp.rf.reg_file_arr[3][20] ));
 sky130_fd_sc_hd__dfxtp_1 _30370_ (.CLK(_00889_),
    .D(_02105_),
    .Q(\rvcpu.dp.rf.reg_file_arr[3][21] ));
 sky130_fd_sc_hd__dfxtp_1 _30371_ (.CLK(_00890_),
    .D(_02106_),
    .Q(\rvcpu.dp.rf.reg_file_arr[3][22] ));
 sky130_fd_sc_hd__dfxtp_1 _30372_ (.CLK(_00891_),
    .D(_02107_),
    .Q(\rvcpu.dp.rf.reg_file_arr[3][23] ));
 sky130_fd_sc_hd__dfxtp_1 _30373_ (.CLK(_00892_),
    .D(_02108_),
    .Q(\rvcpu.dp.rf.reg_file_arr[3][24] ));
 sky130_fd_sc_hd__dfxtp_1 _30374_ (.CLK(_00893_),
    .D(_02109_),
    .Q(\rvcpu.dp.rf.reg_file_arr[3][25] ));
 sky130_fd_sc_hd__dfxtp_1 _30375_ (.CLK(_00894_),
    .D(_02110_),
    .Q(\rvcpu.dp.rf.reg_file_arr[3][26] ));
 sky130_fd_sc_hd__dfxtp_1 _30376_ (.CLK(_00895_),
    .D(_02111_),
    .Q(\rvcpu.dp.rf.reg_file_arr[3][27] ));
 sky130_fd_sc_hd__dfxtp_1 _30377_ (.CLK(_00896_),
    .D(_02112_),
    .Q(\rvcpu.dp.rf.reg_file_arr[3][28] ));
 sky130_fd_sc_hd__dfxtp_1 _30378_ (.CLK(_00897_),
    .D(_02113_),
    .Q(\rvcpu.dp.rf.reg_file_arr[3][29] ));
 sky130_fd_sc_hd__dfxtp_1 _30379_ (.CLK(_00898_),
    .D(_02114_),
    .Q(\rvcpu.dp.rf.reg_file_arr[3][30] ));
 sky130_fd_sc_hd__dfxtp_1 _30380_ (.CLK(_00899_),
    .D(_02115_),
    .Q(\rvcpu.dp.rf.reg_file_arr[3][31] ));
 sky130_fd_sc_hd__dfxtp_1 _30381_ (.CLK(clk),
    .D(_02116_),
    .Q(\datamem.data_ram[58][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30382_ (.CLK(clk),
    .D(_02117_),
    .Q(\datamem.data_ram[58][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30383_ (.CLK(clk),
    .D(_02118_),
    .Q(\datamem.data_ram[58][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30384_ (.CLK(clk),
    .D(_02119_),
    .Q(\datamem.data_ram[58][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30385_ (.CLK(clk),
    .D(_02120_),
    .Q(\datamem.data_ram[58][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30386_ (.CLK(clk),
    .D(_02121_),
    .Q(\datamem.data_ram[58][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30387_ (.CLK(clk),
    .D(_02122_),
    .Q(\datamem.data_ram[58][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30388_ (.CLK(clk),
    .D(_02123_),
    .Q(\datamem.data_ram[58][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30389_ (.CLK(_00900_),
    .D(_02124_),
    .Q(\rvcpu.dp.rf.reg_file_arr[31][0] ));
 sky130_fd_sc_hd__dfxtp_1 _30390_ (.CLK(_00901_),
    .D(_02125_),
    .Q(\rvcpu.dp.rf.reg_file_arr[31][1] ));
 sky130_fd_sc_hd__dfxtp_1 _30391_ (.CLK(_00902_),
    .D(_02126_),
    .Q(\rvcpu.dp.rf.reg_file_arr[31][2] ));
 sky130_fd_sc_hd__dfxtp_1 _30392_ (.CLK(_00903_),
    .D(_02127_),
    .Q(\rvcpu.dp.rf.reg_file_arr[31][3] ));
 sky130_fd_sc_hd__dfxtp_1 _30393_ (.CLK(_00904_),
    .D(_02128_),
    .Q(\rvcpu.dp.rf.reg_file_arr[31][4] ));
 sky130_fd_sc_hd__dfxtp_1 _30394_ (.CLK(_00905_),
    .D(_02129_),
    .Q(\rvcpu.dp.rf.reg_file_arr[31][5] ));
 sky130_fd_sc_hd__dfxtp_1 _30395_ (.CLK(_00906_),
    .D(_02130_),
    .Q(\rvcpu.dp.rf.reg_file_arr[31][6] ));
 sky130_fd_sc_hd__dfxtp_1 _30396_ (.CLK(_00907_),
    .D(_02131_),
    .Q(\rvcpu.dp.rf.reg_file_arr[31][7] ));
 sky130_fd_sc_hd__dfxtp_1 _30397_ (.CLK(_00908_),
    .D(_02132_),
    .Q(\rvcpu.dp.rf.reg_file_arr[31][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30398_ (.CLK(_00909_),
    .D(_02133_),
    .Q(\rvcpu.dp.rf.reg_file_arr[31][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30399_ (.CLK(_00910_),
    .D(_02134_),
    .Q(\rvcpu.dp.rf.reg_file_arr[31][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30400_ (.CLK(_00911_),
    .D(_02135_),
    .Q(\rvcpu.dp.rf.reg_file_arr[31][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30401_ (.CLK(_00912_),
    .D(_02136_),
    .Q(\rvcpu.dp.rf.reg_file_arr[31][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30402_ (.CLK(_00913_),
    .D(_02137_),
    .Q(\rvcpu.dp.rf.reg_file_arr[31][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30403_ (.CLK(_00914_),
    .D(_02138_),
    .Q(\rvcpu.dp.rf.reg_file_arr[31][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30404_ (.CLK(_00915_),
    .D(_02139_),
    .Q(\rvcpu.dp.rf.reg_file_arr[31][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30405_ (.CLK(_00916_),
    .D(_02140_),
    .Q(\rvcpu.dp.rf.reg_file_arr[31][16] ));
 sky130_fd_sc_hd__dfxtp_1 _30406_ (.CLK(_00917_),
    .D(_02141_),
    .Q(\rvcpu.dp.rf.reg_file_arr[31][17] ));
 sky130_fd_sc_hd__dfxtp_1 _30407_ (.CLK(_00918_),
    .D(_02142_),
    .Q(\rvcpu.dp.rf.reg_file_arr[31][18] ));
 sky130_fd_sc_hd__dfxtp_1 _30408_ (.CLK(_00919_),
    .D(_02143_),
    .Q(\rvcpu.dp.rf.reg_file_arr[31][19] ));
 sky130_fd_sc_hd__dfxtp_1 _30409_ (.CLK(_00920_),
    .D(_02144_),
    .Q(\rvcpu.dp.rf.reg_file_arr[31][20] ));
 sky130_fd_sc_hd__dfxtp_1 _30410_ (.CLK(_00921_),
    .D(_02145_),
    .Q(\rvcpu.dp.rf.reg_file_arr[31][21] ));
 sky130_fd_sc_hd__dfxtp_1 _30411_ (.CLK(_00922_),
    .D(_02146_),
    .Q(\rvcpu.dp.rf.reg_file_arr[31][22] ));
 sky130_fd_sc_hd__dfxtp_1 _30412_ (.CLK(_00923_),
    .D(_02147_),
    .Q(\rvcpu.dp.rf.reg_file_arr[31][23] ));
 sky130_fd_sc_hd__dfxtp_1 _30413_ (.CLK(_00924_),
    .D(_02148_),
    .Q(\rvcpu.dp.rf.reg_file_arr[31][24] ));
 sky130_fd_sc_hd__dfxtp_1 _30414_ (.CLK(_00925_),
    .D(_02149_),
    .Q(\rvcpu.dp.rf.reg_file_arr[31][25] ));
 sky130_fd_sc_hd__dfxtp_1 _30415_ (.CLK(_00926_),
    .D(_02150_),
    .Q(\rvcpu.dp.rf.reg_file_arr[31][26] ));
 sky130_fd_sc_hd__dfxtp_1 _30416_ (.CLK(_00927_),
    .D(_02151_),
    .Q(\rvcpu.dp.rf.reg_file_arr[31][27] ));
 sky130_fd_sc_hd__dfxtp_1 _30417_ (.CLK(_00928_),
    .D(_02152_),
    .Q(\rvcpu.dp.rf.reg_file_arr[31][28] ));
 sky130_fd_sc_hd__dfxtp_1 _30418_ (.CLK(_00929_),
    .D(_02153_),
    .Q(\rvcpu.dp.rf.reg_file_arr[31][29] ));
 sky130_fd_sc_hd__dfxtp_1 _30419_ (.CLK(_00930_),
    .D(_02154_),
    .Q(\rvcpu.dp.rf.reg_file_arr[31][30] ));
 sky130_fd_sc_hd__dfxtp_1 _30420_ (.CLK(_00931_),
    .D(_02155_),
    .Q(\rvcpu.dp.rf.reg_file_arr[31][31] ));
 sky130_fd_sc_hd__dfxtp_1 _30421_ (.CLK(_00932_),
    .D(_02156_),
    .Q(\rvcpu.dp.rf.reg_file_arr[29][0] ));
 sky130_fd_sc_hd__dfxtp_1 _30422_ (.CLK(_00933_),
    .D(_02157_),
    .Q(\rvcpu.dp.rf.reg_file_arr[29][1] ));
 sky130_fd_sc_hd__dfxtp_1 _30423_ (.CLK(_00934_),
    .D(_02158_),
    .Q(\rvcpu.dp.rf.reg_file_arr[29][2] ));
 sky130_fd_sc_hd__dfxtp_1 _30424_ (.CLK(_00935_),
    .D(_02159_),
    .Q(\rvcpu.dp.rf.reg_file_arr[29][3] ));
 sky130_fd_sc_hd__dfxtp_1 _30425_ (.CLK(_00936_),
    .D(_02160_),
    .Q(\rvcpu.dp.rf.reg_file_arr[29][4] ));
 sky130_fd_sc_hd__dfxtp_1 _30426_ (.CLK(_00937_),
    .D(_02161_),
    .Q(\rvcpu.dp.rf.reg_file_arr[29][5] ));
 sky130_fd_sc_hd__dfxtp_1 _30427_ (.CLK(_00938_),
    .D(_02162_),
    .Q(\rvcpu.dp.rf.reg_file_arr[29][6] ));
 sky130_fd_sc_hd__dfxtp_1 _30428_ (.CLK(_00939_),
    .D(_02163_),
    .Q(\rvcpu.dp.rf.reg_file_arr[29][7] ));
 sky130_fd_sc_hd__dfxtp_1 _30429_ (.CLK(_00940_),
    .D(_02164_),
    .Q(\rvcpu.dp.rf.reg_file_arr[29][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30430_ (.CLK(_00941_),
    .D(_02165_),
    .Q(\rvcpu.dp.rf.reg_file_arr[29][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30431_ (.CLK(_00942_),
    .D(_02166_),
    .Q(\rvcpu.dp.rf.reg_file_arr[29][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30432_ (.CLK(_00943_),
    .D(_02167_),
    .Q(\rvcpu.dp.rf.reg_file_arr[29][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30433_ (.CLK(_00944_),
    .D(_02168_),
    .Q(\rvcpu.dp.rf.reg_file_arr[29][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30434_ (.CLK(_00945_),
    .D(_02169_),
    .Q(\rvcpu.dp.rf.reg_file_arr[29][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30435_ (.CLK(_00946_),
    .D(_02170_),
    .Q(\rvcpu.dp.rf.reg_file_arr[29][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30436_ (.CLK(_00947_),
    .D(_02171_),
    .Q(\rvcpu.dp.rf.reg_file_arr[29][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30437_ (.CLK(_00948_),
    .D(_02172_),
    .Q(\rvcpu.dp.rf.reg_file_arr[29][16] ));
 sky130_fd_sc_hd__dfxtp_1 _30438_ (.CLK(_00949_),
    .D(_02173_),
    .Q(\rvcpu.dp.rf.reg_file_arr[29][17] ));
 sky130_fd_sc_hd__dfxtp_1 _30439_ (.CLK(_00950_),
    .D(_02174_),
    .Q(\rvcpu.dp.rf.reg_file_arr[29][18] ));
 sky130_fd_sc_hd__dfxtp_1 _30440_ (.CLK(_00951_),
    .D(_02175_),
    .Q(\rvcpu.dp.rf.reg_file_arr[29][19] ));
 sky130_fd_sc_hd__dfxtp_1 _30441_ (.CLK(_00952_),
    .D(_02176_),
    .Q(\rvcpu.dp.rf.reg_file_arr[29][20] ));
 sky130_fd_sc_hd__dfxtp_1 _30442_ (.CLK(_00953_),
    .D(_02177_),
    .Q(\rvcpu.dp.rf.reg_file_arr[29][21] ));
 sky130_fd_sc_hd__dfxtp_1 _30443_ (.CLK(_00954_),
    .D(_02178_),
    .Q(\rvcpu.dp.rf.reg_file_arr[29][22] ));
 sky130_fd_sc_hd__dfxtp_1 _30444_ (.CLK(_00955_),
    .D(_02179_),
    .Q(\rvcpu.dp.rf.reg_file_arr[29][23] ));
 sky130_fd_sc_hd__dfxtp_1 _30445_ (.CLK(_00956_),
    .D(_02180_),
    .Q(\rvcpu.dp.rf.reg_file_arr[29][24] ));
 sky130_fd_sc_hd__dfxtp_1 _30446_ (.CLK(_00957_),
    .D(_02181_),
    .Q(\rvcpu.dp.rf.reg_file_arr[29][25] ));
 sky130_fd_sc_hd__dfxtp_1 _30447_ (.CLK(_00958_),
    .D(_02182_),
    .Q(\rvcpu.dp.rf.reg_file_arr[29][26] ));
 sky130_fd_sc_hd__dfxtp_1 _30448_ (.CLK(_00959_),
    .D(_02183_),
    .Q(\rvcpu.dp.rf.reg_file_arr[29][27] ));
 sky130_fd_sc_hd__dfxtp_1 _30449_ (.CLK(_00960_),
    .D(_02184_),
    .Q(\rvcpu.dp.rf.reg_file_arr[29][28] ));
 sky130_fd_sc_hd__dfxtp_1 _30450_ (.CLK(_00961_),
    .D(_02185_),
    .Q(\rvcpu.dp.rf.reg_file_arr[29][29] ));
 sky130_fd_sc_hd__dfxtp_1 _30451_ (.CLK(_00962_),
    .D(_02186_),
    .Q(\rvcpu.dp.rf.reg_file_arr[29][30] ));
 sky130_fd_sc_hd__dfxtp_1 _30452_ (.CLK(_00963_),
    .D(_02187_),
    .Q(\rvcpu.dp.rf.reg_file_arr[29][31] ));
 sky130_fd_sc_hd__dfxtp_1 _30453_ (.CLK(_00964_),
    .D(_02188_),
    .Q(\rvcpu.dp.rf.reg_file_arr[19][0] ));
 sky130_fd_sc_hd__dfxtp_1 _30454_ (.CLK(_00965_),
    .D(_02189_),
    .Q(\rvcpu.dp.rf.reg_file_arr[19][1] ));
 sky130_fd_sc_hd__dfxtp_1 _30455_ (.CLK(_00966_),
    .D(_02190_),
    .Q(\rvcpu.dp.rf.reg_file_arr[19][2] ));
 sky130_fd_sc_hd__dfxtp_1 _30456_ (.CLK(_00967_),
    .D(_02191_),
    .Q(\rvcpu.dp.rf.reg_file_arr[19][3] ));
 sky130_fd_sc_hd__dfxtp_1 _30457_ (.CLK(_00968_),
    .D(_02192_),
    .Q(\rvcpu.dp.rf.reg_file_arr[19][4] ));
 sky130_fd_sc_hd__dfxtp_1 _30458_ (.CLK(_00969_),
    .D(_02193_),
    .Q(\rvcpu.dp.rf.reg_file_arr[19][5] ));
 sky130_fd_sc_hd__dfxtp_1 _30459_ (.CLK(_00970_),
    .D(_02194_),
    .Q(\rvcpu.dp.rf.reg_file_arr[19][6] ));
 sky130_fd_sc_hd__dfxtp_1 _30460_ (.CLK(_00971_),
    .D(_02195_),
    .Q(\rvcpu.dp.rf.reg_file_arr[19][7] ));
 sky130_fd_sc_hd__dfxtp_1 _30461_ (.CLK(_00972_),
    .D(_02196_),
    .Q(\rvcpu.dp.rf.reg_file_arr[19][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30462_ (.CLK(_00973_),
    .D(_02197_),
    .Q(\rvcpu.dp.rf.reg_file_arr[19][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30463_ (.CLK(_00974_),
    .D(_02198_),
    .Q(\rvcpu.dp.rf.reg_file_arr[19][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30464_ (.CLK(_00975_),
    .D(_02199_),
    .Q(\rvcpu.dp.rf.reg_file_arr[19][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30465_ (.CLK(_00976_),
    .D(_02200_),
    .Q(\rvcpu.dp.rf.reg_file_arr[19][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30466_ (.CLK(_00977_),
    .D(_02201_),
    .Q(\rvcpu.dp.rf.reg_file_arr[19][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30467_ (.CLK(_00978_),
    .D(_02202_),
    .Q(\rvcpu.dp.rf.reg_file_arr[19][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30468_ (.CLK(_00979_),
    .D(_02203_),
    .Q(\rvcpu.dp.rf.reg_file_arr[19][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30469_ (.CLK(_00980_),
    .D(_02204_),
    .Q(\rvcpu.dp.rf.reg_file_arr[19][16] ));
 sky130_fd_sc_hd__dfxtp_1 _30470_ (.CLK(_00981_),
    .D(_02205_),
    .Q(\rvcpu.dp.rf.reg_file_arr[19][17] ));
 sky130_fd_sc_hd__dfxtp_1 _30471_ (.CLK(_00982_),
    .D(_02206_),
    .Q(\rvcpu.dp.rf.reg_file_arr[19][18] ));
 sky130_fd_sc_hd__dfxtp_1 _30472_ (.CLK(_00983_),
    .D(_02207_),
    .Q(\rvcpu.dp.rf.reg_file_arr[19][19] ));
 sky130_fd_sc_hd__dfxtp_1 _30473_ (.CLK(_00984_),
    .D(_02208_),
    .Q(\rvcpu.dp.rf.reg_file_arr[19][20] ));
 sky130_fd_sc_hd__dfxtp_1 _30474_ (.CLK(_00985_),
    .D(_02209_),
    .Q(\rvcpu.dp.rf.reg_file_arr[19][21] ));
 sky130_fd_sc_hd__dfxtp_1 _30475_ (.CLK(_00986_),
    .D(_02210_),
    .Q(\rvcpu.dp.rf.reg_file_arr[19][22] ));
 sky130_fd_sc_hd__dfxtp_1 _30476_ (.CLK(_00987_),
    .D(_02211_),
    .Q(\rvcpu.dp.rf.reg_file_arr[19][23] ));
 sky130_fd_sc_hd__dfxtp_1 _30477_ (.CLK(_00988_),
    .D(_02212_),
    .Q(\rvcpu.dp.rf.reg_file_arr[19][24] ));
 sky130_fd_sc_hd__dfxtp_1 _30478_ (.CLK(_00989_),
    .D(_02213_),
    .Q(\rvcpu.dp.rf.reg_file_arr[19][25] ));
 sky130_fd_sc_hd__dfxtp_1 _30479_ (.CLK(_00990_),
    .D(_02214_),
    .Q(\rvcpu.dp.rf.reg_file_arr[19][26] ));
 sky130_fd_sc_hd__dfxtp_1 _30480_ (.CLK(_00991_),
    .D(_02215_),
    .Q(\rvcpu.dp.rf.reg_file_arr[19][27] ));
 sky130_fd_sc_hd__dfxtp_1 _30481_ (.CLK(_00992_),
    .D(_02216_),
    .Q(\rvcpu.dp.rf.reg_file_arr[19][28] ));
 sky130_fd_sc_hd__dfxtp_1 _30482_ (.CLK(_00993_),
    .D(_02217_),
    .Q(\rvcpu.dp.rf.reg_file_arr[19][29] ));
 sky130_fd_sc_hd__dfxtp_1 _30483_ (.CLK(_00994_),
    .D(_02218_),
    .Q(\rvcpu.dp.rf.reg_file_arr[19][30] ));
 sky130_fd_sc_hd__dfxtp_1 _30484_ (.CLK(_00995_),
    .D(_02219_),
    .Q(\rvcpu.dp.rf.reg_file_arr[19][31] ));
 sky130_fd_sc_hd__dfxtp_1 _30485_ (.CLK(clk),
    .D(_02220_),
    .Q(\datamem.data_ram[57][24] ));
 sky130_fd_sc_hd__dfxtp_1 _30486_ (.CLK(clk),
    .D(_02221_),
    .Q(\datamem.data_ram[57][25] ));
 sky130_fd_sc_hd__dfxtp_1 _30487_ (.CLK(clk),
    .D(_02222_),
    .Q(\datamem.data_ram[57][26] ));
 sky130_fd_sc_hd__dfxtp_1 _30488_ (.CLK(clk),
    .D(_02223_),
    .Q(\datamem.data_ram[57][27] ));
 sky130_fd_sc_hd__dfxtp_1 _30489_ (.CLK(clk),
    .D(_02224_),
    .Q(\datamem.data_ram[57][28] ));
 sky130_fd_sc_hd__dfxtp_1 _30490_ (.CLK(clk),
    .D(_02225_),
    .Q(\datamem.data_ram[57][29] ));
 sky130_fd_sc_hd__dfxtp_1 _30491_ (.CLK(clk),
    .D(_02226_),
    .Q(\datamem.data_ram[57][30] ));
 sky130_fd_sc_hd__dfxtp_1 _30492_ (.CLK(clk),
    .D(_02227_),
    .Q(\datamem.data_ram[57][31] ));
 sky130_fd_sc_hd__dfxtp_1 _30493_ (.CLK(clk),
    .D(_02228_),
    .Q(\datamem.data_ram[57][16] ));
 sky130_fd_sc_hd__dfxtp_1 _30494_ (.CLK(clk),
    .D(_02229_),
    .Q(\datamem.data_ram[57][17] ));
 sky130_fd_sc_hd__dfxtp_1 _30495_ (.CLK(clk),
    .D(_02230_),
    .Q(\datamem.data_ram[57][18] ));
 sky130_fd_sc_hd__dfxtp_1 _30496_ (.CLK(clk),
    .D(_02231_),
    .Q(\datamem.data_ram[57][19] ));
 sky130_fd_sc_hd__dfxtp_1 _30497_ (.CLK(clk),
    .D(_02232_),
    .Q(\datamem.data_ram[57][20] ));
 sky130_fd_sc_hd__dfxtp_1 _30498_ (.CLK(clk),
    .D(_02233_),
    .Q(\datamem.data_ram[57][21] ));
 sky130_fd_sc_hd__dfxtp_1 _30499_ (.CLK(clk),
    .D(_02234_),
    .Q(\datamem.data_ram[57][22] ));
 sky130_fd_sc_hd__dfxtp_1 _30500_ (.CLK(clk),
    .D(_02235_),
    .Q(\datamem.data_ram[57][23] ));
 sky130_fd_sc_hd__dfxtp_1 _30501_ (.CLK(clk),
    .D(_02236_),
    .Q(\datamem.data_ram[57][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30502_ (.CLK(clk),
    .D(_02237_),
    .Q(\datamem.data_ram[57][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30503_ (.CLK(clk),
    .D(_02238_),
    .Q(\datamem.data_ram[57][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30504_ (.CLK(clk),
    .D(_02239_),
    .Q(\datamem.data_ram[57][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30505_ (.CLK(clk),
    .D(_02240_),
    .Q(\datamem.data_ram[57][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30506_ (.CLK(clk),
    .D(_02241_),
    .Q(\datamem.data_ram[57][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30507_ (.CLK(clk),
    .D(_02242_),
    .Q(\datamem.data_ram[57][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30508_ (.CLK(clk),
    .D(_02243_),
    .Q(\datamem.data_ram[57][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30509_ (.CLK(clk),
    .D(_02244_),
    .Q(\datamem.data_ram[56][24] ));
 sky130_fd_sc_hd__dfxtp_1 _30510_ (.CLK(clk),
    .D(_02245_),
    .Q(\datamem.data_ram[56][25] ));
 sky130_fd_sc_hd__dfxtp_1 _30511_ (.CLK(clk),
    .D(_02246_),
    .Q(\datamem.data_ram[56][26] ));
 sky130_fd_sc_hd__dfxtp_1 _30512_ (.CLK(clk),
    .D(_02247_),
    .Q(\datamem.data_ram[56][27] ));
 sky130_fd_sc_hd__dfxtp_1 _30513_ (.CLK(clk),
    .D(_02248_),
    .Q(\datamem.data_ram[56][28] ));
 sky130_fd_sc_hd__dfxtp_1 _30514_ (.CLK(clk),
    .D(_02249_),
    .Q(\datamem.data_ram[56][29] ));
 sky130_fd_sc_hd__dfxtp_1 _30515_ (.CLK(clk),
    .D(_02250_),
    .Q(\datamem.data_ram[56][30] ));
 sky130_fd_sc_hd__dfxtp_1 _30516_ (.CLK(clk),
    .D(_02251_),
    .Q(\datamem.data_ram[56][31] ));
 sky130_fd_sc_hd__dfxtp_1 _30517_ (.CLK(clk),
    .D(_02252_),
    .Q(\datamem.data_ram[56][16] ));
 sky130_fd_sc_hd__dfxtp_1 _30518_ (.CLK(clk),
    .D(_02253_),
    .Q(\datamem.data_ram[56][17] ));
 sky130_fd_sc_hd__dfxtp_1 _30519_ (.CLK(clk),
    .D(_02254_),
    .Q(\datamem.data_ram[56][18] ));
 sky130_fd_sc_hd__dfxtp_1 _30520_ (.CLK(clk),
    .D(_02255_),
    .Q(\datamem.data_ram[56][19] ));
 sky130_fd_sc_hd__dfxtp_1 _30521_ (.CLK(clk),
    .D(_02256_),
    .Q(\datamem.data_ram[56][20] ));
 sky130_fd_sc_hd__dfxtp_1 _30522_ (.CLK(clk),
    .D(_02257_),
    .Q(\datamem.data_ram[56][21] ));
 sky130_fd_sc_hd__dfxtp_1 _30523_ (.CLK(clk),
    .D(_02258_),
    .Q(\datamem.data_ram[56][22] ));
 sky130_fd_sc_hd__dfxtp_1 _30524_ (.CLK(clk),
    .D(_02259_),
    .Q(\datamem.data_ram[56][23] ));
 sky130_fd_sc_hd__dfxtp_1 _30525_ (.CLK(clk),
    .D(_02260_),
    .Q(\datamem.data_ram[56][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30526_ (.CLK(clk),
    .D(_02261_),
    .Q(\datamem.data_ram[56][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30527_ (.CLK(clk),
    .D(_02262_),
    .Q(\datamem.data_ram[56][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30528_ (.CLK(clk),
    .D(_02263_),
    .Q(\datamem.data_ram[56][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30529_ (.CLK(clk),
    .D(_02264_),
    .Q(\datamem.data_ram[56][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30530_ (.CLK(clk),
    .D(_02265_),
    .Q(\datamem.data_ram[56][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30531_ (.CLK(clk),
    .D(_02266_),
    .Q(\datamem.data_ram[56][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30532_ (.CLK(clk),
    .D(_02267_),
    .Q(\datamem.data_ram[56][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30533_ (.CLK(clk),
    .D(_02268_),
    .Q(\datamem.data_ram[55][24] ));
 sky130_fd_sc_hd__dfxtp_1 _30534_ (.CLK(clk),
    .D(_02269_),
    .Q(\datamem.data_ram[55][25] ));
 sky130_fd_sc_hd__dfxtp_1 _30535_ (.CLK(clk),
    .D(_02270_),
    .Q(\datamem.data_ram[55][26] ));
 sky130_fd_sc_hd__dfxtp_1 _30536_ (.CLK(clk),
    .D(_02271_),
    .Q(\datamem.data_ram[55][27] ));
 sky130_fd_sc_hd__dfxtp_1 _30537_ (.CLK(clk),
    .D(_02272_),
    .Q(\datamem.data_ram[55][28] ));
 sky130_fd_sc_hd__dfxtp_1 _30538_ (.CLK(clk),
    .D(_02273_),
    .Q(\datamem.data_ram[55][29] ));
 sky130_fd_sc_hd__dfxtp_1 _30539_ (.CLK(clk),
    .D(_02274_),
    .Q(\datamem.data_ram[55][30] ));
 sky130_fd_sc_hd__dfxtp_1 _30540_ (.CLK(clk),
    .D(_02275_),
    .Q(\datamem.data_ram[55][31] ));
 sky130_fd_sc_hd__dfxtp_1 _30541_ (.CLK(clk),
    .D(_02276_),
    .Q(\datamem.data_ram[55][16] ));
 sky130_fd_sc_hd__dfxtp_1 _30542_ (.CLK(clk),
    .D(_02277_),
    .Q(\datamem.data_ram[55][17] ));
 sky130_fd_sc_hd__dfxtp_1 _30543_ (.CLK(clk),
    .D(_02278_),
    .Q(\datamem.data_ram[55][18] ));
 sky130_fd_sc_hd__dfxtp_1 _30544_ (.CLK(clk),
    .D(_02279_),
    .Q(\datamem.data_ram[55][19] ));
 sky130_fd_sc_hd__dfxtp_1 _30545_ (.CLK(clk),
    .D(_02280_),
    .Q(\datamem.data_ram[55][20] ));
 sky130_fd_sc_hd__dfxtp_1 _30546_ (.CLK(clk),
    .D(_02281_),
    .Q(\datamem.data_ram[55][21] ));
 sky130_fd_sc_hd__dfxtp_1 _30547_ (.CLK(clk),
    .D(_02282_),
    .Q(\datamem.data_ram[55][22] ));
 sky130_fd_sc_hd__dfxtp_1 _30548_ (.CLK(clk),
    .D(_02283_),
    .Q(\datamem.data_ram[55][23] ));
 sky130_fd_sc_hd__dfxtp_1 _30549_ (.CLK(clk),
    .D(_02284_),
    .Q(\datamem.data_ram[55][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30550_ (.CLK(clk),
    .D(_02285_),
    .Q(\datamem.data_ram[55][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30551_ (.CLK(clk),
    .D(_02286_),
    .Q(\datamem.data_ram[55][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30552_ (.CLK(clk),
    .D(_02287_),
    .Q(\datamem.data_ram[55][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30553_ (.CLK(clk),
    .D(_02288_),
    .Q(\datamem.data_ram[55][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30554_ (.CLK(clk),
    .D(_02289_),
    .Q(\datamem.data_ram[55][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30555_ (.CLK(clk),
    .D(_02290_),
    .Q(\datamem.data_ram[55][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30556_ (.CLK(clk),
    .D(_02291_),
    .Q(\datamem.data_ram[55][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30557_ (.CLK(clk),
    .D(_02292_),
    .Q(\datamem.data_ram[54][24] ));
 sky130_fd_sc_hd__dfxtp_1 _30558_ (.CLK(clk),
    .D(_02293_),
    .Q(\datamem.data_ram[54][25] ));
 sky130_fd_sc_hd__dfxtp_1 _30559_ (.CLK(clk),
    .D(_02294_),
    .Q(\datamem.data_ram[54][26] ));
 sky130_fd_sc_hd__dfxtp_1 _30560_ (.CLK(clk),
    .D(_02295_),
    .Q(\datamem.data_ram[54][27] ));
 sky130_fd_sc_hd__dfxtp_1 _30561_ (.CLK(clk),
    .D(_02296_),
    .Q(\datamem.data_ram[54][28] ));
 sky130_fd_sc_hd__dfxtp_1 _30562_ (.CLK(clk),
    .D(_02297_),
    .Q(\datamem.data_ram[54][29] ));
 sky130_fd_sc_hd__dfxtp_1 _30563_ (.CLK(clk),
    .D(_02298_),
    .Q(\datamem.data_ram[54][30] ));
 sky130_fd_sc_hd__dfxtp_1 _30564_ (.CLK(clk),
    .D(_02299_),
    .Q(\datamem.data_ram[54][31] ));
 sky130_fd_sc_hd__dfxtp_1 _30565_ (.CLK(clk),
    .D(_02300_),
    .Q(\datamem.data_ram[54][16] ));
 sky130_fd_sc_hd__dfxtp_1 _30566_ (.CLK(clk),
    .D(_02301_),
    .Q(\datamem.data_ram[54][17] ));
 sky130_fd_sc_hd__dfxtp_1 _30567_ (.CLK(clk),
    .D(_02302_),
    .Q(\datamem.data_ram[54][18] ));
 sky130_fd_sc_hd__dfxtp_1 _30568_ (.CLK(clk),
    .D(_02303_),
    .Q(\datamem.data_ram[54][19] ));
 sky130_fd_sc_hd__dfxtp_1 _30569_ (.CLK(clk),
    .D(_02304_),
    .Q(\datamem.data_ram[54][20] ));
 sky130_fd_sc_hd__dfxtp_1 _30570_ (.CLK(clk),
    .D(_02305_),
    .Q(\datamem.data_ram[54][21] ));
 sky130_fd_sc_hd__dfxtp_1 _30571_ (.CLK(clk),
    .D(_02306_),
    .Q(\datamem.data_ram[54][22] ));
 sky130_fd_sc_hd__dfxtp_1 _30572_ (.CLK(clk),
    .D(_02307_),
    .Q(\datamem.data_ram[54][23] ));
 sky130_fd_sc_hd__dfxtp_1 _30573_ (.CLK(clk),
    .D(_02308_),
    .Q(\datamem.data_ram[54][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30574_ (.CLK(clk),
    .D(_02309_),
    .Q(\datamem.data_ram[54][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30575_ (.CLK(clk),
    .D(_02310_),
    .Q(\datamem.data_ram[54][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30576_ (.CLK(clk),
    .D(_02311_),
    .Q(\datamem.data_ram[54][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30577_ (.CLK(clk),
    .D(_02312_),
    .Q(\datamem.data_ram[54][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30578_ (.CLK(clk),
    .D(_02313_),
    .Q(\datamem.data_ram[54][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30579_ (.CLK(clk),
    .D(_02314_),
    .Q(\datamem.data_ram[54][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30580_ (.CLK(clk),
    .D(_02315_),
    .Q(\datamem.data_ram[54][15] ));
 sky130_fd_sc_hd__dfxtp_2 _30581_ (.CLK(clk),
    .D(_02316_),
    .Q(\datamem.data_ram[53][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30582_ (.CLK(clk),
    .D(_02317_),
    .Q(\datamem.data_ram[53][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30583_ (.CLK(clk),
    .D(_02318_),
    .Q(\datamem.data_ram[53][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30584_ (.CLK(clk),
    .D(_02319_),
    .Q(\datamem.data_ram[53][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30585_ (.CLK(clk),
    .D(_02320_),
    .Q(\datamem.data_ram[53][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30586_ (.CLK(clk),
    .D(_02321_),
    .Q(\datamem.data_ram[53][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30587_ (.CLK(clk),
    .D(_02322_),
    .Q(\datamem.data_ram[53][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30588_ (.CLK(clk),
    .D(_02323_),
    .Q(\datamem.data_ram[53][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30589_ (.CLK(clk),
    .D(_02324_),
    .Q(\datamem.data_ram[53][0] ));
 sky130_fd_sc_hd__dfxtp_1 _30590_ (.CLK(clk),
    .D(_02325_),
    .Q(\datamem.data_ram[53][1] ));
 sky130_fd_sc_hd__dfxtp_1 _30591_ (.CLK(clk),
    .D(_02326_),
    .Q(\datamem.data_ram[53][2] ));
 sky130_fd_sc_hd__dfxtp_2 _30592_ (.CLK(clk),
    .D(_02327_),
    .Q(\datamem.data_ram[53][3] ));
 sky130_fd_sc_hd__dfxtp_1 _30593_ (.CLK(clk),
    .D(_02328_),
    .Q(\datamem.data_ram[53][4] ));
 sky130_fd_sc_hd__dfxtp_1 _30594_ (.CLK(clk),
    .D(_02329_),
    .Q(\datamem.data_ram[53][5] ));
 sky130_fd_sc_hd__dfxtp_1 _30595_ (.CLK(clk),
    .D(_02330_),
    .Q(\datamem.data_ram[53][6] ));
 sky130_fd_sc_hd__dfxtp_2 _30596_ (.CLK(clk),
    .D(_02331_),
    .Q(\datamem.data_ram[53][7] ));
 sky130_fd_sc_hd__dfxtp_1 _30597_ (.CLK(clk),
    .D(_02332_),
    .Q(\datamem.data_ram[53][24] ));
 sky130_fd_sc_hd__dfxtp_1 _30598_ (.CLK(clk),
    .D(_02333_),
    .Q(\datamem.data_ram[53][25] ));
 sky130_fd_sc_hd__dfxtp_1 _30599_ (.CLK(clk),
    .D(_02334_),
    .Q(\datamem.data_ram[53][26] ));
 sky130_fd_sc_hd__dfxtp_1 _30600_ (.CLK(clk),
    .D(_02335_),
    .Q(\datamem.data_ram[53][27] ));
 sky130_fd_sc_hd__dfxtp_1 _30601_ (.CLK(clk),
    .D(_02336_),
    .Q(\datamem.data_ram[53][28] ));
 sky130_fd_sc_hd__dfxtp_1 _30602_ (.CLK(clk),
    .D(_02337_),
    .Q(\datamem.data_ram[53][29] ));
 sky130_fd_sc_hd__dfxtp_1 _30603_ (.CLK(clk),
    .D(_02338_),
    .Q(\datamem.data_ram[53][30] ));
 sky130_fd_sc_hd__dfxtp_1 _30604_ (.CLK(clk),
    .D(_02339_),
    .Q(\datamem.data_ram[53][31] ));
 sky130_fd_sc_hd__dfxtp_1 _30605_ (.CLK(clk),
    .D(_02340_),
    .Q(\datamem.data_ram[52][24] ));
 sky130_fd_sc_hd__dfxtp_1 _30606_ (.CLK(clk),
    .D(_02341_),
    .Q(\datamem.data_ram[52][25] ));
 sky130_fd_sc_hd__dfxtp_1 _30607_ (.CLK(clk),
    .D(_02342_),
    .Q(\datamem.data_ram[52][26] ));
 sky130_fd_sc_hd__dfxtp_1 _30608_ (.CLK(clk),
    .D(_02343_),
    .Q(\datamem.data_ram[52][27] ));
 sky130_fd_sc_hd__dfxtp_2 _30609_ (.CLK(clk),
    .D(_02344_),
    .Q(\datamem.data_ram[52][28] ));
 sky130_fd_sc_hd__dfxtp_1 _30610_ (.CLK(clk),
    .D(_02345_),
    .Q(\datamem.data_ram[52][29] ));
 sky130_fd_sc_hd__dfxtp_1 _30611_ (.CLK(clk),
    .D(_02346_),
    .Q(\datamem.data_ram[52][30] ));
 sky130_fd_sc_hd__dfxtp_1 _30612_ (.CLK(clk),
    .D(_02347_),
    .Q(\datamem.data_ram[52][31] ));
 sky130_fd_sc_hd__dfxtp_1 _30613_ (.CLK(clk),
    .D(_02348_),
    .Q(\datamem.data_ram[52][16] ));
 sky130_fd_sc_hd__dfxtp_1 _30614_ (.CLK(clk),
    .D(_02349_),
    .Q(\datamem.data_ram[52][17] ));
 sky130_fd_sc_hd__dfxtp_1 _30615_ (.CLK(clk),
    .D(_02350_),
    .Q(\datamem.data_ram[52][18] ));
 sky130_fd_sc_hd__dfxtp_1 _30616_ (.CLK(clk),
    .D(_02351_),
    .Q(\datamem.data_ram[52][19] ));
 sky130_fd_sc_hd__dfxtp_1 _30617_ (.CLK(clk),
    .D(_02352_),
    .Q(\datamem.data_ram[52][20] ));
 sky130_fd_sc_hd__dfxtp_1 _30618_ (.CLK(clk),
    .D(_02353_),
    .Q(\datamem.data_ram[52][21] ));
 sky130_fd_sc_hd__dfxtp_1 _30619_ (.CLK(clk),
    .D(_02354_),
    .Q(\datamem.data_ram[52][22] ));
 sky130_fd_sc_hd__dfxtp_1 _30620_ (.CLK(clk),
    .D(_02355_),
    .Q(\datamem.data_ram[52][23] ));
 sky130_fd_sc_hd__dfxtp_2 _30621_ (.CLK(clk),
    .D(_02356_),
    .Q(\datamem.data_ram[52][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30622_ (.CLK(clk),
    .D(_02357_),
    .Q(\datamem.data_ram[52][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30623_ (.CLK(clk),
    .D(_02358_),
    .Q(\datamem.data_ram[52][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30624_ (.CLK(clk),
    .D(_02359_),
    .Q(\datamem.data_ram[52][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30625_ (.CLK(clk),
    .D(_02360_),
    .Q(\datamem.data_ram[52][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30626_ (.CLK(clk),
    .D(_02361_),
    .Q(\datamem.data_ram[52][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30627_ (.CLK(clk),
    .D(_02362_),
    .Q(\datamem.data_ram[52][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30628_ (.CLK(clk),
    .D(_02363_),
    .Q(\datamem.data_ram[52][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30629_ (.CLK(clk),
    .D(_02364_),
    .Q(\datamem.data_ram[51][24] ));
 sky130_fd_sc_hd__dfxtp_1 _30630_ (.CLK(clk),
    .D(_02365_),
    .Q(\datamem.data_ram[51][25] ));
 sky130_fd_sc_hd__dfxtp_1 _30631_ (.CLK(clk),
    .D(_02366_),
    .Q(\datamem.data_ram[51][26] ));
 sky130_fd_sc_hd__dfxtp_1 _30632_ (.CLK(clk),
    .D(_02367_),
    .Q(\datamem.data_ram[51][27] ));
 sky130_fd_sc_hd__dfxtp_1 _30633_ (.CLK(clk),
    .D(_02368_),
    .Q(\datamem.data_ram[51][28] ));
 sky130_fd_sc_hd__dfxtp_1 _30634_ (.CLK(clk),
    .D(_02369_),
    .Q(\datamem.data_ram[51][29] ));
 sky130_fd_sc_hd__dfxtp_1 _30635_ (.CLK(clk),
    .D(_02370_),
    .Q(\datamem.data_ram[51][30] ));
 sky130_fd_sc_hd__dfxtp_1 _30636_ (.CLK(clk),
    .D(_02371_),
    .Q(\datamem.data_ram[51][31] ));
 sky130_fd_sc_hd__dfxtp_1 _30637_ (.CLK(clk),
    .D(_02372_),
    .Q(\datamem.data_ram[51][16] ));
 sky130_fd_sc_hd__dfxtp_1 _30638_ (.CLK(clk),
    .D(_02373_),
    .Q(\datamem.data_ram[51][17] ));
 sky130_fd_sc_hd__dfxtp_1 _30639_ (.CLK(clk),
    .D(_02374_),
    .Q(\datamem.data_ram[51][18] ));
 sky130_fd_sc_hd__dfxtp_1 _30640_ (.CLK(clk),
    .D(_02375_),
    .Q(\datamem.data_ram[51][19] ));
 sky130_fd_sc_hd__dfxtp_1 _30641_ (.CLK(clk),
    .D(_02376_),
    .Q(\datamem.data_ram[51][20] ));
 sky130_fd_sc_hd__dfxtp_1 _30642_ (.CLK(clk),
    .D(_02377_),
    .Q(\datamem.data_ram[51][21] ));
 sky130_fd_sc_hd__dfxtp_1 _30643_ (.CLK(clk),
    .D(_02378_),
    .Q(\datamem.data_ram[51][22] ));
 sky130_fd_sc_hd__dfxtp_1 _30644_ (.CLK(clk),
    .D(_02379_),
    .Q(\datamem.data_ram[51][23] ));
 sky130_fd_sc_hd__dfxtp_1 _30645_ (.CLK(clk),
    .D(_02380_),
    .Q(\datamem.data_ram[51][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30646_ (.CLK(clk),
    .D(_02381_),
    .Q(\datamem.data_ram[51][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30647_ (.CLK(clk),
    .D(_02382_),
    .Q(\datamem.data_ram[51][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30648_ (.CLK(clk),
    .D(_02383_),
    .Q(\datamem.data_ram[51][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30649_ (.CLK(clk),
    .D(_02384_),
    .Q(\datamem.data_ram[51][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30650_ (.CLK(clk),
    .D(_02385_),
    .Q(\datamem.data_ram[51][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30651_ (.CLK(clk),
    .D(_02386_),
    .Q(\datamem.data_ram[51][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30652_ (.CLK(clk),
    .D(_02387_),
    .Q(\datamem.data_ram[51][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30653_ (.CLK(clk),
    .D(_02388_),
    .Q(\datamem.data_ram[50][24] ));
 sky130_fd_sc_hd__dfxtp_1 _30654_ (.CLK(clk),
    .D(_02389_),
    .Q(\datamem.data_ram[50][25] ));
 sky130_fd_sc_hd__dfxtp_1 _30655_ (.CLK(clk),
    .D(_02390_),
    .Q(\datamem.data_ram[50][26] ));
 sky130_fd_sc_hd__dfxtp_1 _30656_ (.CLK(clk),
    .D(_02391_),
    .Q(\datamem.data_ram[50][27] ));
 sky130_fd_sc_hd__dfxtp_1 _30657_ (.CLK(clk),
    .D(_02392_),
    .Q(\datamem.data_ram[50][28] ));
 sky130_fd_sc_hd__dfxtp_1 _30658_ (.CLK(clk),
    .D(_02393_),
    .Q(\datamem.data_ram[50][29] ));
 sky130_fd_sc_hd__dfxtp_1 _30659_ (.CLK(clk),
    .D(_02394_),
    .Q(\datamem.data_ram[50][30] ));
 sky130_fd_sc_hd__dfxtp_1 _30660_ (.CLK(clk),
    .D(_02395_),
    .Q(\datamem.data_ram[50][31] ));
 sky130_fd_sc_hd__dfxtp_1 _30661_ (.CLK(clk),
    .D(_02396_),
    .Q(\datamem.data_ram[50][16] ));
 sky130_fd_sc_hd__dfxtp_1 _30662_ (.CLK(clk),
    .D(_02397_),
    .Q(\datamem.data_ram[50][17] ));
 sky130_fd_sc_hd__dfxtp_1 _30663_ (.CLK(clk),
    .D(_02398_),
    .Q(\datamem.data_ram[50][18] ));
 sky130_fd_sc_hd__dfxtp_1 _30664_ (.CLK(clk),
    .D(_02399_),
    .Q(\datamem.data_ram[50][19] ));
 sky130_fd_sc_hd__dfxtp_1 _30665_ (.CLK(clk),
    .D(_02400_),
    .Q(\datamem.data_ram[50][20] ));
 sky130_fd_sc_hd__dfxtp_1 _30666_ (.CLK(clk),
    .D(_02401_),
    .Q(\datamem.data_ram[50][21] ));
 sky130_fd_sc_hd__dfxtp_1 _30667_ (.CLK(clk),
    .D(_02402_),
    .Q(\datamem.data_ram[50][22] ));
 sky130_fd_sc_hd__dfxtp_1 _30668_ (.CLK(clk),
    .D(_02403_),
    .Q(\datamem.data_ram[50][23] ));
 sky130_fd_sc_hd__dfxtp_1 _30669_ (.CLK(clk),
    .D(_02404_),
    .Q(\datamem.data_ram[50][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30670_ (.CLK(clk),
    .D(_02405_),
    .Q(\datamem.data_ram[50][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30671_ (.CLK(clk),
    .D(_02406_),
    .Q(\datamem.data_ram[50][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30672_ (.CLK(clk),
    .D(_02407_),
    .Q(\datamem.data_ram[50][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30673_ (.CLK(clk),
    .D(_02408_),
    .Q(\datamem.data_ram[50][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30674_ (.CLK(clk),
    .D(_02409_),
    .Q(\datamem.data_ram[50][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30675_ (.CLK(clk),
    .D(_02410_),
    .Q(\datamem.data_ram[50][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30676_ (.CLK(clk),
    .D(_02411_),
    .Q(\datamem.data_ram[50][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30677_ (.CLK(clk),
    .D(_02412_),
    .Q(\datamem.data_ram[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _30678_ (.CLK(clk),
    .D(_02413_),
    .Q(\datamem.data_ram[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _30679_ (.CLK(clk),
    .D(_02414_),
    .Q(\datamem.data_ram[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _30680_ (.CLK(clk),
    .D(_02415_),
    .Q(\datamem.data_ram[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _30681_ (.CLK(clk),
    .D(_02416_),
    .Q(\datamem.data_ram[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _30682_ (.CLK(clk),
    .D(_02417_),
    .Q(\datamem.data_ram[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _30683_ (.CLK(clk),
    .D(_02418_),
    .Q(\datamem.data_ram[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _30684_ (.CLK(clk),
    .D(_02419_),
    .Q(\datamem.data_ram[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _30685_ (.CLK(clk),
    .D(_02420_),
    .Q(\datamem.data_ram[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30686_ (.CLK(clk),
    .D(_02421_),
    .Q(\datamem.data_ram[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30687_ (.CLK(clk),
    .D(_02422_),
    .Q(\datamem.data_ram[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30688_ (.CLK(clk),
    .D(_02423_),
    .Q(\datamem.data_ram[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30689_ (.CLK(clk),
    .D(_02424_),
    .Q(\datamem.data_ram[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30690_ (.CLK(clk),
    .D(_02425_),
    .Q(\datamem.data_ram[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30691_ (.CLK(clk),
    .D(_02426_),
    .Q(\datamem.data_ram[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30692_ (.CLK(clk),
    .D(_02427_),
    .Q(\datamem.data_ram[4][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30693_ (.CLK(clk),
    .D(_02428_),
    .Q(\datamem.data_ram[4][16] ));
 sky130_fd_sc_hd__dfxtp_1 _30694_ (.CLK(clk),
    .D(_02429_),
    .Q(\datamem.data_ram[4][17] ));
 sky130_fd_sc_hd__dfxtp_1 _30695_ (.CLK(clk),
    .D(_02430_),
    .Q(\datamem.data_ram[4][18] ));
 sky130_fd_sc_hd__dfxtp_1 _30696_ (.CLK(clk),
    .D(_02431_),
    .Q(\datamem.data_ram[4][19] ));
 sky130_fd_sc_hd__dfxtp_1 _30697_ (.CLK(clk),
    .D(_02432_),
    .Q(\datamem.data_ram[4][20] ));
 sky130_fd_sc_hd__dfxtp_1 _30698_ (.CLK(clk),
    .D(_02433_),
    .Q(\datamem.data_ram[4][21] ));
 sky130_fd_sc_hd__dfxtp_1 _30699_ (.CLK(clk),
    .D(_02434_),
    .Q(\datamem.data_ram[4][22] ));
 sky130_fd_sc_hd__dfxtp_1 _30700_ (.CLK(clk),
    .D(_02435_),
    .Q(\datamem.data_ram[4][23] ));
 sky130_fd_sc_hd__dfxtp_1 _30701_ (.CLK(clk),
    .D(_02436_),
    .Q(\datamem.data_ram[49][24] ));
 sky130_fd_sc_hd__dfxtp_1 _30702_ (.CLK(clk),
    .D(_02437_),
    .Q(\datamem.data_ram[49][25] ));
 sky130_fd_sc_hd__dfxtp_1 _30703_ (.CLK(clk),
    .D(_02438_),
    .Q(\datamem.data_ram[49][26] ));
 sky130_fd_sc_hd__dfxtp_1 _30704_ (.CLK(clk),
    .D(_02439_),
    .Q(\datamem.data_ram[49][27] ));
 sky130_fd_sc_hd__dfxtp_1 _30705_ (.CLK(clk),
    .D(_02440_),
    .Q(\datamem.data_ram[49][28] ));
 sky130_fd_sc_hd__dfxtp_1 _30706_ (.CLK(clk),
    .D(_02441_),
    .Q(\datamem.data_ram[49][29] ));
 sky130_fd_sc_hd__dfxtp_1 _30707_ (.CLK(clk),
    .D(_02442_),
    .Q(\datamem.data_ram[49][30] ));
 sky130_fd_sc_hd__dfxtp_1 _30708_ (.CLK(clk),
    .D(_02443_),
    .Q(\datamem.data_ram[49][31] ));
 sky130_fd_sc_hd__dfxtp_1 _30709_ (.CLK(clk),
    .D(_02444_),
    .Q(\datamem.data_ram[49][16] ));
 sky130_fd_sc_hd__dfxtp_1 _30710_ (.CLK(clk),
    .D(_02445_),
    .Q(\datamem.data_ram[49][17] ));
 sky130_fd_sc_hd__dfxtp_1 _30711_ (.CLK(clk),
    .D(_02446_),
    .Q(\datamem.data_ram[49][18] ));
 sky130_fd_sc_hd__dfxtp_1 _30712_ (.CLK(clk),
    .D(_02447_),
    .Q(\datamem.data_ram[49][19] ));
 sky130_fd_sc_hd__dfxtp_1 _30713_ (.CLK(clk),
    .D(_02448_),
    .Q(\datamem.data_ram[49][20] ));
 sky130_fd_sc_hd__dfxtp_1 _30714_ (.CLK(clk),
    .D(_02449_),
    .Q(\datamem.data_ram[49][21] ));
 sky130_fd_sc_hd__dfxtp_1 _30715_ (.CLK(clk),
    .D(_02450_),
    .Q(\datamem.data_ram[49][22] ));
 sky130_fd_sc_hd__dfxtp_1 _30716_ (.CLK(clk),
    .D(_02451_),
    .Q(\datamem.data_ram[49][23] ));
 sky130_fd_sc_hd__dfxtp_1 _30717_ (.CLK(clk),
    .D(_02452_),
    .Q(\datamem.data_ram[49][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30718_ (.CLK(clk),
    .D(_02453_),
    .Q(\datamem.data_ram[49][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30719_ (.CLK(clk),
    .D(_02454_),
    .Q(\datamem.data_ram[49][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30720_ (.CLK(clk),
    .D(_02455_),
    .Q(\datamem.data_ram[49][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30721_ (.CLK(clk),
    .D(_02456_),
    .Q(\datamem.data_ram[49][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30722_ (.CLK(clk),
    .D(_02457_),
    .Q(\datamem.data_ram[49][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30723_ (.CLK(clk),
    .D(_02458_),
    .Q(\datamem.data_ram[49][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30724_ (.CLK(clk),
    .D(_02459_),
    .Q(\datamem.data_ram[49][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30725_ (.CLK(clk),
    .D(_02460_),
    .Q(\datamem.data_ram[48][24] ));
 sky130_fd_sc_hd__dfxtp_1 _30726_ (.CLK(clk),
    .D(_02461_),
    .Q(\datamem.data_ram[48][25] ));
 sky130_fd_sc_hd__dfxtp_1 _30727_ (.CLK(clk),
    .D(_02462_),
    .Q(\datamem.data_ram[48][26] ));
 sky130_fd_sc_hd__dfxtp_1 _30728_ (.CLK(clk),
    .D(_02463_),
    .Q(\datamem.data_ram[48][27] ));
 sky130_fd_sc_hd__dfxtp_1 _30729_ (.CLK(clk),
    .D(_02464_),
    .Q(\datamem.data_ram[48][28] ));
 sky130_fd_sc_hd__dfxtp_1 _30730_ (.CLK(clk),
    .D(_02465_),
    .Q(\datamem.data_ram[48][29] ));
 sky130_fd_sc_hd__dfxtp_1 _30731_ (.CLK(clk),
    .D(_02466_),
    .Q(\datamem.data_ram[48][30] ));
 sky130_fd_sc_hd__dfxtp_1 _30732_ (.CLK(clk),
    .D(_02467_),
    .Q(\datamem.data_ram[48][31] ));
 sky130_fd_sc_hd__dfxtp_1 _30733_ (.CLK(clk),
    .D(_02468_),
    .Q(\datamem.data_ram[47][24] ));
 sky130_fd_sc_hd__dfxtp_1 _30734_ (.CLK(clk),
    .D(_02469_),
    .Q(\datamem.data_ram[47][25] ));
 sky130_fd_sc_hd__dfxtp_1 _30735_ (.CLK(clk),
    .D(_02470_),
    .Q(\datamem.data_ram[47][26] ));
 sky130_fd_sc_hd__dfxtp_1 _30736_ (.CLK(clk),
    .D(_02471_),
    .Q(\datamem.data_ram[47][27] ));
 sky130_fd_sc_hd__dfxtp_1 _30737_ (.CLK(clk),
    .D(_02472_),
    .Q(\datamem.data_ram[47][28] ));
 sky130_fd_sc_hd__dfxtp_1 _30738_ (.CLK(clk),
    .D(_02473_),
    .Q(\datamem.data_ram[47][29] ));
 sky130_fd_sc_hd__dfxtp_1 _30739_ (.CLK(clk),
    .D(_02474_),
    .Q(\datamem.data_ram[47][30] ));
 sky130_fd_sc_hd__dfxtp_1 _30740_ (.CLK(clk),
    .D(_02475_),
    .Q(\datamem.data_ram[47][31] ));
 sky130_fd_sc_hd__dfxtp_1 _30741_ (.CLK(clk),
    .D(_02476_),
    .Q(\datamem.data_ram[48][16] ));
 sky130_fd_sc_hd__dfxtp_1 _30742_ (.CLK(clk),
    .D(_02477_),
    .Q(\datamem.data_ram[48][17] ));
 sky130_fd_sc_hd__dfxtp_1 _30743_ (.CLK(clk),
    .D(_02478_),
    .Q(\datamem.data_ram[48][18] ));
 sky130_fd_sc_hd__dfxtp_1 _30744_ (.CLK(clk),
    .D(_02479_),
    .Q(\datamem.data_ram[48][19] ));
 sky130_fd_sc_hd__dfxtp_1 _30745_ (.CLK(clk),
    .D(_02480_),
    .Q(\datamem.data_ram[48][20] ));
 sky130_fd_sc_hd__dfxtp_1 _30746_ (.CLK(clk),
    .D(_02481_),
    .Q(\datamem.data_ram[48][21] ));
 sky130_fd_sc_hd__dfxtp_1 _30747_ (.CLK(clk),
    .D(_02482_),
    .Q(\datamem.data_ram[48][22] ));
 sky130_fd_sc_hd__dfxtp_1 _30748_ (.CLK(clk),
    .D(_02483_),
    .Q(\datamem.data_ram[48][23] ));
 sky130_fd_sc_hd__dfxtp_1 _30749_ (.CLK(clk),
    .D(_02484_),
    .Q(\datamem.data_ram[48][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30750_ (.CLK(clk),
    .D(_02485_),
    .Q(\datamem.data_ram[48][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30751_ (.CLK(clk),
    .D(_02486_),
    .Q(\datamem.data_ram[48][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30752_ (.CLK(clk),
    .D(_02487_),
    .Q(\datamem.data_ram[48][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30753_ (.CLK(clk),
    .D(_02488_),
    .Q(\datamem.data_ram[48][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30754_ (.CLK(clk),
    .D(_02489_),
    .Q(\datamem.data_ram[48][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30755_ (.CLK(clk),
    .D(_02490_),
    .Q(\datamem.data_ram[48][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30756_ (.CLK(clk),
    .D(_02491_),
    .Q(\datamem.data_ram[48][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30757_ (.CLK(clk),
    .D(_02492_),
    .Q(\datamem.data_ram[47][16] ));
 sky130_fd_sc_hd__dfxtp_1 _30758_ (.CLK(clk),
    .D(_02493_),
    .Q(\datamem.data_ram[47][17] ));
 sky130_fd_sc_hd__dfxtp_1 _30759_ (.CLK(clk),
    .D(_02494_),
    .Q(\datamem.data_ram[47][18] ));
 sky130_fd_sc_hd__dfxtp_1 _30760_ (.CLK(clk),
    .D(_02495_),
    .Q(\datamem.data_ram[47][19] ));
 sky130_fd_sc_hd__dfxtp_1 _30761_ (.CLK(clk),
    .D(_02496_),
    .Q(\datamem.data_ram[47][20] ));
 sky130_fd_sc_hd__dfxtp_1 _30762_ (.CLK(clk),
    .D(_02497_),
    .Q(\datamem.data_ram[47][21] ));
 sky130_fd_sc_hd__dfxtp_1 _30763_ (.CLK(clk),
    .D(_02498_),
    .Q(\datamem.data_ram[47][22] ));
 sky130_fd_sc_hd__dfxtp_1 _30764_ (.CLK(clk),
    .D(_02499_),
    .Q(\datamem.data_ram[47][23] ));
 sky130_fd_sc_hd__dfxtp_1 _30765_ (.CLK(clk),
    .D(_02500_),
    .Q(\datamem.data_ram[47][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30766_ (.CLK(clk),
    .D(_02501_),
    .Q(\datamem.data_ram[47][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30767_ (.CLK(clk),
    .D(_02502_),
    .Q(\datamem.data_ram[47][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30768_ (.CLK(clk),
    .D(_02503_),
    .Q(\datamem.data_ram[47][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30769_ (.CLK(clk),
    .D(_02504_),
    .Q(\datamem.data_ram[47][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30770_ (.CLK(clk),
    .D(_02505_),
    .Q(\datamem.data_ram[47][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30771_ (.CLK(clk),
    .D(_02506_),
    .Q(\datamem.data_ram[47][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30772_ (.CLK(clk),
    .D(_02507_),
    .Q(\datamem.data_ram[47][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30773_ (.CLK(clk),
    .D(_02508_),
    .Q(\datamem.data_ram[46][24] ));
 sky130_fd_sc_hd__dfxtp_1 _30774_ (.CLK(clk),
    .D(_02509_),
    .Q(\datamem.data_ram[46][25] ));
 sky130_fd_sc_hd__dfxtp_1 _30775_ (.CLK(clk),
    .D(_02510_),
    .Q(\datamem.data_ram[46][26] ));
 sky130_fd_sc_hd__dfxtp_1 _30776_ (.CLK(clk),
    .D(_02511_),
    .Q(\datamem.data_ram[46][27] ));
 sky130_fd_sc_hd__dfxtp_1 _30777_ (.CLK(clk),
    .D(_02512_),
    .Q(\datamem.data_ram[46][28] ));
 sky130_fd_sc_hd__dfxtp_1 _30778_ (.CLK(clk),
    .D(_02513_),
    .Q(\datamem.data_ram[46][29] ));
 sky130_fd_sc_hd__dfxtp_1 _30779_ (.CLK(clk),
    .D(_02514_),
    .Q(\datamem.data_ram[46][30] ));
 sky130_fd_sc_hd__dfxtp_1 _30780_ (.CLK(clk),
    .D(_02515_),
    .Q(\datamem.data_ram[46][31] ));
 sky130_fd_sc_hd__dfxtp_1 _30781_ (.CLK(clk),
    .D(_02516_),
    .Q(\datamem.data_ram[46][16] ));
 sky130_fd_sc_hd__dfxtp_1 _30782_ (.CLK(clk),
    .D(_02517_),
    .Q(\datamem.data_ram[46][17] ));
 sky130_fd_sc_hd__dfxtp_1 _30783_ (.CLK(clk),
    .D(_02518_),
    .Q(\datamem.data_ram[46][18] ));
 sky130_fd_sc_hd__dfxtp_1 _30784_ (.CLK(clk),
    .D(_02519_),
    .Q(\datamem.data_ram[46][19] ));
 sky130_fd_sc_hd__dfxtp_1 _30785_ (.CLK(clk),
    .D(_02520_),
    .Q(\datamem.data_ram[46][20] ));
 sky130_fd_sc_hd__dfxtp_1 _30786_ (.CLK(clk),
    .D(_02521_),
    .Q(\datamem.data_ram[46][21] ));
 sky130_fd_sc_hd__dfxtp_1 _30787_ (.CLK(clk),
    .D(_02522_),
    .Q(\datamem.data_ram[46][22] ));
 sky130_fd_sc_hd__dfxtp_1 _30788_ (.CLK(clk),
    .D(_02523_),
    .Q(\datamem.data_ram[46][23] ));
 sky130_fd_sc_hd__dfxtp_1 _30789_ (.CLK(clk),
    .D(_02524_),
    .Q(\datamem.data_ram[46][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30790_ (.CLK(clk),
    .D(_02525_),
    .Q(\datamem.data_ram[46][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30791_ (.CLK(clk),
    .D(_02526_),
    .Q(\datamem.data_ram[46][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30792_ (.CLK(clk),
    .D(_02527_),
    .Q(\datamem.data_ram[46][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30793_ (.CLK(clk),
    .D(_02528_),
    .Q(\datamem.data_ram[46][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30794_ (.CLK(clk),
    .D(_02529_),
    .Q(\datamem.data_ram[46][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30795_ (.CLK(clk),
    .D(_02530_),
    .Q(\datamem.data_ram[46][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30796_ (.CLK(clk),
    .D(_02531_),
    .Q(\datamem.data_ram[46][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30797_ (.CLK(clk),
    .D(_02532_),
    .Q(\datamem.data_ram[45][24] ));
 sky130_fd_sc_hd__dfxtp_1 _30798_ (.CLK(clk),
    .D(_02533_),
    .Q(\datamem.data_ram[45][25] ));
 sky130_fd_sc_hd__dfxtp_1 _30799_ (.CLK(clk),
    .D(_02534_),
    .Q(\datamem.data_ram[45][26] ));
 sky130_fd_sc_hd__dfxtp_1 _30800_ (.CLK(clk),
    .D(_02535_),
    .Q(\datamem.data_ram[45][27] ));
 sky130_fd_sc_hd__dfxtp_1 _30801_ (.CLK(clk),
    .D(_02536_),
    .Q(\datamem.data_ram[45][28] ));
 sky130_fd_sc_hd__dfxtp_1 _30802_ (.CLK(clk),
    .D(_02537_),
    .Q(\datamem.data_ram[45][29] ));
 sky130_fd_sc_hd__dfxtp_1 _30803_ (.CLK(clk),
    .D(_02538_),
    .Q(\datamem.data_ram[45][30] ));
 sky130_fd_sc_hd__dfxtp_1 _30804_ (.CLK(clk),
    .D(_02539_),
    .Q(\datamem.data_ram[45][31] ));
 sky130_fd_sc_hd__dfxtp_1 _30805_ (.CLK(clk),
    .D(_02540_),
    .Q(\datamem.data_ram[45][16] ));
 sky130_fd_sc_hd__dfxtp_1 _30806_ (.CLK(clk),
    .D(_02541_),
    .Q(\datamem.data_ram[45][17] ));
 sky130_fd_sc_hd__dfxtp_1 _30807_ (.CLK(clk),
    .D(_02542_),
    .Q(\datamem.data_ram[45][18] ));
 sky130_fd_sc_hd__dfxtp_1 _30808_ (.CLK(clk),
    .D(_02543_),
    .Q(\datamem.data_ram[45][19] ));
 sky130_fd_sc_hd__dfxtp_1 _30809_ (.CLK(clk),
    .D(_02544_),
    .Q(\datamem.data_ram[45][20] ));
 sky130_fd_sc_hd__dfxtp_1 _30810_ (.CLK(clk),
    .D(_02545_),
    .Q(\datamem.data_ram[45][21] ));
 sky130_fd_sc_hd__dfxtp_1 _30811_ (.CLK(clk),
    .D(_02546_),
    .Q(\datamem.data_ram[45][22] ));
 sky130_fd_sc_hd__dfxtp_1 _30812_ (.CLK(clk),
    .D(_02547_),
    .Q(\datamem.data_ram[45][23] ));
 sky130_fd_sc_hd__dfxtp_1 _30813_ (.CLK(clk),
    .D(_02548_),
    .Q(\datamem.data_ram[45][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30814_ (.CLK(clk),
    .D(_02549_),
    .Q(\datamem.data_ram[45][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30815_ (.CLK(clk),
    .D(_02550_),
    .Q(\datamem.data_ram[45][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30816_ (.CLK(clk),
    .D(_02551_),
    .Q(\datamem.data_ram[45][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30817_ (.CLK(clk),
    .D(_02552_),
    .Q(\datamem.data_ram[45][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30818_ (.CLK(clk),
    .D(_02553_),
    .Q(\datamem.data_ram[45][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30819_ (.CLK(clk),
    .D(_02554_),
    .Q(\datamem.data_ram[45][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30820_ (.CLK(clk),
    .D(_02555_),
    .Q(\datamem.data_ram[45][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30821_ (.CLK(clk),
    .D(_02556_),
    .Q(\datamem.data_ram[44][24] ));
 sky130_fd_sc_hd__dfxtp_1 _30822_ (.CLK(clk),
    .D(_02557_),
    .Q(\datamem.data_ram[44][25] ));
 sky130_fd_sc_hd__dfxtp_1 _30823_ (.CLK(clk),
    .D(_02558_),
    .Q(\datamem.data_ram[44][26] ));
 sky130_fd_sc_hd__dfxtp_1 _30824_ (.CLK(clk),
    .D(_02559_),
    .Q(\datamem.data_ram[44][27] ));
 sky130_fd_sc_hd__dfxtp_1 _30825_ (.CLK(clk),
    .D(_02560_),
    .Q(\datamem.data_ram[44][28] ));
 sky130_fd_sc_hd__dfxtp_1 _30826_ (.CLK(clk),
    .D(_02561_),
    .Q(\datamem.data_ram[44][29] ));
 sky130_fd_sc_hd__dfxtp_1 _30827_ (.CLK(clk),
    .D(_02562_),
    .Q(\datamem.data_ram[44][30] ));
 sky130_fd_sc_hd__dfxtp_1 _30828_ (.CLK(clk),
    .D(_02563_),
    .Q(\datamem.data_ram[44][31] ));
 sky130_fd_sc_hd__dfxtp_1 _30829_ (.CLK(clk),
    .D(_02564_),
    .Q(\datamem.data_ram[44][16] ));
 sky130_fd_sc_hd__dfxtp_1 _30830_ (.CLK(clk),
    .D(_02565_),
    .Q(\datamem.data_ram[44][17] ));
 sky130_fd_sc_hd__dfxtp_1 _30831_ (.CLK(clk),
    .D(_02566_),
    .Q(\datamem.data_ram[44][18] ));
 sky130_fd_sc_hd__dfxtp_1 _30832_ (.CLK(clk),
    .D(_02567_),
    .Q(\datamem.data_ram[44][19] ));
 sky130_fd_sc_hd__dfxtp_1 _30833_ (.CLK(clk),
    .D(_02568_),
    .Q(\datamem.data_ram[44][20] ));
 sky130_fd_sc_hd__dfxtp_1 _30834_ (.CLK(clk),
    .D(_02569_),
    .Q(\datamem.data_ram[44][21] ));
 sky130_fd_sc_hd__dfxtp_1 _30835_ (.CLK(clk),
    .D(_02570_),
    .Q(\datamem.data_ram[44][22] ));
 sky130_fd_sc_hd__dfxtp_1 _30836_ (.CLK(clk),
    .D(_02571_),
    .Q(\datamem.data_ram[44][23] ));
 sky130_fd_sc_hd__dfxtp_1 _30837_ (.CLK(clk),
    .D(_02572_),
    .Q(\datamem.data_ram[44][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30838_ (.CLK(clk),
    .D(_02573_),
    .Q(\datamem.data_ram[44][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30839_ (.CLK(clk),
    .D(_02574_),
    .Q(\datamem.data_ram[44][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30840_ (.CLK(clk),
    .D(_02575_),
    .Q(\datamem.data_ram[44][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30841_ (.CLK(clk),
    .D(_02576_),
    .Q(\datamem.data_ram[44][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30842_ (.CLK(clk),
    .D(_02577_),
    .Q(\datamem.data_ram[44][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30843_ (.CLK(clk),
    .D(_02578_),
    .Q(\datamem.data_ram[44][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30844_ (.CLK(clk),
    .D(_02579_),
    .Q(\datamem.data_ram[44][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30845_ (.CLK(clk),
    .D(_02580_),
    .Q(\datamem.data_ram[43][24] ));
 sky130_fd_sc_hd__dfxtp_1 _30846_ (.CLK(clk),
    .D(_02581_),
    .Q(\datamem.data_ram[43][25] ));
 sky130_fd_sc_hd__dfxtp_1 _30847_ (.CLK(clk),
    .D(_02582_),
    .Q(\datamem.data_ram[43][26] ));
 sky130_fd_sc_hd__dfxtp_1 _30848_ (.CLK(clk),
    .D(_02583_),
    .Q(\datamem.data_ram[43][27] ));
 sky130_fd_sc_hd__dfxtp_1 _30849_ (.CLK(clk),
    .D(_02584_),
    .Q(\datamem.data_ram[43][28] ));
 sky130_fd_sc_hd__dfxtp_1 _30850_ (.CLK(clk),
    .D(_02585_),
    .Q(\datamem.data_ram[43][29] ));
 sky130_fd_sc_hd__dfxtp_1 _30851_ (.CLK(clk),
    .D(_02586_),
    .Q(\datamem.data_ram[43][30] ));
 sky130_fd_sc_hd__dfxtp_1 _30852_ (.CLK(clk),
    .D(_02587_),
    .Q(\datamem.data_ram[43][31] ));
 sky130_fd_sc_hd__dfxtp_1 _30853_ (.CLK(clk),
    .D(_02588_),
    .Q(\datamem.data_ram[43][16] ));
 sky130_fd_sc_hd__dfxtp_1 _30854_ (.CLK(clk),
    .D(_02589_),
    .Q(\datamem.data_ram[43][17] ));
 sky130_fd_sc_hd__dfxtp_1 _30855_ (.CLK(clk),
    .D(_02590_),
    .Q(\datamem.data_ram[43][18] ));
 sky130_fd_sc_hd__dfxtp_1 _30856_ (.CLK(clk),
    .D(_02591_),
    .Q(\datamem.data_ram[43][19] ));
 sky130_fd_sc_hd__dfxtp_1 _30857_ (.CLK(clk),
    .D(_02592_),
    .Q(\datamem.data_ram[43][20] ));
 sky130_fd_sc_hd__dfxtp_1 _30858_ (.CLK(clk),
    .D(_02593_),
    .Q(\datamem.data_ram[43][21] ));
 sky130_fd_sc_hd__dfxtp_1 _30859_ (.CLK(clk),
    .D(_02594_),
    .Q(\datamem.data_ram[43][22] ));
 sky130_fd_sc_hd__dfxtp_1 _30860_ (.CLK(clk),
    .D(_02595_),
    .Q(\datamem.data_ram[43][23] ));
 sky130_fd_sc_hd__dfxtp_1 _30861_ (.CLK(clk),
    .D(_02596_),
    .Q(\datamem.data_ram[43][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30862_ (.CLK(clk),
    .D(_02597_),
    .Q(\datamem.data_ram[43][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30863_ (.CLK(clk),
    .D(_02598_),
    .Q(\datamem.data_ram[43][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30864_ (.CLK(clk),
    .D(_02599_),
    .Q(\datamem.data_ram[43][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30865_ (.CLK(clk),
    .D(_02600_),
    .Q(\datamem.data_ram[43][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30866_ (.CLK(clk),
    .D(_02601_),
    .Q(\datamem.data_ram[43][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30867_ (.CLK(clk),
    .D(_02602_),
    .Q(\datamem.data_ram[43][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30868_ (.CLK(clk),
    .D(_02603_),
    .Q(\datamem.data_ram[43][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30869_ (.CLK(clk),
    .D(_02604_),
    .Q(\datamem.data_ram[42][0] ));
 sky130_fd_sc_hd__dfxtp_1 _30870_ (.CLK(clk),
    .D(_02605_),
    .Q(\datamem.data_ram[42][1] ));
 sky130_fd_sc_hd__dfxtp_1 _30871_ (.CLK(clk),
    .D(_02606_),
    .Q(\datamem.data_ram[42][2] ));
 sky130_fd_sc_hd__dfxtp_1 _30872_ (.CLK(clk),
    .D(_02607_),
    .Q(\datamem.data_ram[42][3] ));
 sky130_fd_sc_hd__dfxtp_1 _30873_ (.CLK(clk),
    .D(_02608_),
    .Q(\datamem.data_ram[42][4] ));
 sky130_fd_sc_hd__dfxtp_1 _30874_ (.CLK(clk),
    .D(_02609_),
    .Q(\datamem.data_ram[42][5] ));
 sky130_fd_sc_hd__dfxtp_1 _30875_ (.CLK(clk),
    .D(_02610_),
    .Q(\datamem.data_ram[42][6] ));
 sky130_fd_sc_hd__dfxtp_1 _30876_ (.CLK(clk),
    .D(_02611_),
    .Q(\datamem.data_ram[42][7] ));
 sky130_fd_sc_hd__dfxtp_1 _30877_ (.CLK(clk),
    .D(_02612_),
    .Q(\datamem.data_ram[42][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30878_ (.CLK(clk),
    .D(_02613_),
    .Q(\datamem.data_ram[42][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30879_ (.CLK(clk),
    .D(_02614_),
    .Q(\datamem.data_ram[42][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30880_ (.CLK(clk),
    .D(_02615_),
    .Q(\datamem.data_ram[42][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30881_ (.CLK(clk),
    .D(_02616_),
    .Q(\datamem.data_ram[42][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30882_ (.CLK(clk),
    .D(_02617_),
    .Q(\datamem.data_ram[42][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30883_ (.CLK(clk),
    .D(_02618_),
    .Q(\datamem.data_ram[42][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30884_ (.CLK(clk),
    .D(_02619_),
    .Q(\datamem.data_ram[42][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30885_ (.CLK(clk),
    .D(_02620_),
    .Q(\datamem.data_ram[42][24] ));
 sky130_fd_sc_hd__dfxtp_1 _30886_ (.CLK(clk),
    .D(_02621_),
    .Q(\datamem.data_ram[42][25] ));
 sky130_fd_sc_hd__dfxtp_1 _30887_ (.CLK(clk),
    .D(_02622_),
    .Q(\datamem.data_ram[42][26] ));
 sky130_fd_sc_hd__dfxtp_1 _30888_ (.CLK(clk),
    .D(_02623_),
    .Q(\datamem.data_ram[42][27] ));
 sky130_fd_sc_hd__dfxtp_1 _30889_ (.CLK(clk),
    .D(_02624_),
    .Q(\datamem.data_ram[42][28] ));
 sky130_fd_sc_hd__dfxtp_1 _30890_ (.CLK(clk),
    .D(_02625_),
    .Q(\datamem.data_ram[42][29] ));
 sky130_fd_sc_hd__dfxtp_1 _30891_ (.CLK(clk),
    .D(_02626_),
    .Q(\datamem.data_ram[42][30] ));
 sky130_fd_sc_hd__dfxtp_1 _30892_ (.CLK(clk),
    .D(_02627_),
    .Q(\datamem.data_ram[42][31] ));
 sky130_fd_sc_hd__dfxtp_1 _30893_ (.CLK(clk),
    .D(_02628_),
    .Q(\datamem.data_ram[41][16] ));
 sky130_fd_sc_hd__dfxtp_1 _30894_ (.CLK(clk),
    .D(_02629_),
    .Q(\datamem.data_ram[41][17] ));
 sky130_fd_sc_hd__dfxtp_1 _30895_ (.CLK(clk),
    .D(_02630_),
    .Q(\datamem.data_ram[41][18] ));
 sky130_fd_sc_hd__dfxtp_1 _30896_ (.CLK(clk),
    .D(_02631_),
    .Q(\datamem.data_ram[41][19] ));
 sky130_fd_sc_hd__dfxtp_1 _30897_ (.CLK(clk),
    .D(_02632_),
    .Q(\datamem.data_ram[41][20] ));
 sky130_fd_sc_hd__dfxtp_1 _30898_ (.CLK(clk),
    .D(_02633_),
    .Q(\datamem.data_ram[41][21] ));
 sky130_fd_sc_hd__dfxtp_1 _30899_ (.CLK(clk),
    .D(_02634_),
    .Q(\datamem.data_ram[41][22] ));
 sky130_fd_sc_hd__dfxtp_1 _30900_ (.CLK(clk),
    .D(_02635_),
    .Q(\datamem.data_ram[41][23] ));
 sky130_fd_sc_hd__dfxtp_1 _30901_ (.CLK(clk),
    .D(_02636_),
    .Q(\datamem.data_ram[41][24] ));
 sky130_fd_sc_hd__dfxtp_1 _30902_ (.CLK(clk),
    .D(_02637_),
    .Q(\datamem.data_ram[41][25] ));
 sky130_fd_sc_hd__dfxtp_1 _30903_ (.CLK(clk),
    .D(_02638_),
    .Q(\datamem.data_ram[41][26] ));
 sky130_fd_sc_hd__dfxtp_1 _30904_ (.CLK(clk),
    .D(_02639_),
    .Q(\datamem.data_ram[41][27] ));
 sky130_fd_sc_hd__dfxtp_1 _30905_ (.CLK(clk),
    .D(_02640_),
    .Q(\datamem.data_ram[41][28] ));
 sky130_fd_sc_hd__dfxtp_1 _30906_ (.CLK(clk),
    .D(_02641_),
    .Q(\datamem.data_ram[41][29] ));
 sky130_fd_sc_hd__dfxtp_1 _30907_ (.CLK(clk),
    .D(_02642_),
    .Q(\datamem.data_ram[41][30] ));
 sky130_fd_sc_hd__dfxtp_1 _30908_ (.CLK(clk),
    .D(_02643_),
    .Q(\datamem.data_ram[41][31] ));
 sky130_fd_sc_hd__dfxtp_1 _30909_ (.CLK(clk),
    .D(_02644_),
    .Q(\datamem.data_ram[41][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30910_ (.CLK(clk),
    .D(_02645_),
    .Q(\datamem.data_ram[41][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30911_ (.CLK(clk),
    .D(_02646_),
    .Q(\datamem.data_ram[41][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30912_ (.CLK(clk),
    .D(_02647_),
    .Q(\datamem.data_ram[41][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30913_ (.CLK(clk),
    .D(_02648_),
    .Q(\datamem.data_ram[41][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30914_ (.CLK(clk),
    .D(_02649_),
    .Q(\datamem.data_ram[41][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30915_ (.CLK(clk),
    .D(_02650_),
    .Q(\datamem.data_ram[41][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30916_ (.CLK(clk),
    .D(_02651_),
    .Q(\datamem.data_ram[41][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30917_ (.CLK(clk),
    .D(_02652_),
    .Q(\datamem.data_ram[40][24] ));
 sky130_fd_sc_hd__dfxtp_1 _30918_ (.CLK(clk),
    .D(_02653_),
    .Q(\datamem.data_ram[40][25] ));
 sky130_fd_sc_hd__dfxtp_1 _30919_ (.CLK(clk),
    .D(_02654_),
    .Q(\datamem.data_ram[40][26] ));
 sky130_fd_sc_hd__dfxtp_1 _30920_ (.CLK(clk),
    .D(_02655_),
    .Q(\datamem.data_ram[40][27] ));
 sky130_fd_sc_hd__dfxtp_1 _30921_ (.CLK(clk),
    .D(_02656_),
    .Q(\datamem.data_ram[40][28] ));
 sky130_fd_sc_hd__dfxtp_1 _30922_ (.CLK(clk),
    .D(_02657_),
    .Q(\datamem.data_ram[40][29] ));
 sky130_fd_sc_hd__dfxtp_1 _30923_ (.CLK(clk),
    .D(_02658_),
    .Q(\datamem.data_ram[40][30] ));
 sky130_fd_sc_hd__dfxtp_1 _30924_ (.CLK(clk),
    .D(_02659_),
    .Q(\datamem.data_ram[40][31] ));
 sky130_fd_sc_hd__dfxtp_1 _30925_ (.CLK(clk),
    .D(_02660_),
    .Q(\datamem.data_ram[40][16] ));
 sky130_fd_sc_hd__dfxtp_1 _30926_ (.CLK(clk),
    .D(_02661_),
    .Q(\datamem.data_ram[40][17] ));
 sky130_fd_sc_hd__dfxtp_1 _30927_ (.CLK(clk),
    .D(_02662_),
    .Q(\datamem.data_ram[40][18] ));
 sky130_fd_sc_hd__dfxtp_1 _30928_ (.CLK(clk),
    .D(_02663_),
    .Q(\datamem.data_ram[40][19] ));
 sky130_fd_sc_hd__dfxtp_1 _30929_ (.CLK(clk),
    .D(_02664_),
    .Q(\datamem.data_ram[40][20] ));
 sky130_fd_sc_hd__dfxtp_1 _30930_ (.CLK(clk),
    .D(_02665_),
    .Q(\datamem.data_ram[40][21] ));
 sky130_fd_sc_hd__dfxtp_1 _30931_ (.CLK(clk),
    .D(_02666_),
    .Q(\datamem.data_ram[40][22] ));
 sky130_fd_sc_hd__dfxtp_1 _30932_ (.CLK(clk),
    .D(_02667_),
    .Q(\datamem.data_ram[40][23] ));
 sky130_fd_sc_hd__dfxtp_1 _30933_ (.CLK(clk),
    .D(_02668_),
    .Q(\datamem.data_ram[40][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30934_ (.CLK(clk),
    .D(_02669_),
    .Q(\datamem.data_ram[40][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30935_ (.CLK(clk),
    .D(_02670_),
    .Q(\datamem.data_ram[40][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30936_ (.CLK(clk),
    .D(_02671_),
    .Q(\datamem.data_ram[40][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30937_ (.CLK(clk),
    .D(_02672_),
    .Q(\datamem.data_ram[40][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30938_ (.CLK(clk),
    .D(_02673_),
    .Q(\datamem.data_ram[40][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30939_ (.CLK(clk),
    .D(_02674_),
    .Q(\datamem.data_ram[40][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30940_ (.CLK(clk),
    .D(_02675_),
    .Q(\datamem.data_ram[40][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30941_ (.CLK(clk),
    .D(_02676_),
    .Q(\datamem.data_ram[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _30942_ (.CLK(clk),
    .D(_02677_),
    .Q(\datamem.data_ram[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _30943_ (.CLK(clk),
    .D(_02678_),
    .Q(\datamem.data_ram[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _30944_ (.CLK(clk),
    .D(_02679_),
    .Q(\datamem.data_ram[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _30945_ (.CLK(clk),
    .D(_02680_),
    .Q(\datamem.data_ram[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _30946_ (.CLK(clk),
    .D(_02681_),
    .Q(\datamem.data_ram[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _30947_ (.CLK(clk),
    .D(_02682_),
    .Q(\datamem.data_ram[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _30948_ (.CLK(clk),
    .D(_02683_),
    .Q(\datamem.data_ram[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _30949_ (.CLK(clk),
    .D(_02684_),
    .Q(\datamem.data_ram[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30950_ (.CLK(clk),
    .D(_02685_),
    .Q(\datamem.data_ram[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30951_ (.CLK(clk),
    .D(_02686_),
    .Q(\datamem.data_ram[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30952_ (.CLK(clk),
    .D(_02687_),
    .Q(\datamem.data_ram[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30953_ (.CLK(clk),
    .D(_02688_),
    .Q(\datamem.data_ram[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30954_ (.CLK(clk),
    .D(_02689_),
    .Q(\datamem.data_ram[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30955_ (.CLK(clk),
    .D(_02690_),
    .Q(\datamem.data_ram[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30956_ (.CLK(clk),
    .D(_02691_),
    .Q(\datamem.data_ram[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30957_ (.CLK(clk),
    .D(_02692_),
    .Q(\datamem.data_ram[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 _30958_ (.CLK(clk),
    .D(_02693_),
    .Q(\datamem.data_ram[3][17] ));
 sky130_fd_sc_hd__dfxtp_1 _30959_ (.CLK(clk),
    .D(_02694_),
    .Q(\datamem.data_ram[3][18] ));
 sky130_fd_sc_hd__dfxtp_1 _30960_ (.CLK(clk),
    .D(_02695_),
    .Q(\datamem.data_ram[3][19] ));
 sky130_fd_sc_hd__dfxtp_1 _30961_ (.CLK(clk),
    .D(_02696_),
    .Q(\datamem.data_ram[3][20] ));
 sky130_fd_sc_hd__dfxtp_1 _30962_ (.CLK(clk),
    .D(_02697_),
    .Q(\datamem.data_ram[3][21] ));
 sky130_fd_sc_hd__dfxtp_1 _30963_ (.CLK(clk),
    .D(_02698_),
    .Q(\datamem.data_ram[3][22] ));
 sky130_fd_sc_hd__dfxtp_1 _30964_ (.CLK(clk),
    .D(_02699_),
    .Q(\datamem.data_ram[3][23] ));
 sky130_fd_sc_hd__dfxtp_1 _30965_ (.CLK(clk),
    .D(_02700_),
    .Q(\datamem.data_ram[39][24] ));
 sky130_fd_sc_hd__dfxtp_1 _30966_ (.CLK(clk),
    .D(_02701_),
    .Q(\datamem.data_ram[39][25] ));
 sky130_fd_sc_hd__dfxtp_1 _30967_ (.CLK(clk),
    .D(_02702_),
    .Q(\datamem.data_ram[39][26] ));
 sky130_fd_sc_hd__dfxtp_1 _30968_ (.CLK(clk),
    .D(_02703_),
    .Q(\datamem.data_ram[39][27] ));
 sky130_fd_sc_hd__dfxtp_1 _30969_ (.CLK(clk),
    .D(_02704_),
    .Q(\datamem.data_ram[39][28] ));
 sky130_fd_sc_hd__dfxtp_1 _30970_ (.CLK(clk),
    .D(_02705_),
    .Q(\datamem.data_ram[39][29] ));
 sky130_fd_sc_hd__dfxtp_1 _30971_ (.CLK(clk),
    .D(_02706_),
    .Q(\datamem.data_ram[39][30] ));
 sky130_fd_sc_hd__dfxtp_1 _30972_ (.CLK(clk),
    .D(_02707_),
    .Q(\datamem.data_ram[39][31] ));
 sky130_fd_sc_hd__dfxtp_1 _30973_ (.CLK(clk),
    .D(_02708_),
    .Q(\datamem.data_ram[39][16] ));
 sky130_fd_sc_hd__dfxtp_1 _30974_ (.CLK(clk),
    .D(_02709_),
    .Q(\datamem.data_ram[39][17] ));
 sky130_fd_sc_hd__dfxtp_1 _30975_ (.CLK(clk),
    .D(_02710_),
    .Q(\datamem.data_ram[39][18] ));
 sky130_fd_sc_hd__dfxtp_1 _30976_ (.CLK(clk),
    .D(_02711_),
    .Q(\datamem.data_ram[39][19] ));
 sky130_fd_sc_hd__dfxtp_1 _30977_ (.CLK(clk),
    .D(_02712_),
    .Q(\datamem.data_ram[39][20] ));
 sky130_fd_sc_hd__dfxtp_1 _30978_ (.CLK(clk),
    .D(_02713_),
    .Q(\datamem.data_ram[39][21] ));
 sky130_fd_sc_hd__dfxtp_1 _30979_ (.CLK(clk),
    .D(_02714_),
    .Q(\datamem.data_ram[39][22] ));
 sky130_fd_sc_hd__dfxtp_1 _30980_ (.CLK(clk),
    .D(_02715_),
    .Q(\datamem.data_ram[39][23] ));
 sky130_fd_sc_hd__dfxtp_1 _30981_ (.CLK(clk),
    .D(_02716_),
    .Q(\datamem.data_ram[39][0] ));
 sky130_fd_sc_hd__dfxtp_1 _30982_ (.CLK(clk),
    .D(_02717_),
    .Q(\datamem.data_ram[39][1] ));
 sky130_fd_sc_hd__dfxtp_1 _30983_ (.CLK(clk),
    .D(_02718_),
    .Q(\datamem.data_ram[39][2] ));
 sky130_fd_sc_hd__dfxtp_1 _30984_ (.CLK(clk),
    .D(_02719_),
    .Q(\datamem.data_ram[39][3] ));
 sky130_fd_sc_hd__dfxtp_1 _30985_ (.CLK(clk),
    .D(_02720_),
    .Q(\datamem.data_ram[39][4] ));
 sky130_fd_sc_hd__dfxtp_1 _30986_ (.CLK(clk),
    .D(_02721_),
    .Q(\datamem.data_ram[39][5] ));
 sky130_fd_sc_hd__dfxtp_1 _30987_ (.CLK(clk),
    .D(_02722_),
    .Q(\datamem.data_ram[39][6] ));
 sky130_fd_sc_hd__dfxtp_1 _30988_ (.CLK(clk),
    .D(_02723_),
    .Q(\datamem.data_ram[39][7] ));
 sky130_fd_sc_hd__dfxtp_1 _30989_ (.CLK(clk),
    .D(_02724_),
    .Q(\datamem.data_ram[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _30990_ (.CLK(clk),
    .D(_02725_),
    .Q(\datamem.data_ram[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _30991_ (.CLK(clk),
    .D(_02726_),
    .Q(\datamem.data_ram[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _30992_ (.CLK(clk),
    .D(_02727_),
    .Q(\datamem.data_ram[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _30993_ (.CLK(clk),
    .D(_02728_),
    .Q(\datamem.data_ram[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _30994_ (.CLK(clk),
    .D(_02729_),
    .Q(\datamem.data_ram[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _30995_ (.CLK(clk),
    .D(_02730_),
    .Q(\datamem.data_ram[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _30996_ (.CLK(clk),
    .D(_02731_),
    .Q(\datamem.data_ram[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _30997_ (.CLK(clk),
    .D(_02732_),
    .Q(\datamem.data_ram[22][0] ));
 sky130_fd_sc_hd__dfxtp_1 _30998_ (.CLK(clk),
    .D(_02733_),
    .Q(\datamem.data_ram[22][1] ));
 sky130_fd_sc_hd__dfxtp_1 _30999_ (.CLK(clk),
    .D(_02734_),
    .Q(\datamem.data_ram[22][2] ));
 sky130_fd_sc_hd__dfxtp_1 _31000_ (.CLK(clk),
    .D(_02735_),
    .Q(\datamem.data_ram[22][3] ));
 sky130_fd_sc_hd__dfxtp_1 _31001_ (.CLK(clk),
    .D(_02736_),
    .Q(\datamem.data_ram[22][4] ));
 sky130_fd_sc_hd__dfxtp_1 _31002_ (.CLK(clk),
    .D(_02737_),
    .Q(\datamem.data_ram[22][5] ));
 sky130_fd_sc_hd__dfxtp_1 _31003_ (.CLK(clk),
    .D(_02738_),
    .Q(\datamem.data_ram[22][6] ));
 sky130_fd_sc_hd__dfxtp_1 _31004_ (.CLK(clk),
    .D(_02739_),
    .Q(\datamem.data_ram[22][7] ));
 sky130_fd_sc_hd__dfxtp_1 _31005_ (.CLK(clk),
    .D(_02740_),
    .Q(\datamem.data_ram[11][16] ));
 sky130_fd_sc_hd__dfxtp_1 _31006_ (.CLK(clk),
    .D(_02741_),
    .Q(\datamem.data_ram[11][17] ));
 sky130_fd_sc_hd__dfxtp_1 _31007_ (.CLK(clk),
    .D(_02742_),
    .Q(\datamem.data_ram[11][18] ));
 sky130_fd_sc_hd__dfxtp_1 _31008_ (.CLK(clk),
    .D(_02743_),
    .Q(\datamem.data_ram[11][19] ));
 sky130_fd_sc_hd__dfxtp_1 _31009_ (.CLK(clk),
    .D(_02744_),
    .Q(\datamem.data_ram[11][20] ));
 sky130_fd_sc_hd__dfxtp_1 _31010_ (.CLK(clk),
    .D(_02745_),
    .Q(\datamem.data_ram[11][21] ));
 sky130_fd_sc_hd__dfxtp_1 _31011_ (.CLK(clk),
    .D(_02746_),
    .Q(\datamem.data_ram[11][22] ));
 sky130_fd_sc_hd__dfxtp_1 _31012_ (.CLK(clk),
    .D(_02747_),
    .Q(\datamem.data_ram[11][23] ));
 sky130_fd_sc_hd__dfxtp_1 _31013_ (.CLK(clk),
    .D(_02748_),
    .Q(\datamem.data_ram[42][16] ));
 sky130_fd_sc_hd__dfxtp_1 _31014_ (.CLK(clk),
    .D(_02749_),
    .Q(\datamem.data_ram[42][17] ));
 sky130_fd_sc_hd__dfxtp_1 _31015_ (.CLK(clk),
    .D(_02750_),
    .Q(\datamem.data_ram[42][18] ));
 sky130_fd_sc_hd__dfxtp_1 _31016_ (.CLK(clk),
    .D(_02751_),
    .Q(\datamem.data_ram[42][19] ));
 sky130_fd_sc_hd__dfxtp_1 _31017_ (.CLK(clk),
    .D(_02752_),
    .Q(\datamem.data_ram[42][20] ));
 sky130_fd_sc_hd__dfxtp_1 _31018_ (.CLK(clk),
    .D(_02753_),
    .Q(\datamem.data_ram[42][21] ));
 sky130_fd_sc_hd__dfxtp_1 _31019_ (.CLK(clk),
    .D(_02754_),
    .Q(\datamem.data_ram[42][22] ));
 sky130_fd_sc_hd__dfxtp_1 _31020_ (.CLK(clk),
    .D(_02755_),
    .Q(\datamem.data_ram[42][23] ));
 sky130_fd_sc_hd__dfxtp_1 _31021_ (.CLK(clk),
    .D(_02756_),
    .Q(\datamem.data_ram[40][0] ));
 sky130_fd_sc_hd__dfxtp_1 _31022_ (.CLK(clk),
    .D(_02757_),
    .Q(\datamem.data_ram[40][1] ));
 sky130_fd_sc_hd__dfxtp_1 _31023_ (.CLK(clk),
    .D(_02758_),
    .Q(\datamem.data_ram[40][2] ));
 sky130_fd_sc_hd__dfxtp_1 _31024_ (.CLK(clk),
    .D(_02759_),
    .Q(\datamem.data_ram[40][3] ));
 sky130_fd_sc_hd__dfxtp_1 _31025_ (.CLK(clk),
    .D(_02760_),
    .Q(\datamem.data_ram[40][4] ));
 sky130_fd_sc_hd__dfxtp_1 _31026_ (.CLK(clk),
    .D(_02761_),
    .Q(\datamem.data_ram[40][5] ));
 sky130_fd_sc_hd__dfxtp_1 _31027_ (.CLK(clk),
    .D(_02762_),
    .Q(\datamem.data_ram[40][6] ));
 sky130_fd_sc_hd__dfxtp_1 _31028_ (.CLK(clk),
    .D(_02763_),
    .Q(\datamem.data_ram[40][7] ));
 sky130_fd_sc_hd__dfxtp_1 _31029_ (.CLK(clk),
    .D(_02764_),
    .Q(\datamem.data_ram[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _31030_ (.CLK(clk),
    .D(_02765_),
    .Q(\datamem.data_ram[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _31031_ (.CLK(clk),
    .D(_02766_),
    .Q(\datamem.data_ram[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _31032_ (.CLK(clk),
    .D(_02767_),
    .Q(\datamem.data_ram[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _31033_ (.CLK(clk),
    .D(_02768_),
    .Q(\datamem.data_ram[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _31034_ (.CLK(clk),
    .D(_02769_),
    .Q(\datamem.data_ram[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _31035_ (.CLK(clk),
    .D(_02770_),
    .Q(\datamem.data_ram[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _31036_ (.CLK(clk),
    .D(_02771_),
    .Q(\datamem.data_ram[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _31037_ (.CLK(clk),
    .D(_02772_),
    .Q(\datamem.data_ram[41][0] ));
 sky130_fd_sc_hd__dfxtp_1 _31038_ (.CLK(clk),
    .D(_02773_),
    .Q(\datamem.data_ram[41][1] ));
 sky130_fd_sc_hd__dfxtp_1 _31039_ (.CLK(clk),
    .D(_02774_),
    .Q(\datamem.data_ram[41][2] ));
 sky130_fd_sc_hd__dfxtp_1 _31040_ (.CLK(clk),
    .D(_02775_),
    .Q(\datamem.data_ram[41][3] ));
 sky130_fd_sc_hd__dfxtp_1 _31041_ (.CLK(clk),
    .D(_02776_),
    .Q(\datamem.data_ram[41][4] ));
 sky130_fd_sc_hd__dfxtp_1 _31042_ (.CLK(clk),
    .D(_02777_),
    .Q(\datamem.data_ram[41][5] ));
 sky130_fd_sc_hd__dfxtp_1 _31043_ (.CLK(clk),
    .D(_02778_),
    .Q(\datamem.data_ram[41][6] ));
 sky130_fd_sc_hd__dfxtp_1 _31044_ (.CLK(clk),
    .D(_02779_),
    .Q(\datamem.data_ram[41][7] ));
 sky130_fd_sc_hd__dfxtp_1 _31045_ (.CLK(clk),
    .D(_02780_),
    .Q(\datamem.data_ram[9][24] ));
 sky130_fd_sc_hd__dfxtp_1 _31046_ (.CLK(clk),
    .D(_02781_),
    .Q(\datamem.data_ram[9][25] ));
 sky130_fd_sc_hd__dfxtp_1 _31047_ (.CLK(clk),
    .D(_02782_),
    .Q(\datamem.data_ram[9][26] ));
 sky130_fd_sc_hd__dfxtp_1 _31048_ (.CLK(clk),
    .D(_02783_),
    .Q(\datamem.data_ram[9][27] ));
 sky130_fd_sc_hd__dfxtp_1 _31049_ (.CLK(clk),
    .D(_02784_),
    .Q(\datamem.data_ram[9][28] ));
 sky130_fd_sc_hd__dfxtp_1 _31050_ (.CLK(clk),
    .D(_02785_),
    .Q(\datamem.data_ram[9][29] ));
 sky130_fd_sc_hd__dfxtp_1 _31051_ (.CLK(clk),
    .D(_02786_),
    .Q(\datamem.data_ram[9][30] ));
 sky130_fd_sc_hd__dfxtp_1 _31052_ (.CLK(clk),
    .D(_02787_),
    .Q(\datamem.data_ram[9][31] ));
 sky130_fd_sc_hd__dfxtp_1 _31053_ (.CLK(clk),
    .D(_02788_),
    .Q(\datamem.data_ram[38][0] ));
 sky130_fd_sc_hd__dfxtp_1 _31054_ (.CLK(clk),
    .D(_02789_),
    .Q(\datamem.data_ram[38][1] ));
 sky130_fd_sc_hd__dfxtp_1 _31055_ (.CLK(clk),
    .D(_02790_),
    .Q(\datamem.data_ram[38][2] ));
 sky130_fd_sc_hd__dfxtp_1 _31056_ (.CLK(clk),
    .D(_02791_),
    .Q(\datamem.data_ram[38][3] ));
 sky130_fd_sc_hd__dfxtp_1 _31057_ (.CLK(clk),
    .D(_02792_),
    .Q(\datamem.data_ram[38][4] ));
 sky130_fd_sc_hd__dfxtp_1 _31058_ (.CLK(clk),
    .D(_02793_),
    .Q(\datamem.data_ram[38][5] ));
 sky130_fd_sc_hd__dfxtp_1 _31059_ (.CLK(clk),
    .D(_02794_),
    .Q(\datamem.data_ram[38][6] ));
 sky130_fd_sc_hd__dfxtp_1 _31060_ (.CLK(clk),
    .D(_02795_),
    .Q(\datamem.data_ram[38][7] ));
 sky130_fd_sc_hd__dfxtp_1 _31061_ (.CLK(clk),
    .D(_02796_),
    .Q(\datamem.data_ram[8][8] ));
 sky130_fd_sc_hd__dfxtp_1 _31062_ (.CLK(clk),
    .D(_02797_),
    .Q(\datamem.data_ram[8][9] ));
 sky130_fd_sc_hd__dfxtp_1 _31063_ (.CLK(clk),
    .D(_02798_),
    .Q(\datamem.data_ram[8][10] ));
 sky130_fd_sc_hd__dfxtp_1 _31064_ (.CLK(clk),
    .D(_02799_),
    .Q(\datamem.data_ram[8][11] ));
 sky130_fd_sc_hd__dfxtp_1 _31065_ (.CLK(clk),
    .D(_02800_),
    .Q(\datamem.data_ram[8][12] ));
 sky130_fd_sc_hd__dfxtp_1 _31066_ (.CLK(clk),
    .D(_02801_),
    .Q(\datamem.data_ram[8][13] ));
 sky130_fd_sc_hd__dfxtp_1 _31067_ (.CLK(clk),
    .D(_02802_),
    .Q(\datamem.data_ram[8][14] ));
 sky130_fd_sc_hd__dfxtp_1 _31068_ (.CLK(clk),
    .D(_02803_),
    .Q(\datamem.data_ram[8][15] ));
 sky130_fd_sc_hd__dfxtp_1 _31069_ (.CLK(clk),
    .D(_02804_),
    .Q(\datamem.data_ram[9][16] ));
 sky130_fd_sc_hd__dfxtp_1 _31070_ (.CLK(clk),
    .D(_02805_),
    .Q(\datamem.data_ram[9][17] ));
 sky130_fd_sc_hd__dfxtp_1 _31071_ (.CLK(clk),
    .D(_02806_),
    .Q(\datamem.data_ram[9][18] ));
 sky130_fd_sc_hd__dfxtp_1 _31072_ (.CLK(clk),
    .D(_02807_),
    .Q(\datamem.data_ram[9][19] ));
 sky130_fd_sc_hd__dfxtp_1 _31073_ (.CLK(clk),
    .D(_02808_),
    .Q(\datamem.data_ram[9][20] ));
 sky130_fd_sc_hd__dfxtp_1 _31074_ (.CLK(clk),
    .D(_02809_),
    .Q(\datamem.data_ram[9][21] ));
 sky130_fd_sc_hd__dfxtp_1 _31075_ (.CLK(clk),
    .D(_02810_),
    .Q(\datamem.data_ram[9][22] ));
 sky130_fd_sc_hd__dfxtp_1 _31076_ (.CLK(clk),
    .D(_02811_),
    .Q(\datamem.data_ram[9][23] ));
 sky130_fd_sc_hd__dfxtp_1 _31077_ (.CLK(clk),
    .D(_02812_),
    .Q(\datamem.data_ram[20][0] ));
 sky130_fd_sc_hd__dfxtp_1 _31078_ (.CLK(clk),
    .D(_02813_),
    .Q(\datamem.data_ram[20][1] ));
 sky130_fd_sc_hd__dfxtp_1 _31079_ (.CLK(clk),
    .D(_02814_),
    .Q(\datamem.data_ram[20][2] ));
 sky130_fd_sc_hd__dfxtp_1 _31080_ (.CLK(clk),
    .D(_02815_),
    .Q(\datamem.data_ram[20][3] ));
 sky130_fd_sc_hd__dfxtp_1 _31081_ (.CLK(clk),
    .D(_02816_),
    .Q(\datamem.data_ram[20][4] ));
 sky130_fd_sc_hd__dfxtp_1 _31082_ (.CLK(clk),
    .D(_02817_),
    .Q(\datamem.data_ram[20][5] ));
 sky130_fd_sc_hd__dfxtp_1 _31083_ (.CLK(clk),
    .D(_02818_),
    .Q(\datamem.data_ram[20][6] ));
 sky130_fd_sc_hd__dfxtp_1 _31084_ (.CLK(clk),
    .D(_02819_),
    .Q(\datamem.data_ram[20][7] ));
 sky130_fd_sc_hd__dfxtp_1 _31085_ (.CLK(clk),
    .D(_02820_),
    .Q(\datamem.data_ram[21][0] ));
 sky130_fd_sc_hd__dfxtp_1 _31086_ (.CLK(clk),
    .D(_02821_),
    .Q(\datamem.data_ram[21][1] ));
 sky130_fd_sc_hd__dfxtp_1 _31087_ (.CLK(clk),
    .D(_02822_),
    .Q(\datamem.data_ram[21][2] ));
 sky130_fd_sc_hd__dfxtp_1 _31088_ (.CLK(clk),
    .D(_02823_),
    .Q(\datamem.data_ram[21][3] ));
 sky130_fd_sc_hd__dfxtp_1 _31089_ (.CLK(clk),
    .D(_02824_),
    .Q(\datamem.data_ram[21][4] ));
 sky130_fd_sc_hd__dfxtp_1 _31090_ (.CLK(clk),
    .D(_02825_),
    .Q(\datamem.data_ram[21][5] ));
 sky130_fd_sc_hd__dfxtp_1 _31091_ (.CLK(clk),
    .D(_02826_),
    .Q(\datamem.data_ram[21][6] ));
 sky130_fd_sc_hd__dfxtp_1 _31092_ (.CLK(clk),
    .D(_02827_),
    .Q(\datamem.data_ram[21][7] ));
 sky130_fd_sc_hd__dfxtp_1 _31093_ (.CLK(clk),
    .D(_02828_),
    .Q(\datamem.data_ram[9][8] ));
 sky130_fd_sc_hd__dfxtp_1 _31094_ (.CLK(clk),
    .D(_02829_),
    .Q(\datamem.data_ram[9][9] ));
 sky130_fd_sc_hd__dfxtp_1 _31095_ (.CLK(clk),
    .D(_02830_),
    .Q(\datamem.data_ram[9][10] ));
 sky130_fd_sc_hd__dfxtp_1 _31096_ (.CLK(clk),
    .D(_02831_),
    .Q(\datamem.data_ram[9][11] ));
 sky130_fd_sc_hd__dfxtp_1 _31097_ (.CLK(clk),
    .D(_02832_),
    .Q(\datamem.data_ram[9][12] ));
 sky130_fd_sc_hd__dfxtp_1 _31098_ (.CLK(clk),
    .D(_02833_),
    .Q(\datamem.data_ram[9][13] ));
 sky130_fd_sc_hd__dfxtp_1 _31099_ (.CLK(clk),
    .D(_02834_),
    .Q(\datamem.data_ram[9][14] ));
 sky130_fd_sc_hd__dfxtp_1 _31100_ (.CLK(clk),
    .D(_02835_),
    .Q(\datamem.data_ram[9][15] ));
 sky130_fd_sc_hd__dfxtp_1 _31101_ (.CLK(clk),
    .D(_02836_),
    .Q(\datamem.data_ram[19][0] ));
 sky130_fd_sc_hd__dfxtp_1 _31102_ (.CLK(clk),
    .D(_02837_),
    .Q(\datamem.data_ram[19][1] ));
 sky130_fd_sc_hd__dfxtp_1 _31103_ (.CLK(clk),
    .D(_02838_),
    .Q(\datamem.data_ram[19][2] ));
 sky130_fd_sc_hd__dfxtp_1 _31104_ (.CLK(clk),
    .D(_02839_),
    .Q(\datamem.data_ram[19][3] ));
 sky130_fd_sc_hd__dfxtp_1 _31105_ (.CLK(clk),
    .D(_02840_),
    .Q(\datamem.data_ram[19][4] ));
 sky130_fd_sc_hd__dfxtp_1 _31106_ (.CLK(clk),
    .D(_02841_),
    .Q(\datamem.data_ram[19][5] ));
 sky130_fd_sc_hd__dfxtp_1 _31107_ (.CLK(clk),
    .D(_02842_),
    .Q(\datamem.data_ram[19][6] ));
 sky130_fd_sc_hd__dfxtp_1 _31108_ (.CLK(clk),
    .D(_02843_),
    .Q(\datamem.data_ram[19][7] ));
 sky130_fd_sc_hd__dfxtp_1 _31109_ (.CLK(clk),
    .D(_02844_),
    .Q(\datamem.data_ram[43][0] ));
 sky130_fd_sc_hd__dfxtp_1 _31110_ (.CLK(clk),
    .D(_02845_),
    .Q(\datamem.data_ram[43][1] ));
 sky130_fd_sc_hd__dfxtp_1 _31111_ (.CLK(clk),
    .D(_02846_),
    .Q(\datamem.data_ram[43][2] ));
 sky130_fd_sc_hd__dfxtp_1 _31112_ (.CLK(clk),
    .D(_02847_),
    .Q(\datamem.data_ram[43][3] ));
 sky130_fd_sc_hd__dfxtp_1 _31113_ (.CLK(clk),
    .D(_02848_),
    .Q(\datamem.data_ram[43][4] ));
 sky130_fd_sc_hd__dfxtp_1 _31114_ (.CLK(clk),
    .D(_02849_),
    .Q(\datamem.data_ram[43][5] ));
 sky130_fd_sc_hd__dfxtp_1 _31115_ (.CLK(clk),
    .D(_02850_),
    .Q(\datamem.data_ram[43][6] ));
 sky130_fd_sc_hd__dfxtp_1 _31116_ (.CLK(clk),
    .D(_02851_),
    .Q(\datamem.data_ram[43][7] ));
 sky130_fd_sc_hd__dfxtp_1 _31117_ (.CLK(clk),
    .D(_02852_),
    .Q(\datamem.data_ram[35][0] ));
 sky130_fd_sc_hd__dfxtp_1 _31118_ (.CLK(clk),
    .D(_02853_),
    .Q(\datamem.data_ram[35][1] ));
 sky130_fd_sc_hd__dfxtp_1 _31119_ (.CLK(clk),
    .D(_02854_),
    .Q(\datamem.data_ram[35][2] ));
 sky130_fd_sc_hd__dfxtp_1 _31120_ (.CLK(clk),
    .D(_02855_),
    .Q(\datamem.data_ram[35][3] ));
 sky130_fd_sc_hd__dfxtp_1 _31121_ (.CLK(clk),
    .D(_02856_),
    .Q(\datamem.data_ram[35][4] ));
 sky130_fd_sc_hd__dfxtp_1 _31122_ (.CLK(clk),
    .D(_02857_),
    .Q(\datamem.data_ram[35][5] ));
 sky130_fd_sc_hd__dfxtp_1 _31123_ (.CLK(clk),
    .D(_02858_),
    .Q(\datamem.data_ram[35][6] ));
 sky130_fd_sc_hd__dfxtp_1 _31124_ (.CLK(clk),
    .D(_02859_),
    .Q(\datamem.data_ram[35][7] ));
 sky130_fd_sc_hd__dfxtp_1 _31125_ (.CLK(clk),
    .D(_02860_),
    .Q(\datamem.data_ram[25][0] ));
 sky130_fd_sc_hd__dfxtp_1 _31126_ (.CLK(clk),
    .D(_02861_),
    .Q(\datamem.data_ram[25][1] ));
 sky130_fd_sc_hd__dfxtp_1 _31127_ (.CLK(clk),
    .D(_02862_),
    .Q(\datamem.data_ram[25][2] ));
 sky130_fd_sc_hd__dfxtp_1 _31128_ (.CLK(clk),
    .D(_02863_),
    .Q(\datamem.data_ram[25][3] ));
 sky130_fd_sc_hd__dfxtp_1 _31129_ (.CLK(clk),
    .D(_02864_),
    .Q(\datamem.data_ram[25][4] ));
 sky130_fd_sc_hd__dfxtp_1 _31130_ (.CLK(clk),
    .D(_02865_),
    .Q(\datamem.data_ram[25][5] ));
 sky130_fd_sc_hd__dfxtp_1 _31131_ (.CLK(clk),
    .D(_02866_),
    .Q(\datamem.data_ram[25][6] ));
 sky130_fd_sc_hd__dfxtp_1 _31132_ (.CLK(clk),
    .D(_02867_),
    .Q(\datamem.data_ram[25][7] ));
 sky130_fd_sc_hd__dfxtp_1 _31133_ (.CLK(clk),
    .D(_02868_),
    .Q(\datamem.data_ram[4][24] ));
 sky130_fd_sc_hd__dfxtp_1 _31134_ (.CLK(clk),
    .D(_02869_),
    .Q(\datamem.data_ram[4][25] ));
 sky130_fd_sc_hd__dfxtp_1 _31135_ (.CLK(clk),
    .D(_02870_),
    .Q(\datamem.data_ram[4][26] ));
 sky130_fd_sc_hd__dfxtp_1 _31136_ (.CLK(clk),
    .D(_02871_),
    .Q(\datamem.data_ram[4][27] ));
 sky130_fd_sc_hd__dfxtp_1 _31137_ (.CLK(clk),
    .D(_02872_),
    .Q(\datamem.data_ram[4][28] ));
 sky130_fd_sc_hd__dfxtp_1 _31138_ (.CLK(clk),
    .D(_02873_),
    .Q(\datamem.data_ram[4][29] ));
 sky130_fd_sc_hd__dfxtp_1 _31139_ (.CLK(clk),
    .D(_02874_),
    .Q(\datamem.data_ram[4][30] ));
 sky130_fd_sc_hd__dfxtp_1 _31140_ (.CLK(clk),
    .D(_02875_),
    .Q(\datamem.data_ram[4][31] ));
 sky130_fd_sc_hd__dfxtp_4 _31141_ (.CLK(clk),
    .D(\rvcpu.ALUResultE[0] ),
    .Q(\rvcpu.dp.plem.ALUResultM[0] ));
 sky130_fd_sc_hd__dfxtp_4 _31142_ (.CLK(clk),
    .D(\rvcpu.ALUResultE[1] ),
    .Q(\rvcpu.dp.plem.ALUResultM[1] ));
 sky130_fd_sc_hd__dfxtp_4 _31143_ (.CLK(clk),
    .D(\rvcpu.ALUResultE[2] ),
    .Q(\rvcpu.dp.plem.ALUResultM[2] ));
 sky130_fd_sc_hd__dfxtp_4 _31144_ (.CLK(clk),
    .D(\rvcpu.ALUResultE[3] ),
    .Q(\rvcpu.dp.plem.ALUResultM[3] ));
 sky130_fd_sc_hd__dfxtp_4 _31145_ (.CLK(clk),
    .D(\rvcpu.ALUResultE[4] ),
    .Q(\rvcpu.dp.plem.ALUResultM[4] ));
 sky130_fd_sc_hd__dfxtp_4 _31146_ (.CLK(clk),
    .D(\rvcpu.ALUResultE[5] ),
    .Q(\rvcpu.dp.plem.ALUResultM[5] ));
 sky130_fd_sc_hd__dfxtp_4 _31147_ (.CLK(clk),
    .D(\rvcpu.ALUResultE[6] ),
    .Q(\rvcpu.dp.plem.ALUResultM[6] ));
 sky130_fd_sc_hd__dfxtp_4 _31148_ (.CLK(clk),
    .D(\rvcpu.ALUResultE[7] ),
    .Q(\rvcpu.dp.plem.ALUResultM[7] ));
 sky130_fd_sc_hd__dfxtp_2 _31149_ (.CLK(clk),
    .D(\rvcpu.ALUResultE[8] ),
    .Q(\rvcpu.dp.plem.ALUResultM[8] ));
 sky130_fd_sc_hd__dfxtp_1 _31150_ (.CLK(clk),
    .D(\rvcpu.ALUResultE[9] ),
    .Q(\rvcpu.dp.plem.ALUResultM[9] ));
 sky130_fd_sc_hd__dfxtp_1 _31151_ (.CLK(clk),
    .D(\rvcpu.ALUResultE[10] ),
    .Q(\rvcpu.dp.plem.ALUResultM[10] ));
 sky130_fd_sc_hd__dfxtp_1 _31152_ (.CLK(clk),
    .D(\rvcpu.ALUResultE[11] ),
    .Q(\rvcpu.dp.plem.ALUResultM[11] ));
 sky130_fd_sc_hd__dfxtp_1 _31153_ (.CLK(clk),
    .D(\rvcpu.ALUResultE[12] ),
    .Q(\rvcpu.dp.plem.ALUResultM[12] ));
 sky130_fd_sc_hd__dfxtp_1 _31154_ (.CLK(clk),
    .D(\rvcpu.ALUResultE[13] ),
    .Q(\rvcpu.dp.plem.ALUResultM[13] ));
 sky130_fd_sc_hd__dfxtp_2 _31155_ (.CLK(clk),
    .D(\rvcpu.ALUResultE[14] ),
    .Q(\rvcpu.dp.plem.ALUResultM[14] ));
 sky130_fd_sc_hd__dfxtp_1 _31156_ (.CLK(clk),
    .D(\rvcpu.ALUResultE[15] ),
    .Q(\rvcpu.dp.plem.ALUResultM[15] ));
 sky130_fd_sc_hd__dfxtp_1 _31157_ (.CLK(clk),
    .D(\rvcpu.ALUResultE[16] ),
    .Q(\rvcpu.dp.plem.ALUResultM[16] ));
 sky130_fd_sc_hd__dfxtp_1 _31158_ (.CLK(clk),
    .D(\rvcpu.ALUResultE[17] ),
    .Q(\rvcpu.dp.plem.ALUResultM[17] ));
 sky130_fd_sc_hd__dfxtp_1 _31159_ (.CLK(clk),
    .D(\rvcpu.ALUResultE[18] ),
    .Q(\rvcpu.dp.plem.ALUResultM[18] ));
 sky130_fd_sc_hd__dfxtp_1 _31160_ (.CLK(clk),
    .D(\rvcpu.ALUResultE[19] ),
    .Q(\rvcpu.dp.plem.ALUResultM[19] ));
 sky130_fd_sc_hd__dfxtp_1 _31161_ (.CLK(clk),
    .D(\rvcpu.ALUResultE[20] ),
    .Q(\rvcpu.dp.plem.ALUResultM[20] ));
 sky130_fd_sc_hd__dfxtp_1 _31162_ (.CLK(clk),
    .D(\rvcpu.ALUResultE[21] ),
    .Q(\rvcpu.dp.plem.ALUResultM[21] ));
 sky130_fd_sc_hd__dfxtp_1 _31163_ (.CLK(clk),
    .D(\rvcpu.ALUResultE[22] ),
    .Q(\rvcpu.dp.plem.ALUResultM[22] ));
 sky130_fd_sc_hd__dfxtp_1 _31164_ (.CLK(clk),
    .D(\rvcpu.ALUResultE[23] ),
    .Q(\rvcpu.dp.plem.ALUResultM[23] ));
 sky130_fd_sc_hd__dfxtp_1 _31165_ (.CLK(clk),
    .D(\rvcpu.ALUResultE[24] ),
    .Q(\rvcpu.dp.plem.ALUResultM[24] ));
 sky130_fd_sc_hd__dfxtp_1 _31166_ (.CLK(clk),
    .D(\rvcpu.ALUResultE[25] ),
    .Q(\rvcpu.dp.plem.ALUResultM[25] ));
 sky130_fd_sc_hd__dfxtp_1 _31167_ (.CLK(clk),
    .D(\rvcpu.ALUResultE[26] ),
    .Q(\rvcpu.dp.plem.ALUResultM[26] ));
 sky130_fd_sc_hd__dfxtp_1 _31168_ (.CLK(clk),
    .D(\rvcpu.ALUResultE[27] ),
    .Q(\rvcpu.dp.plem.ALUResultM[27] ));
 sky130_fd_sc_hd__dfxtp_1 _31169_ (.CLK(clk),
    .D(\rvcpu.ALUResultE[28] ),
    .Q(\rvcpu.dp.plem.ALUResultM[28] ));
 sky130_fd_sc_hd__dfxtp_1 _31170_ (.CLK(clk),
    .D(\rvcpu.ALUResultE[29] ),
    .Q(\rvcpu.dp.plem.ALUResultM[29] ));
 sky130_fd_sc_hd__dfxtp_1 _31171_ (.CLK(clk),
    .D(\rvcpu.ALUResultE[30] ),
    .Q(\rvcpu.dp.plem.ALUResultM[30] ));
 sky130_fd_sc_hd__dfxtp_1 _31172_ (.CLK(clk),
    .D(\rvcpu.ALUResultE[31] ),
    .Q(\rvcpu.dp.plem.ALUResultM[31] ));
 sky130_fd_sc_hd__dfxtp_1 _31173_ (.CLK(clk),
    .D(_02876_),
    .Q(\datamem.data_ram[5][24] ));
 sky130_fd_sc_hd__dfxtp_1 _31174_ (.CLK(clk),
    .D(_02877_),
    .Q(\datamem.data_ram[5][25] ));
 sky130_fd_sc_hd__dfxtp_1 _31175_ (.CLK(clk),
    .D(_02878_),
    .Q(\datamem.data_ram[5][26] ));
 sky130_fd_sc_hd__dfxtp_1 _31176_ (.CLK(clk),
    .D(_02879_),
    .Q(\datamem.data_ram[5][27] ));
 sky130_fd_sc_hd__dfxtp_1 _31177_ (.CLK(clk),
    .D(_02880_),
    .Q(\datamem.data_ram[5][28] ));
 sky130_fd_sc_hd__dfxtp_1 _31178_ (.CLK(clk),
    .D(_02881_),
    .Q(\datamem.data_ram[5][29] ));
 sky130_fd_sc_hd__dfxtp_1 _31179_ (.CLK(clk),
    .D(_02882_),
    .Q(\datamem.data_ram[5][30] ));
 sky130_fd_sc_hd__dfxtp_1 _31180_ (.CLK(clk),
    .D(_02883_),
    .Q(\datamem.data_ram[5][31] ));
 sky130_fd_sc_hd__dfxtp_1 _31181_ (.CLK(clk),
    .D(_02884_),
    .Q(\rvcpu.dp.plfd.PCPlus4D[2] ));
 sky130_fd_sc_hd__dfxtp_1 _31182_ (.CLK(clk),
    .D(_02885_),
    .Q(\rvcpu.dp.plfd.PCPlus4D[3] ));
 sky130_fd_sc_hd__dfxtp_1 _31183_ (.CLK(clk),
    .D(_02886_),
    .Q(\rvcpu.dp.plfd.PCPlus4D[4] ));
 sky130_fd_sc_hd__dfxtp_1 _31184_ (.CLK(clk),
    .D(_02887_),
    .Q(\rvcpu.dp.plfd.PCPlus4D[5] ));
 sky130_fd_sc_hd__dfxtp_1 _31185_ (.CLK(clk),
    .D(_02888_),
    .Q(\rvcpu.dp.plfd.PCPlus4D[6] ));
 sky130_fd_sc_hd__dfxtp_1 _31186_ (.CLK(clk),
    .D(_02889_),
    .Q(\rvcpu.dp.plfd.PCPlus4D[7] ));
 sky130_fd_sc_hd__dfxtp_1 _31187_ (.CLK(clk),
    .D(_02890_),
    .Q(\rvcpu.dp.plfd.PCPlus4D[8] ));
 sky130_fd_sc_hd__dfxtp_1 _31188_ (.CLK(clk),
    .D(_02891_),
    .Q(\rvcpu.dp.plfd.PCPlus4D[9] ));
 sky130_fd_sc_hd__dfxtp_1 _31189_ (.CLK(clk),
    .D(_02892_),
    .Q(\rvcpu.dp.plfd.PCPlus4D[10] ));
 sky130_fd_sc_hd__dfxtp_1 _31190_ (.CLK(clk),
    .D(_02893_),
    .Q(\rvcpu.dp.plfd.PCPlus4D[11] ));
 sky130_fd_sc_hd__dfxtp_1 _31191_ (.CLK(clk),
    .D(_02894_),
    .Q(\rvcpu.dp.plfd.PCPlus4D[12] ));
 sky130_fd_sc_hd__dfxtp_1 _31192_ (.CLK(clk),
    .D(_02895_),
    .Q(\rvcpu.dp.plfd.PCPlus4D[13] ));
 sky130_fd_sc_hd__dfxtp_1 _31193_ (.CLK(clk),
    .D(_02896_),
    .Q(\rvcpu.dp.plfd.PCPlus4D[14] ));
 sky130_fd_sc_hd__dfxtp_1 _31194_ (.CLK(clk),
    .D(_02897_),
    .Q(\rvcpu.dp.plfd.PCPlus4D[15] ));
 sky130_fd_sc_hd__dfxtp_1 _31195_ (.CLK(clk),
    .D(_02898_),
    .Q(\rvcpu.dp.plfd.PCPlus4D[16] ));
 sky130_fd_sc_hd__dfxtp_1 _31196_ (.CLK(clk),
    .D(_02899_),
    .Q(\rvcpu.dp.plfd.PCPlus4D[17] ));
 sky130_fd_sc_hd__dfxtp_1 _31197_ (.CLK(clk),
    .D(_02900_),
    .Q(\rvcpu.dp.plfd.PCPlus4D[18] ));
 sky130_fd_sc_hd__dfxtp_1 _31198_ (.CLK(clk),
    .D(_02901_),
    .Q(\rvcpu.dp.plfd.PCPlus4D[19] ));
 sky130_fd_sc_hd__dfxtp_1 _31199_ (.CLK(clk),
    .D(_02902_),
    .Q(\rvcpu.dp.plfd.PCPlus4D[20] ));
 sky130_fd_sc_hd__dfxtp_1 _31200_ (.CLK(clk),
    .D(_02903_),
    .Q(\rvcpu.dp.plfd.PCPlus4D[21] ));
 sky130_fd_sc_hd__dfxtp_1 _31201_ (.CLK(clk),
    .D(_02904_),
    .Q(\rvcpu.dp.plfd.PCPlus4D[22] ));
 sky130_fd_sc_hd__dfxtp_1 _31202_ (.CLK(clk),
    .D(_02905_),
    .Q(\rvcpu.dp.plfd.PCPlus4D[23] ));
 sky130_fd_sc_hd__dfxtp_1 _31203_ (.CLK(clk),
    .D(_02906_),
    .Q(\rvcpu.dp.plfd.PCPlus4D[24] ));
 sky130_fd_sc_hd__dfxtp_1 _31204_ (.CLK(clk),
    .D(_02907_),
    .Q(\rvcpu.dp.plfd.PCPlus4D[25] ));
 sky130_fd_sc_hd__dfxtp_1 _31205_ (.CLK(clk),
    .D(_02908_),
    .Q(\rvcpu.dp.plfd.PCPlus4D[26] ));
 sky130_fd_sc_hd__dfxtp_1 _31206_ (.CLK(clk),
    .D(_02909_),
    .Q(\rvcpu.dp.plfd.PCPlus4D[27] ));
 sky130_fd_sc_hd__dfxtp_1 _31207_ (.CLK(clk),
    .D(_02910_),
    .Q(\rvcpu.dp.plfd.PCPlus4D[28] ));
 sky130_fd_sc_hd__dfxtp_1 _31208_ (.CLK(clk),
    .D(_02911_),
    .Q(\rvcpu.dp.plfd.PCPlus4D[29] ));
 sky130_fd_sc_hd__dfxtp_1 _31209_ (.CLK(clk),
    .D(_02912_),
    .Q(\rvcpu.dp.plfd.PCPlus4D[30] ));
 sky130_fd_sc_hd__dfxtp_1 _31210_ (.CLK(clk),
    .D(_02913_),
    .Q(\rvcpu.dp.plfd.PCPlus4D[31] ));
 sky130_fd_sc_hd__dfxtp_1 _31211_ (.CLK(clk),
    .D(_02914_),
    .Q(\rvcpu.dp.plfd.PCD[0] ));
 sky130_fd_sc_hd__dfxtp_1 _31212_ (.CLK(clk),
    .D(_02915_),
    .Q(\rvcpu.dp.plfd.PCD[1] ));
 sky130_fd_sc_hd__dfxtp_1 _31213_ (.CLK(clk),
    .D(_02916_),
    .Q(\rvcpu.dp.plfd.PCD[2] ));
 sky130_fd_sc_hd__dfxtp_1 _31214_ (.CLK(clk),
    .D(_02917_),
    .Q(\rvcpu.dp.plfd.PCD[3] ));
 sky130_fd_sc_hd__dfxtp_1 _31215_ (.CLK(clk),
    .D(_02918_),
    .Q(\rvcpu.dp.plfd.PCD[4] ));
 sky130_fd_sc_hd__dfxtp_1 _31216_ (.CLK(clk),
    .D(_02919_),
    .Q(\rvcpu.dp.plfd.PCD[5] ));
 sky130_fd_sc_hd__dfxtp_1 _31217_ (.CLK(clk),
    .D(_02920_),
    .Q(\rvcpu.dp.plfd.PCD[6] ));
 sky130_fd_sc_hd__dfxtp_1 _31218_ (.CLK(clk),
    .D(_02921_),
    .Q(\rvcpu.dp.plfd.PCD[7] ));
 sky130_fd_sc_hd__dfxtp_1 _31219_ (.CLK(clk),
    .D(_02922_),
    .Q(\rvcpu.dp.plfd.PCD[8] ));
 sky130_fd_sc_hd__dfxtp_1 _31220_ (.CLK(clk),
    .D(_02923_),
    .Q(\rvcpu.dp.plfd.PCD[9] ));
 sky130_fd_sc_hd__dfxtp_1 _31221_ (.CLK(clk),
    .D(_02924_),
    .Q(\rvcpu.dp.plfd.PCD[10] ));
 sky130_fd_sc_hd__dfxtp_1 _31222_ (.CLK(clk),
    .D(_02925_),
    .Q(\rvcpu.dp.plfd.PCD[11] ));
 sky130_fd_sc_hd__dfxtp_1 _31223_ (.CLK(clk),
    .D(_02926_),
    .Q(\rvcpu.dp.plfd.PCD[12] ));
 sky130_fd_sc_hd__dfxtp_1 _31224_ (.CLK(clk),
    .D(_02927_),
    .Q(\rvcpu.dp.plfd.PCD[13] ));
 sky130_fd_sc_hd__dfxtp_1 _31225_ (.CLK(clk),
    .D(_02928_),
    .Q(\rvcpu.dp.plfd.PCD[14] ));
 sky130_fd_sc_hd__dfxtp_1 _31226_ (.CLK(clk),
    .D(_02929_),
    .Q(\rvcpu.dp.plfd.PCD[15] ));
 sky130_fd_sc_hd__dfxtp_1 _31227_ (.CLK(clk),
    .D(_02930_),
    .Q(\rvcpu.dp.plfd.PCD[16] ));
 sky130_fd_sc_hd__dfxtp_1 _31228_ (.CLK(clk),
    .D(_02931_),
    .Q(\rvcpu.dp.plfd.PCD[17] ));
 sky130_fd_sc_hd__dfxtp_1 _31229_ (.CLK(clk),
    .D(_02932_),
    .Q(\rvcpu.dp.plfd.PCD[18] ));
 sky130_fd_sc_hd__dfxtp_1 _31230_ (.CLK(clk),
    .D(_02933_),
    .Q(\rvcpu.dp.plfd.PCD[19] ));
 sky130_fd_sc_hd__dfxtp_1 _31231_ (.CLK(clk),
    .D(_02934_),
    .Q(\rvcpu.dp.plfd.PCD[20] ));
 sky130_fd_sc_hd__dfxtp_1 _31232_ (.CLK(clk),
    .D(_02935_),
    .Q(\rvcpu.dp.plfd.PCD[21] ));
 sky130_fd_sc_hd__dfxtp_1 _31233_ (.CLK(clk),
    .D(_02936_),
    .Q(\rvcpu.dp.plfd.PCD[22] ));
 sky130_fd_sc_hd__dfxtp_1 _31234_ (.CLK(clk),
    .D(_02937_),
    .Q(\rvcpu.dp.plfd.PCD[23] ));
 sky130_fd_sc_hd__dfxtp_1 _31235_ (.CLK(clk),
    .D(_02938_),
    .Q(\rvcpu.dp.plfd.PCD[24] ));
 sky130_fd_sc_hd__dfxtp_1 _31236_ (.CLK(clk),
    .D(_02939_),
    .Q(\rvcpu.dp.plfd.PCD[25] ));
 sky130_fd_sc_hd__dfxtp_1 _31237_ (.CLK(clk),
    .D(_02940_),
    .Q(\rvcpu.dp.plfd.PCD[26] ));
 sky130_fd_sc_hd__dfxtp_1 _31238_ (.CLK(clk),
    .D(_02941_),
    .Q(\rvcpu.dp.plfd.PCD[27] ));
 sky130_fd_sc_hd__dfxtp_1 _31239_ (.CLK(clk),
    .D(_02942_),
    .Q(\rvcpu.dp.plfd.PCD[28] ));
 sky130_fd_sc_hd__dfxtp_1 _31240_ (.CLK(clk),
    .D(_02943_),
    .Q(\rvcpu.dp.plfd.PCD[29] ));
 sky130_fd_sc_hd__dfxtp_1 _31241_ (.CLK(clk),
    .D(_02944_),
    .Q(\rvcpu.dp.plfd.PCD[30] ));
 sky130_fd_sc_hd__dfxtp_1 _31242_ (.CLK(clk),
    .D(_02945_),
    .Q(\rvcpu.dp.plfd.PCD[31] ));
 sky130_fd_sc_hd__dfxtp_1 _31243_ (.CLK(clk),
    .D(_02946_),
    .Q(\rvcpu.dp.plfd.InstrD[0] ));
 sky130_fd_sc_hd__dfxtp_1 _31244_ (.CLK(clk),
    .D(_02947_),
    .Q(\rvcpu.dp.plfd.InstrD[2] ));
 sky130_fd_sc_hd__dfxtp_1 _31245_ (.CLK(clk),
    .D(_02948_),
    .Q(\rvcpu.dp.plfd.InstrD[3] ));
 sky130_fd_sc_hd__dfxtp_1 _31246_ (.CLK(clk),
    .D(_02949_),
    .Q(\rvcpu.dp.plfd.InstrD[4] ));
 sky130_fd_sc_hd__dfxtp_2 _31247_ (.CLK(clk),
    .D(_02950_),
    .Q(\rvcpu.c.ad.opb5 ));
 sky130_fd_sc_hd__dfxtp_2 _31248_ (.CLK(clk),
    .D(_02951_),
    .Q(\rvcpu.dp.plfd.InstrD[6] ));
 sky130_fd_sc_hd__dfxtp_1 _31249_ (.CLK(clk),
    .D(_02952_),
    .Q(\rvcpu.dp.plfd.InstrD[7] ));
 sky130_fd_sc_hd__dfxtp_1 _31250_ (.CLK(clk),
    .D(_02953_),
    .Q(\rvcpu.dp.plfd.InstrD[8] ));
 sky130_fd_sc_hd__dfxtp_1 _31251_ (.CLK(clk),
    .D(_02954_),
    .Q(\rvcpu.dp.plfd.InstrD[9] ));
 sky130_fd_sc_hd__dfxtp_1 _31252_ (.CLK(clk),
    .D(_02955_),
    .Q(\rvcpu.dp.plfd.InstrD[10] ));
 sky130_fd_sc_hd__dfxtp_1 _31253_ (.CLK(clk),
    .D(_02956_),
    .Q(\rvcpu.dp.plfd.InstrD[11] ));
 sky130_fd_sc_hd__dfxtp_1 _31254_ (.CLK(clk),
    .D(_02957_),
    .Q(\rvcpu.dp.plfd.InstrD[12] ));
 sky130_fd_sc_hd__dfxtp_1 _31255_ (.CLK(clk),
    .D(_02958_),
    .Q(\rvcpu.dp.plfd.InstrD[13] ));
 sky130_fd_sc_hd__dfxtp_2 _31256_ (.CLK(clk),
    .D(_02959_),
    .Q(\rvcpu.dp.plfd.InstrD[14] ));
 sky130_fd_sc_hd__dfxtp_4 _31257_ (.CLK(clk),
    .D(_02960_),
    .Q(\rvcpu.dp.plfd.InstrD[15] ));
 sky130_fd_sc_hd__dfxtp_4 _31258_ (.CLK(clk),
    .D(_02961_),
    .Q(\rvcpu.dp.plfd.InstrD[16] ));
 sky130_fd_sc_hd__dfxtp_4 _31259_ (.CLK(clk),
    .D(_02962_),
    .Q(\rvcpu.dp.plfd.InstrD[17] ));
 sky130_fd_sc_hd__dfxtp_2 _31260_ (.CLK(clk),
    .D(_02963_),
    .Q(\rvcpu.dp.plfd.InstrD[18] ));
 sky130_fd_sc_hd__dfxtp_4 _31261_ (.CLK(clk),
    .D(_02964_),
    .Q(\rvcpu.dp.plfd.InstrD[19] ));
 sky130_fd_sc_hd__dfxtp_1 _31262_ (.CLK(clk),
    .D(_02965_),
    .Q(\rvcpu.dp.plfd.InstrD[20] ));
 sky130_fd_sc_hd__dfxtp_1 _31263_ (.CLK(clk),
    .D(_02966_),
    .Q(\rvcpu.dp.plfd.InstrD[21] ));
 sky130_fd_sc_hd__dfxtp_2 _31264_ (.CLK(clk),
    .D(_02967_),
    .Q(\rvcpu.dp.plfd.InstrD[22] ));
 sky130_fd_sc_hd__dfxtp_2 _31265_ (.CLK(clk),
    .D(_02968_),
    .Q(\rvcpu.dp.plfd.InstrD[23] ));
 sky130_fd_sc_hd__dfxtp_4 _31266_ (.CLK(clk),
    .D(_02969_),
    .Q(\rvcpu.dp.plfd.InstrD[24] ));
 sky130_fd_sc_hd__dfxtp_1 _31267_ (.CLK(clk),
    .D(_02970_),
    .Q(\rvcpu.dp.plfd.InstrD[25] ));
 sky130_fd_sc_hd__dfxtp_1 _31268_ (.CLK(clk),
    .D(_02971_),
    .Q(\rvcpu.dp.plfd.InstrD[26] ));
 sky130_fd_sc_hd__dfxtp_1 _31269_ (.CLK(clk),
    .D(_02972_),
    .Q(\rvcpu.dp.plfd.InstrD[27] ));
 sky130_fd_sc_hd__dfxtp_1 _31270_ (.CLK(clk),
    .D(_02973_),
    .Q(\rvcpu.dp.plfd.InstrD[28] ));
 sky130_fd_sc_hd__dfxtp_1 _31271_ (.CLK(clk),
    .D(_02974_),
    .Q(\rvcpu.dp.plfd.InstrD[29] ));
 sky130_fd_sc_hd__dfxtp_1 _31272_ (.CLK(clk),
    .D(_02975_),
    .Q(\rvcpu.c.ad.funct7b5 ));
 sky130_fd_sc_hd__dfxtp_1 _31273_ (.CLK(clk),
    .D(_02976_),
    .Q(\rvcpu.dp.plfd.InstrD[31] ));
 sky130_fd_sc_hd__dfxtp_1 _31274_ (.CLK(clk),
    .D(_02977_),
    .Q(\datamem.data_ram[24][0] ));
 sky130_fd_sc_hd__dfxtp_1 _31275_ (.CLK(clk),
    .D(_02978_),
    .Q(\datamem.data_ram[24][1] ));
 sky130_fd_sc_hd__dfxtp_1 _31276_ (.CLK(clk),
    .D(_02979_),
    .Q(\datamem.data_ram[24][2] ));
 sky130_fd_sc_hd__dfxtp_1 _31277_ (.CLK(clk),
    .D(_02980_),
    .Q(\datamem.data_ram[24][3] ));
 sky130_fd_sc_hd__dfxtp_1 _31278_ (.CLK(clk),
    .D(_02981_),
    .Q(\datamem.data_ram[24][4] ));
 sky130_fd_sc_hd__dfxtp_1 _31279_ (.CLK(clk),
    .D(_02982_),
    .Q(\datamem.data_ram[24][5] ));
 sky130_fd_sc_hd__dfxtp_1 _31280_ (.CLK(clk),
    .D(_02983_),
    .Q(\datamem.data_ram[24][6] ));
 sky130_fd_sc_hd__dfxtp_1 _31281_ (.CLK(clk),
    .D(_02984_),
    .Q(\datamem.data_ram[24][7] ));
 sky130_fd_sc_hd__dfxtp_1 _31282_ (.CLK(clk),
    .D(_02985_),
    .Q(\datamem.data_ram[34][0] ));
 sky130_fd_sc_hd__dfxtp_1 _31283_ (.CLK(clk),
    .D(_02986_),
    .Q(\datamem.data_ram[34][1] ));
 sky130_fd_sc_hd__dfxtp_1 _31284_ (.CLK(clk),
    .D(_02987_),
    .Q(\datamem.data_ram[34][2] ));
 sky130_fd_sc_hd__dfxtp_1 _31285_ (.CLK(clk),
    .D(_02988_),
    .Q(\datamem.data_ram[34][3] ));
 sky130_fd_sc_hd__dfxtp_1 _31286_ (.CLK(clk),
    .D(_02989_),
    .Q(\datamem.data_ram[34][4] ));
 sky130_fd_sc_hd__dfxtp_1 _31287_ (.CLK(clk),
    .D(_02990_),
    .Q(\datamem.data_ram[34][5] ));
 sky130_fd_sc_hd__dfxtp_1 _31288_ (.CLK(clk),
    .D(_02991_),
    .Q(\datamem.data_ram[34][6] ));
 sky130_fd_sc_hd__dfxtp_1 _31289_ (.CLK(clk),
    .D(_02992_),
    .Q(\datamem.data_ram[34][7] ));
 sky130_fd_sc_hd__dfxtp_1 _31290_ (.CLK(clk),
    .D(_02993_),
    .Q(\rvcpu.dp.plde.MemWriteE ));
 sky130_fd_sc_hd__dfxtp_1 _31291_ (.CLK(clk),
    .D(_02994_),
    .Q(\rvcpu.dp.plde.unsignE ));
 sky130_fd_sc_hd__dfxtp_2 _31292_ (.CLK(clk),
    .D(_02995_),
    .Q(\rvcpu.dp.plde.JalrE ));
 sky130_fd_sc_hd__dfxtp_1 _31293_ (.CLK(clk),
    .D(_02996_),
    .Q(\rvcpu.dp.plde.JumpE ));
 sky130_fd_sc_hd__dfxtp_1 _31294_ (.CLK(clk),
    .D(_02997_),
    .Q(\rvcpu.dp.plde.BranchE ));
 sky130_fd_sc_hd__dfxtp_1 _31295_ (.CLK(clk),
    .D(_02998_),
    .Q(\rvcpu.dp.plde.RegWriteE ));
 sky130_fd_sc_hd__dfxtp_1 _31296_ (.CLK(clk),
    .D(_02999_),
    .Q(\rvcpu.dp.plde.PCPlus4E[2] ));
 sky130_fd_sc_hd__dfxtp_1 _31297_ (.CLK(clk),
    .D(_03000_),
    .Q(\rvcpu.dp.plde.PCPlus4E[3] ));
 sky130_fd_sc_hd__dfxtp_1 _31298_ (.CLK(clk),
    .D(_03001_),
    .Q(\rvcpu.dp.plde.PCPlus4E[4] ));
 sky130_fd_sc_hd__dfxtp_1 _31299_ (.CLK(clk),
    .D(_03002_),
    .Q(\rvcpu.dp.plde.PCPlus4E[5] ));
 sky130_fd_sc_hd__dfxtp_1 _31300_ (.CLK(clk),
    .D(_03003_),
    .Q(\rvcpu.dp.plde.PCPlus4E[6] ));
 sky130_fd_sc_hd__dfxtp_1 _31301_ (.CLK(clk),
    .D(_03004_),
    .Q(\rvcpu.dp.plde.PCPlus4E[7] ));
 sky130_fd_sc_hd__dfxtp_1 _31302_ (.CLK(clk),
    .D(_03005_),
    .Q(\rvcpu.dp.plde.PCPlus4E[8] ));
 sky130_fd_sc_hd__dfxtp_1 _31303_ (.CLK(clk),
    .D(_03006_),
    .Q(\rvcpu.dp.plde.PCPlus4E[9] ));
 sky130_fd_sc_hd__dfxtp_1 _31304_ (.CLK(clk),
    .D(_03007_),
    .Q(\rvcpu.dp.plde.PCPlus4E[10] ));
 sky130_fd_sc_hd__dfxtp_1 _31305_ (.CLK(clk),
    .D(_03008_),
    .Q(\rvcpu.dp.plde.PCPlus4E[11] ));
 sky130_fd_sc_hd__dfxtp_1 _31306_ (.CLK(clk),
    .D(_03009_),
    .Q(\rvcpu.dp.plde.PCPlus4E[12] ));
 sky130_fd_sc_hd__dfxtp_1 _31307_ (.CLK(clk),
    .D(_03010_),
    .Q(\rvcpu.dp.plde.PCPlus4E[13] ));
 sky130_fd_sc_hd__dfxtp_1 _31308_ (.CLK(clk),
    .D(_03011_),
    .Q(\rvcpu.dp.plde.PCPlus4E[14] ));
 sky130_fd_sc_hd__dfxtp_1 _31309_ (.CLK(clk),
    .D(_03012_),
    .Q(\rvcpu.dp.plde.PCPlus4E[15] ));
 sky130_fd_sc_hd__dfxtp_1 _31310_ (.CLK(clk),
    .D(_03013_),
    .Q(\rvcpu.dp.plde.PCPlus4E[16] ));
 sky130_fd_sc_hd__dfxtp_1 _31311_ (.CLK(clk),
    .D(_03014_),
    .Q(\rvcpu.dp.plde.PCPlus4E[17] ));
 sky130_fd_sc_hd__dfxtp_1 _31312_ (.CLK(clk),
    .D(_03015_),
    .Q(\rvcpu.dp.plde.PCPlus4E[18] ));
 sky130_fd_sc_hd__dfxtp_1 _31313_ (.CLK(clk),
    .D(_03016_),
    .Q(\rvcpu.dp.plde.PCPlus4E[19] ));
 sky130_fd_sc_hd__dfxtp_1 _31314_ (.CLK(clk),
    .D(_03017_),
    .Q(\rvcpu.dp.plde.PCPlus4E[20] ));
 sky130_fd_sc_hd__dfxtp_1 _31315_ (.CLK(clk),
    .D(_03018_),
    .Q(\rvcpu.dp.plde.PCPlus4E[21] ));
 sky130_fd_sc_hd__dfxtp_1 _31316_ (.CLK(clk),
    .D(_03019_),
    .Q(\rvcpu.dp.plde.PCPlus4E[22] ));
 sky130_fd_sc_hd__dfxtp_1 _31317_ (.CLK(clk),
    .D(_03020_),
    .Q(\rvcpu.dp.plde.PCPlus4E[23] ));
 sky130_fd_sc_hd__dfxtp_1 _31318_ (.CLK(clk),
    .D(_03021_),
    .Q(\rvcpu.dp.plde.PCPlus4E[24] ));
 sky130_fd_sc_hd__dfxtp_1 _31319_ (.CLK(clk),
    .D(_03022_),
    .Q(\rvcpu.dp.plde.PCPlus4E[25] ));
 sky130_fd_sc_hd__dfxtp_1 _31320_ (.CLK(clk),
    .D(_03023_),
    .Q(\rvcpu.dp.plde.PCPlus4E[26] ));
 sky130_fd_sc_hd__dfxtp_1 _31321_ (.CLK(clk),
    .D(_03024_),
    .Q(\rvcpu.dp.plde.PCPlus4E[27] ));
 sky130_fd_sc_hd__dfxtp_1 _31322_ (.CLK(clk),
    .D(_03025_),
    .Q(\rvcpu.dp.plde.PCPlus4E[28] ));
 sky130_fd_sc_hd__dfxtp_1 _31323_ (.CLK(clk),
    .D(_03026_),
    .Q(\rvcpu.dp.plde.PCPlus4E[29] ));
 sky130_fd_sc_hd__dfxtp_1 _31324_ (.CLK(clk),
    .D(_03027_),
    .Q(\rvcpu.dp.plde.PCPlus4E[30] ));
 sky130_fd_sc_hd__dfxtp_1 _31325_ (.CLK(clk),
    .D(_03028_),
    .Q(\rvcpu.dp.plde.PCPlus4E[31] ));
 sky130_fd_sc_hd__dfxtp_2 _31326_ (.CLK(clk),
    .D(_03029_),
    .Q(\rvcpu.dp.plde.funct3E[0] ));
 sky130_fd_sc_hd__dfxtp_2 _31327_ (.CLK(clk),
    .D(_03030_),
    .Q(\rvcpu.dp.plde.funct3E[1] ));
 sky130_fd_sc_hd__dfxtp_2 _31328_ (.CLK(clk),
    .D(_03031_),
    .Q(\rvcpu.dp.plde.funct3E[2] ));
 sky130_fd_sc_hd__dfxtp_1 _31329_ (.CLK(clk),
    .D(_03032_),
    .Q(\rvcpu.dp.plde.RdE[0] ));
 sky130_fd_sc_hd__dfxtp_1 _31330_ (.CLK(clk),
    .D(_03033_),
    .Q(\rvcpu.dp.plde.RdE[1] ));
 sky130_fd_sc_hd__dfxtp_1 _31331_ (.CLK(clk),
    .D(_03034_),
    .Q(\rvcpu.dp.plde.RdE[2] ));
 sky130_fd_sc_hd__dfxtp_1 _31332_ (.CLK(clk),
    .D(_03035_),
    .Q(\rvcpu.dp.plde.RdE[3] ));
 sky130_fd_sc_hd__dfxtp_1 _31333_ (.CLK(clk),
    .D(_03036_),
    .Q(\rvcpu.dp.plde.RdE[4] ));
 sky130_fd_sc_hd__dfxtp_1 _31334_ (.CLK(clk),
    .D(_03037_),
    .Q(\rvcpu.dp.plde.Rs2E[0] ));
 sky130_fd_sc_hd__dfxtp_1 _31335_ (.CLK(clk),
    .D(_03038_),
    .Q(\rvcpu.dp.plde.Rs2E[1] ));
 sky130_fd_sc_hd__dfxtp_1 _31336_ (.CLK(clk),
    .D(_03039_),
    .Q(\rvcpu.dp.plde.Rs2E[2] ));
 sky130_fd_sc_hd__dfxtp_1 _31337_ (.CLK(clk),
    .D(_03040_),
    .Q(\rvcpu.dp.plde.Rs2E[3] ));
 sky130_fd_sc_hd__dfxtp_1 _31338_ (.CLK(clk),
    .D(_03041_),
    .Q(\rvcpu.dp.plde.Rs2E[4] ));
 sky130_fd_sc_hd__dfxtp_1 _31339_ (.CLK(clk),
    .D(_03042_),
    .Q(\rvcpu.dp.plde.Rs1E[0] ));
 sky130_fd_sc_hd__dfxtp_1 _31340_ (.CLK(clk),
    .D(_03043_),
    .Q(\rvcpu.dp.plde.Rs1E[1] ));
 sky130_fd_sc_hd__dfxtp_1 _31341_ (.CLK(clk),
    .D(_03044_),
    .Q(\rvcpu.dp.plde.Rs1E[2] ));
 sky130_fd_sc_hd__dfxtp_1 _31342_ (.CLK(clk),
    .D(_03045_),
    .Q(\rvcpu.dp.plde.Rs1E[3] ));
 sky130_fd_sc_hd__dfxtp_1 _31343_ (.CLK(clk),
    .D(_03046_),
    .Q(\rvcpu.dp.plde.Rs1E[4] ));
 sky130_fd_sc_hd__dfxtp_2 _31344_ (.CLK(clk),
    .D(_03047_),
    .Q(\rvcpu.dp.plde.ALUControlE[0] ));
 sky130_fd_sc_hd__dfxtp_2 _31345_ (.CLK(clk),
    .D(_03048_),
    .Q(\rvcpu.dp.plde.ALUControlE[1] ));
 sky130_fd_sc_hd__dfxtp_1 _31346_ (.CLK(clk),
    .D(_03049_),
    .Q(\rvcpu.dp.plde.ALUControlE[2] ));
 sky130_fd_sc_hd__dfxtp_1 _31347_ (.CLK(clk),
    .D(_03050_),
    .Q(\rvcpu.dp.plde.ALUControlE[3] ));
 sky130_fd_sc_hd__dfxtp_2 _31348_ (.CLK(clk),
    .D(_03051_),
    .Q(\rvcpu.dp.plde.luiE ));
 sky130_fd_sc_hd__dfxtp_1 _31349_ (.CLK(clk),
    .D(_03052_),
    .Q(\rvcpu.dp.hu.ResultSrcE0 ));
 sky130_fd_sc_hd__dfxtp_1 _31350_ (.CLK(clk),
    .D(_03053_),
    .Q(\rvcpu.dp.plde.ResultSrcE[1] ));
 sky130_fd_sc_hd__dfxtp_4 _31351_ (.CLK(clk),
    .D(_03054_),
    .Q(\rvcpu.dp.plde.ImmExtE[0] ));
 sky130_fd_sc_hd__dfxtp_4 _31352_ (.CLK(clk),
    .D(_03055_),
    .Q(\rvcpu.dp.plde.ImmExtE[1] ));
 sky130_fd_sc_hd__dfxtp_2 _31353_ (.CLK(clk),
    .D(_03056_),
    .Q(\rvcpu.dp.plde.ImmExtE[2] ));
 sky130_fd_sc_hd__dfxtp_2 _31354_ (.CLK(clk),
    .D(_03057_),
    .Q(\rvcpu.dp.plde.ImmExtE[3] ));
 sky130_fd_sc_hd__dfxtp_4 _31355_ (.CLK(clk),
    .D(_03058_),
    .Q(\rvcpu.dp.plde.ImmExtE[4] ));
 sky130_fd_sc_hd__dfxtp_2 _31356_ (.CLK(clk),
    .D(_03059_),
    .Q(\rvcpu.dp.plde.ImmExtE[5] ));
 sky130_fd_sc_hd__dfxtp_2 _31357_ (.CLK(clk),
    .D(_03060_),
    .Q(\rvcpu.dp.plde.ImmExtE[6] ));
 sky130_fd_sc_hd__dfxtp_2 _31358_ (.CLK(clk),
    .D(_03061_),
    .Q(\rvcpu.dp.plde.ImmExtE[7] ));
 sky130_fd_sc_hd__dfxtp_2 _31359_ (.CLK(clk),
    .D(_03062_),
    .Q(\rvcpu.dp.plde.ImmExtE[8] ));
 sky130_fd_sc_hd__dfxtp_4 _31360_ (.CLK(clk),
    .D(_03063_),
    .Q(\rvcpu.dp.plde.ImmExtE[9] ));
 sky130_fd_sc_hd__dfxtp_2 _31361_ (.CLK(clk),
    .D(_03064_),
    .Q(\rvcpu.dp.plde.ImmExtE[10] ));
 sky130_fd_sc_hd__dfxtp_2 _31362_ (.CLK(clk),
    .D(_03065_),
    .Q(\rvcpu.dp.plde.ImmExtE[11] ));
 sky130_fd_sc_hd__dfxtp_2 _31363_ (.CLK(clk),
    .D(_03066_),
    .Q(\rvcpu.dp.plde.ImmExtE[12] ));
 sky130_fd_sc_hd__dfxtp_2 _31364_ (.CLK(clk),
    .D(_03067_),
    .Q(\rvcpu.dp.plde.ImmExtE[13] ));
 sky130_fd_sc_hd__dfxtp_2 _31365_ (.CLK(clk),
    .D(_03068_),
    .Q(\rvcpu.dp.plde.ImmExtE[14] ));
 sky130_fd_sc_hd__dfxtp_2 _31366_ (.CLK(clk),
    .D(_03069_),
    .Q(\rvcpu.dp.plde.ImmExtE[15] ));
 sky130_fd_sc_hd__dfxtp_2 _31367_ (.CLK(clk),
    .D(_03070_),
    .Q(\rvcpu.dp.plde.ImmExtE[16] ));
 sky130_fd_sc_hd__dfxtp_2 _31368_ (.CLK(clk),
    .D(_03071_),
    .Q(\rvcpu.dp.plde.ImmExtE[17] ));
 sky130_fd_sc_hd__dfxtp_2 _31369_ (.CLK(clk),
    .D(_03072_),
    .Q(\rvcpu.dp.plde.ImmExtE[18] ));
 sky130_fd_sc_hd__dfxtp_2 _31370_ (.CLK(clk),
    .D(_03073_),
    .Q(\rvcpu.dp.plde.ImmExtE[19] ));
 sky130_fd_sc_hd__dfxtp_1 _31371_ (.CLK(clk),
    .D(_03074_),
    .Q(\rvcpu.dp.plde.ImmExtE[20] ));
 sky130_fd_sc_hd__dfxtp_1 _31372_ (.CLK(clk),
    .D(_03075_),
    .Q(\rvcpu.dp.plde.ImmExtE[21] ));
 sky130_fd_sc_hd__dfxtp_1 _31373_ (.CLK(clk),
    .D(_03076_),
    .Q(\rvcpu.dp.plde.ImmExtE[22] ));
 sky130_fd_sc_hd__dfxtp_1 _31374_ (.CLK(clk),
    .D(_03077_),
    .Q(\rvcpu.dp.plde.ImmExtE[23] ));
 sky130_fd_sc_hd__dfxtp_1 _31375_ (.CLK(clk),
    .D(_03078_),
    .Q(\rvcpu.dp.plde.ImmExtE[24] ));
 sky130_fd_sc_hd__dfxtp_1 _31376_ (.CLK(clk),
    .D(_03079_),
    .Q(\rvcpu.dp.plde.ImmExtE[25] ));
 sky130_fd_sc_hd__dfxtp_2 _31377_ (.CLK(clk),
    .D(_03080_),
    .Q(\rvcpu.dp.plde.ImmExtE[26] ));
 sky130_fd_sc_hd__dfxtp_1 _31378_ (.CLK(clk),
    .D(_03081_),
    .Q(\rvcpu.dp.plde.ImmExtE[27] ));
 sky130_fd_sc_hd__dfxtp_1 _31379_ (.CLK(clk),
    .D(_03082_),
    .Q(\rvcpu.dp.plde.ImmExtE[28] ));
 sky130_fd_sc_hd__dfxtp_1 _31380_ (.CLK(clk),
    .D(_03083_),
    .Q(\rvcpu.dp.plde.ImmExtE[29] ));
 sky130_fd_sc_hd__dfxtp_1 _31381_ (.CLK(clk),
    .D(_03084_),
    .Q(\rvcpu.dp.plde.ImmExtE[30] ));
 sky130_fd_sc_hd__dfxtp_1 _31382_ (.CLK(clk),
    .D(_03085_),
    .Q(\rvcpu.dp.plde.ImmExtE[31] ));
 sky130_fd_sc_hd__dfxtp_1 _31383_ (.CLK(clk),
    .D(_03086_),
    .Q(\rvcpu.dp.plde.PCE[0] ));
 sky130_fd_sc_hd__dfxtp_1 _31384_ (.CLK(clk),
    .D(_03087_),
    .Q(\rvcpu.dp.plde.PCE[1] ));
 sky130_fd_sc_hd__dfxtp_1 _31385_ (.CLK(clk),
    .D(_03088_),
    .Q(\rvcpu.dp.plde.PCE[2] ));
 sky130_fd_sc_hd__dfxtp_1 _31386_ (.CLK(clk),
    .D(_03089_),
    .Q(\rvcpu.dp.plde.PCE[3] ));
 sky130_fd_sc_hd__dfxtp_1 _31387_ (.CLK(clk),
    .D(_03090_),
    .Q(\rvcpu.dp.plde.PCE[4] ));
 sky130_fd_sc_hd__dfxtp_1 _31388_ (.CLK(clk),
    .D(_03091_),
    .Q(\rvcpu.dp.plde.PCE[5] ));
 sky130_fd_sc_hd__dfxtp_1 _31389_ (.CLK(clk),
    .D(_03092_),
    .Q(\rvcpu.dp.plde.PCE[6] ));
 sky130_fd_sc_hd__dfxtp_1 _31390_ (.CLK(clk),
    .D(_03093_),
    .Q(\rvcpu.dp.plde.PCE[7] ));
 sky130_fd_sc_hd__dfxtp_1 _31391_ (.CLK(clk),
    .D(_03094_),
    .Q(\rvcpu.dp.plde.PCE[8] ));
 sky130_fd_sc_hd__dfxtp_1 _31392_ (.CLK(clk),
    .D(_03095_),
    .Q(\rvcpu.dp.plde.PCE[9] ));
 sky130_fd_sc_hd__dfxtp_1 _31393_ (.CLK(clk),
    .D(_03096_),
    .Q(\rvcpu.dp.plde.PCE[10] ));
 sky130_fd_sc_hd__dfxtp_1 _31394_ (.CLK(clk),
    .D(_03097_),
    .Q(\rvcpu.dp.plde.PCE[11] ));
 sky130_fd_sc_hd__dfxtp_1 _31395_ (.CLK(clk),
    .D(_03098_),
    .Q(\rvcpu.dp.plde.PCE[12] ));
 sky130_fd_sc_hd__dfxtp_1 _31396_ (.CLK(clk),
    .D(_03099_),
    .Q(\rvcpu.dp.plde.PCE[13] ));
 sky130_fd_sc_hd__dfxtp_1 _31397_ (.CLK(clk),
    .D(_03100_),
    .Q(\rvcpu.dp.plde.PCE[14] ));
 sky130_fd_sc_hd__dfxtp_1 _31398_ (.CLK(clk),
    .D(_03101_),
    .Q(\rvcpu.dp.plde.PCE[15] ));
 sky130_fd_sc_hd__dfxtp_1 _31399_ (.CLK(clk),
    .D(_03102_),
    .Q(\rvcpu.dp.plde.PCE[16] ));
 sky130_fd_sc_hd__dfxtp_1 _31400_ (.CLK(clk),
    .D(_03103_),
    .Q(\rvcpu.dp.plde.PCE[17] ));
 sky130_fd_sc_hd__dfxtp_1 _31401_ (.CLK(clk),
    .D(_03104_),
    .Q(\rvcpu.dp.plde.PCE[18] ));
 sky130_fd_sc_hd__dfxtp_1 _31402_ (.CLK(clk),
    .D(_03105_),
    .Q(\rvcpu.dp.plde.PCE[19] ));
 sky130_fd_sc_hd__dfxtp_1 _31403_ (.CLK(clk),
    .D(_03106_),
    .Q(\rvcpu.dp.plde.PCE[20] ));
 sky130_fd_sc_hd__dfxtp_1 _31404_ (.CLK(clk),
    .D(_03107_),
    .Q(\rvcpu.dp.plde.PCE[21] ));
 sky130_fd_sc_hd__dfxtp_1 _31405_ (.CLK(clk),
    .D(_03108_),
    .Q(\rvcpu.dp.plde.PCE[22] ));
 sky130_fd_sc_hd__dfxtp_1 _31406_ (.CLK(clk),
    .D(_03109_),
    .Q(\rvcpu.dp.plde.PCE[23] ));
 sky130_fd_sc_hd__dfxtp_1 _31407_ (.CLK(clk),
    .D(_03110_),
    .Q(\rvcpu.dp.plde.PCE[24] ));
 sky130_fd_sc_hd__dfxtp_1 _31408_ (.CLK(clk),
    .D(_03111_),
    .Q(\rvcpu.dp.plde.PCE[25] ));
 sky130_fd_sc_hd__dfxtp_1 _31409_ (.CLK(clk),
    .D(_03112_),
    .Q(\rvcpu.dp.plde.PCE[26] ));
 sky130_fd_sc_hd__dfxtp_1 _31410_ (.CLK(clk),
    .D(_03113_),
    .Q(\rvcpu.dp.plde.PCE[27] ));
 sky130_fd_sc_hd__dfxtp_1 _31411_ (.CLK(clk),
    .D(_03114_),
    .Q(\rvcpu.dp.plde.PCE[28] ));
 sky130_fd_sc_hd__dfxtp_1 _31412_ (.CLK(clk),
    .D(_03115_),
    .Q(\rvcpu.dp.plde.PCE[29] ));
 sky130_fd_sc_hd__dfxtp_1 _31413_ (.CLK(clk),
    .D(_03116_),
    .Q(\rvcpu.dp.plde.PCE[30] ));
 sky130_fd_sc_hd__dfxtp_1 _31414_ (.CLK(clk),
    .D(_03117_),
    .Q(\rvcpu.dp.plde.PCE[31] ));
 sky130_fd_sc_hd__dfxtp_1 _31415_ (.CLK(clk),
    .D(_03118_),
    .Q(\datamem.data_ram[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _31416_ (.CLK(clk),
    .D(_03119_),
    .Q(\datamem.data_ram[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _31417_ (.CLK(clk),
    .D(_03120_),
    .Q(\datamem.data_ram[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _31418_ (.CLK(clk),
    .D(_03121_),
    .Q(\datamem.data_ram[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _31419_ (.CLK(clk),
    .D(_03122_),
    .Q(\datamem.data_ram[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _31420_ (.CLK(clk),
    .D(_03123_),
    .Q(\datamem.data_ram[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _31421_ (.CLK(clk),
    .D(_03124_),
    .Q(\datamem.data_ram[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _31422_ (.CLK(clk),
    .D(_03125_),
    .Q(\datamem.data_ram[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _31423_ (.CLK(clk),
    .D(_03126_),
    .Q(\datamem.data_ram[44][0] ));
 sky130_fd_sc_hd__dfxtp_1 _31424_ (.CLK(clk),
    .D(_03127_),
    .Q(\datamem.data_ram[44][1] ));
 sky130_fd_sc_hd__dfxtp_1 _31425_ (.CLK(clk),
    .D(_03128_),
    .Q(\datamem.data_ram[44][2] ));
 sky130_fd_sc_hd__dfxtp_1 _31426_ (.CLK(clk),
    .D(_03129_),
    .Q(\datamem.data_ram[44][3] ));
 sky130_fd_sc_hd__dfxtp_1 _31427_ (.CLK(clk),
    .D(_03130_),
    .Q(\datamem.data_ram[44][4] ));
 sky130_fd_sc_hd__dfxtp_1 _31428_ (.CLK(clk),
    .D(_03131_),
    .Q(\datamem.data_ram[44][5] ));
 sky130_fd_sc_hd__dfxtp_1 _31429_ (.CLK(clk),
    .D(_03132_),
    .Q(\datamem.data_ram[44][6] ));
 sky130_fd_sc_hd__dfxtp_1 _31430_ (.CLK(clk),
    .D(_03133_),
    .Q(\datamem.data_ram[44][7] ));
 sky130_fd_sc_hd__dfxtp_1 _31431_ (.CLK(clk),
    .D(_03134_),
    .Q(\datamem.data_ram[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _31432_ (.CLK(clk),
    .D(_03135_),
    .Q(\datamem.data_ram[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _31433_ (.CLK(clk),
    .D(_03136_),
    .Q(\datamem.data_ram[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _31434_ (.CLK(clk),
    .D(_03137_),
    .Q(\datamem.data_ram[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _31435_ (.CLK(clk),
    .D(_03138_),
    .Q(\datamem.data_ram[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _31436_ (.CLK(clk),
    .D(_03139_),
    .Q(\datamem.data_ram[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _31437_ (.CLK(clk),
    .D(_03140_),
    .Q(\datamem.data_ram[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _31438_ (.CLK(clk),
    .D(_03141_),
    .Q(\datamem.data_ram[14][7] ));
 sky130_fd_sc_hd__dlxtn_1 _31439_ (.D(_00002_),
    .GATE_N(_00003_),
    .Q(\rvcpu.dp.Cout ));
 sky130_fd_sc_hd__dfxtp_1 _31440_ (.CLK(clk),
    .D(\rvcpu.dp.hu.ResultSrcE0 ),
    .Q(\rvcpu.dp.plem.ResultSrcM[0] ));
 sky130_fd_sc_hd__dfxtp_1 _31441_ (.CLK(clk),
    .D(\rvcpu.dp.plde.ResultSrcE[1] ),
    .Q(\rvcpu.dp.plem.ResultSrcM[1] ));
 sky130_fd_sc_hd__dfxtp_2 _31442_ (.CLK(clk),
    .D(\rvcpu.dp.SrcBFW_Mux.y[0] ),
    .Q(\rvcpu.dp.plem.WriteDataM[0] ));
 sky130_fd_sc_hd__dfxtp_2 _31443_ (.CLK(clk),
    .D(\rvcpu.dp.SrcBFW_Mux.y[1] ),
    .Q(\rvcpu.dp.plem.WriteDataM[1] ));
 sky130_fd_sc_hd__dfxtp_2 _31444_ (.CLK(clk),
    .D(\rvcpu.dp.SrcBFW_Mux.y[2] ),
    .Q(\rvcpu.dp.plem.WriteDataM[2] ));
 sky130_fd_sc_hd__dfxtp_2 _31445_ (.CLK(clk),
    .D(\rvcpu.dp.SrcBFW_Mux.y[3] ),
    .Q(\rvcpu.dp.plem.WriteDataM[3] ));
 sky130_fd_sc_hd__dfxtp_2 _31446_ (.CLK(clk),
    .D(\rvcpu.dp.SrcBFW_Mux.y[4] ),
    .Q(\rvcpu.dp.plem.WriteDataM[4] ));
 sky130_fd_sc_hd__dfxtp_2 _31447_ (.CLK(clk),
    .D(\rvcpu.dp.SrcBFW_Mux.y[5] ),
    .Q(\rvcpu.dp.plem.WriteDataM[5] ));
 sky130_fd_sc_hd__dfxtp_2 _31448_ (.CLK(clk),
    .D(\rvcpu.dp.SrcBFW_Mux.y[6] ),
    .Q(\rvcpu.dp.plem.WriteDataM[6] ));
 sky130_fd_sc_hd__dfxtp_2 _31449_ (.CLK(clk),
    .D(\rvcpu.dp.SrcBFW_Mux.y[7] ),
    .Q(\rvcpu.dp.plem.WriteDataM[7] ));
 sky130_fd_sc_hd__dfxtp_1 _31450_ (.CLK(clk),
    .D(\rvcpu.dp.SrcBFW_Mux.y[8] ),
    .Q(\rvcpu.dp.plem.WriteDataM[8] ));
 sky130_fd_sc_hd__dfxtp_1 _31451_ (.CLK(clk),
    .D(\rvcpu.dp.SrcBFW_Mux.y[9] ),
    .Q(\rvcpu.dp.plem.WriteDataM[9] ));
 sky130_fd_sc_hd__dfxtp_1 _31452_ (.CLK(clk),
    .D(\rvcpu.dp.SrcBFW_Mux.y[10] ),
    .Q(\rvcpu.dp.plem.WriteDataM[10] ));
 sky130_fd_sc_hd__dfxtp_1 _31453_ (.CLK(clk),
    .D(\rvcpu.dp.SrcBFW_Mux.y[11] ),
    .Q(\rvcpu.dp.plem.WriteDataM[11] ));
 sky130_fd_sc_hd__dfxtp_1 _31454_ (.CLK(clk),
    .D(\rvcpu.dp.SrcBFW_Mux.y[12] ),
    .Q(\rvcpu.dp.plem.WriteDataM[12] ));
 sky130_fd_sc_hd__dfxtp_1 _31455_ (.CLK(clk),
    .D(\rvcpu.dp.SrcBFW_Mux.y[13] ),
    .Q(\rvcpu.dp.plem.WriteDataM[13] ));
 sky130_fd_sc_hd__dfxtp_1 _31456_ (.CLK(clk),
    .D(\rvcpu.dp.SrcBFW_Mux.y[14] ),
    .Q(\rvcpu.dp.plem.WriteDataM[14] ));
 sky130_fd_sc_hd__dfxtp_1 _31457_ (.CLK(clk),
    .D(\rvcpu.dp.SrcBFW_Mux.y[15] ),
    .Q(\rvcpu.dp.plem.WriteDataM[15] ));
 sky130_fd_sc_hd__dfxtp_1 _31458_ (.CLK(clk),
    .D(\rvcpu.dp.SrcBFW_Mux.y[16] ),
    .Q(\rvcpu.dp.plem.WriteDataM[16] ));
 sky130_fd_sc_hd__dfxtp_1 _31459_ (.CLK(clk),
    .D(\rvcpu.dp.SrcBFW_Mux.y[17] ),
    .Q(\rvcpu.dp.plem.WriteDataM[17] ));
 sky130_fd_sc_hd__dfxtp_1 _31460_ (.CLK(clk),
    .D(\rvcpu.dp.SrcBFW_Mux.y[18] ),
    .Q(\rvcpu.dp.plem.WriteDataM[18] ));
 sky130_fd_sc_hd__dfxtp_1 _31461_ (.CLK(clk),
    .D(\rvcpu.dp.SrcBFW_Mux.y[19] ),
    .Q(\rvcpu.dp.plem.WriteDataM[19] ));
 sky130_fd_sc_hd__dfxtp_1 _31462_ (.CLK(clk),
    .D(\rvcpu.dp.SrcBFW_Mux.y[20] ),
    .Q(\rvcpu.dp.plem.WriteDataM[20] ));
 sky130_fd_sc_hd__dfxtp_1 _31463_ (.CLK(clk),
    .D(\rvcpu.dp.SrcBFW_Mux.y[21] ),
    .Q(\rvcpu.dp.plem.WriteDataM[21] ));
 sky130_fd_sc_hd__dfxtp_1 _31464_ (.CLK(clk),
    .D(\rvcpu.dp.SrcBFW_Mux.y[22] ),
    .Q(\rvcpu.dp.plem.WriteDataM[22] ));
 sky130_fd_sc_hd__dfxtp_1 _31465_ (.CLK(clk),
    .D(\rvcpu.dp.SrcBFW_Mux.y[23] ),
    .Q(\rvcpu.dp.plem.WriteDataM[23] ));
 sky130_fd_sc_hd__dfxtp_1 _31466_ (.CLK(clk),
    .D(\rvcpu.dp.SrcBFW_Mux.y[24] ),
    .Q(\rvcpu.dp.plem.WriteDataM[24] ));
 sky130_fd_sc_hd__dfxtp_1 _31467_ (.CLK(clk),
    .D(\rvcpu.dp.SrcBFW_Mux.y[25] ),
    .Q(\rvcpu.dp.plem.WriteDataM[25] ));
 sky130_fd_sc_hd__dfxtp_1 _31468_ (.CLK(clk),
    .D(\rvcpu.dp.SrcBFW_Mux.y[26] ),
    .Q(\rvcpu.dp.plem.WriteDataM[26] ));
 sky130_fd_sc_hd__dfxtp_1 _31469_ (.CLK(clk),
    .D(\rvcpu.dp.SrcBFW_Mux.y[27] ),
    .Q(\rvcpu.dp.plem.WriteDataM[27] ));
 sky130_fd_sc_hd__dfxtp_1 _31470_ (.CLK(clk),
    .D(\rvcpu.dp.SrcBFW_Mux.y[28] ),
    .Q(\rvcpu.dp.plem.WriteDataM[28] ));
 sky130_fd_sc_hd__dfxtp_1 _31471_ (.CLK(clk),
    .D(\rvcpu.dp.SrcBFW_Mux.y[29] ),
    .Q(\rvcpu.dp.plem.WriteDataM[29] ));
 sky130_fd_sc_hd__dfxtp_1 _31472_ (.CLK(clk),
    .D(\rvcpu.dp.SrcBFW_Mux.y[30] ),
    .Q(\rvcpu.dp.plem.WriteDataM[30] ));
 sky130_fd_sc_hd__dfxtp_1 _31473_ (.CLK(clk),
    .D(\rvcpu.dp.SrcBFW_Mux.y[31] ),
    .Q(\rvcpu.dp.plem.WriteDataM[31] ));
 sky130_fd_sc_hd__dfxtp_1 _31474_ (.CLK(clk),
    .D(\rvcpu.dp.lAuiPCE[0] ),
    .Q(\rvcpu.dp.plem.lAuiPCM[0] ));
 sky130_fd_sc_hd__dfxtp_1 _31475_ (.CLK(clk),
    .D(\rvcpu.dp.lAuiPCE[1] ),
    .Q(\rvcpu.dp.plem.lAuiPCM[1] ));
 sky130_fd_sc_hd__dfxtp_1 _31476_ (.CLK(clk),
    .D(\rvcpu.dp.lAuiPCE[2] ),
    .Q(\rvcpu.dp.plem.lAuiPCM[2] ));
 sky130_fd_sc_hd__dfxtp_1 _31477_ (.CLK(clk),
    .D(\rvcpu.dp.lAuiPCE[3] ),
    .Q(\rvcpu.dp.plem.lAuiPCM[3] ));
 sky130_fd_sc_hd__dfxtp_1 _31478_ (.CLK(clk),
    .D(\rvcpu.dp.lAuiPCE[4] ),
    .Q(\rvcpu.dp.plem.lAuiPCM[4] ));
 sky130_fd_sc_hd__dfxtp_1 _31479_ (.CLK(clk),
    .D(\rvcpu.dp.lAuiPCE[5] ),
    .Q(\rvcpu.dp.plem.lAuiPCM[5] ));
 sky130_fd_sc_hd__dfxtp_1 _31480_ (.CLK(clk),
    .D(\rvcpu.dp.lAuiPCE[6] ),
    .Q(\rvcpu.dp.plem.lAuiPCM[6] ));
 sky130_fd_sc_hd__dfxtp_1 _31481_ (.CLK(clk),
    .D(\rvcpu.dp.lAuiPCE[7] ),
    .Q(\rvcpu.dp.plem.lAuiPCM[7] ));
 sky130_fd_sc_hd__dfxtp_1 _31482_ (.CLK(clk),
    .D(\rvcpu.dp.lAuiPCE[8] ),
    .Q(\rvcpu.dp.plem.lAuiPCM[8] ));
 sky130_fd_sc_hd__dfxtp_1 _31483_ (.CLK(clk),
    .D(\rvcpu.dp.lAuiPCE[9] ),
    .Q(\rvcpu.dp.plem.lAuiPCM[9] ));
 sky130_fd_sc_hd__dfxtp_1 _31484_ (.CLK(clk),
    .D(\rvcpu.dp.lAuiPCE[10] ),
    .Q(\rvcpu.dp.plem.lAuiPCM[10] ));
 sky130_fd_sc_hd__dfxtp_1 _31485_ (.CLK(clk),
    .D(\rvcpu.dp.lAuiPCE[11] ),
    .Q(\rvcpu.dp.plem.lAuiPCM[11] ));
 sky130_fd_sc_hd__dfxtp_1 _31486_ (.CLK(clk),
    .D(\rvcpu.dp.lAuiPCE[12] ),
    .Q(\rvcpu.dp.plem.lAuiPCM[12] ));
 sky130_fd_sc_hd__dfxtp_1 _31487_ (.CLK(clk),
    .D(\rvcpu.dp.lAuiPCE[13] ),
    .Q(\rvcpu.dp.plem.lAuiPCM[13] ));
 sky130_fd_sc_hd__dfxtp_1 _31488_ (.CLK(clk),
    .D(\rvcpu.dp.lAuiPCE[14] ),
    .Q(\rvcpu.dp.plem.lAuiPCM[14] ));
 sky130_fd_sc_hd__dfxtp_1 _31489_ (.CLK(clk),
    .D(\rvcpu.dp.lAuiPCE[15] ),
    .Q(\rvcpu.dp.plem.lAuiPCM[15] ));
 sky130_fd_sc_hd__dfxtp_1 _31490_ (.CLK(clk),
    .D(\rvcpu.dp.lAuiPCE[16] ),
    .Q(\rvcpu.dp.plem.lAuiPCM[16] ));
 sky130_fd_sc_hd__dfxtp_1 _31491_ (.CLK(clk),
    .D(\rvcpu.dp.lAuiPCE[17] ),
    .Q(\rvcpu.dp.plem.lAuiPCM[17] ));
 sky130_fd_sc_hd__dfxtp_1 _31492_ (.CLK(clk),
    .D(\rvcpu.dp.lAuiPCE[18] ),
    .Q(\rvcpu.dp.plem.lAuiPCM[18] ));
 sky130_fd_sc_hd__dfxtp_1 _31493_ (.CLK(clk),
    .D(\rvcpu.dp.lAuiPCE[19] ),
    .Q(\rvcpu.dp.plem.lAuiPCM[19] ));
 sky130_fd_sc_hd__dfxtp_1 _31494_ (.CLK(clk),
    .D(\rvcpu.dp.lAuiPCE[20] ),
    .Q(\rvcpu.dp.plem.lAuiPCM[20] ));
 sky130_fd_sc_hd__dfxtp_1 _31495_ (.CLK(clk),
    .D(\rvcpu.dp.lAuiPCE[21] ),
    .Q(\rvcpu.dp.plem.lAuiPCM[21] ));
 sky130_fd_sc_hd__dfxtp_1 _31496_ (.CLK(clk),
    .D(\rvcpu.dp.lAuiPCE[22] ),
    .Q(\rvcpu.dp.plem.lAuiPCM[22] ));
 sky130_fd_sc_hd__dfxtp_1 _31497_ (.CLK(clk),
    .D(\rvcpu.dp.lAuiPCE[23] ),
    .Q(\rvcpu.dp.plem.lAuiPCM[23] ));
 sky130_fd_sc_hd__dfxtp_1 _31498_ (.CLK(clk),
    .D(\rvcpu.dp.lAuiPCE[24] ),
    .Q(\rvcpu.dp.plem.lAuiPCM[24] ));
 sky130_fd_sc_hd__dfxtp_1 _31499_ (.CLK(clk),
    .D(\rvcpu.dp.lAuiPCE[25] ),
    .Q(\rvcpu.dp.plem.lAuiPCM[25] ));
 sky130_fd_sc_hd__dfxtp_1 _31500_ (.CLK(clk),
    .D(\rvcpu.dp.lAuiPCE[26] ),
    .Q(\rvcpu.dp.plem.lAuiPCM[26] ));
 sky130_fd_sc_hd__dfxtp_1 _31501_ (.CLK(clk),
    .D(\rvcpu.dp.lAuiPCE[27] ),
    .Q(\rvcpu.dp.plem.lAuiPCM[27] ));
 sky130_fd_sc_hd__dfxtp_1 _31502_ (.CLK(clk),
    .D(\rvcpu.dp.lAuiPCE[28] ),
    .Q(\rvcpu.dp.plem.lAuiPCM[28] ));
 sky130_fd_sc_hd__dfxtp_1 _31503_ (.CLK(clk),
    .D(\rvcpu.dp.lAuiPCE[29] ),
    .Q(\rvcpu.dp.plem.lAuiPCM[29] ));
 sky130_fd_sc_hd__dfxtp_1 _31504_ (.CLK(clk),
    .D(\rvcpu.dp.lAuiPCE[30] ),
    .Q(\rvcpu.dp.plem.lAuiPCM[30] ));
 sky130_fd_sc_hd__dfxtp_1 _31505_ (.CLK(clk),
    .D(\rvcpu.dp.lAuiPCE[31] ),
    .Q(\rvcpu.dp.plem.lAuiPCM[31] ));
 sky130_fd_sc_hd__dfxtp_1 _31506_ (.CLK(clk),
    .D(\rvcpu.dp.plde.PCE[0] ),
    .Q(\rvcpu.dp.plem.PCPlus4M[0] ));
 sky130_fd_sc_hd__dfxtp_1 _31507_ (.CLK(clk),
    .D(\rvcpu.dp.plde.PCE[1] ),
    .Q(\rvcpu.dp.plem.PCPlus4M[1] ));
 sky130_fd_sc_hd__dfxtp_1 _31508_ (.CLK(clk),
    .D(\rvcpu.dp.plde.PCPlus4E[2] ),
    .Q(\rvcpu.dp.plem.PCPlus4M[2] ));
 sky130_fd_sc_hd__dfxtp_1 _31509_ (.CLK(clk),
    .D(\rvcpu.dp.plde.PCPlus4E[3] ),
    .Q(\rvcpu.dp.plem.PCPlus4M[3] ));
 sky130_fd_sc_hd__dfxtp_1 _31510_ (.CLK(clk),
    .D(\rvcpu.dp.plde.PCPlus4E[4] ),
    .Q(\rvcpu.dp.plem.PCPlus4M[4] ));
 sky130_fd_sc_hd__dfxtp_1 _31511_ (.CLK(clk),
    .D(\rvcpu.dp.plde.PCPlus4E[5] ),
    .Q(\rvcpu.dp.plem.PCPlus4M[5] ));
 sky130_fd_sc_hd__dfxtp_1 _31512_ (.CLK(clk),
    .D(\rvcpu.dp.plde.PCPlus4E[6] ),
    .Q(\rvcpu.dp.plem.PCPlus4M[6] ));
 sky130_fd_sc_hd__dfxtp_1 _31513_ (.CLK(clk),
    .D(\rvcpu.dp.plde.PCPlus4E[7] ),
    .Q(\rvcpu.dp.plem.PCPlus4M[7] ));
 sky130_fd_sc_hd__dfxtp_1 _31514_ (.CLK(clk),
    .D(\rvcpu.dp.plde.PCPlus4E[8] ),
    .Q(\rvcpu.dp.plem.PCPlus4M[8] ));
 sky130_fd_sc_hd__dfxtp_1 _31515_ (.CLK(clk),
    .D(\rvcpu.dp.plde.PCPlus4E[9] ),
    .Q(\rvcpu.dp.plem.PCPlus4M[9] ));
 sky130_fd_sc_hd__dfxtp_1 _31516_ (.CLK(clk),
    .D(\rvcpu.dp.plde.PCPlus4E[10] ),
    .Q(\rvcpu.dp.plem.PCPlus4M[10] ));
 sky130_fd_sc_hd__dfxtp_1 _31517_ (.CLK(clk),
    .D(\rvcpu.dp.plde.PCPlus4E[11] ),
    .Q(\rvcpu.dp.plem.PCPlus4M[11] ));
 sky130_fd_sc_hd__dfxtp_1 _31518_ (.CLK(clk),
    .D(\rvcpu.dp.plde.PCPlus4E[12] ),
    .Q(\rvcpu.dp.plem.PCPlus4M[12] ));
 sky130_fd_sc_hd__dfxtp_1 _31519_ (.CLK(clk),
    .D(\rvcpu.dp.plde.PCPlus4E[13] ),
    .Q(\rvcpu.dp.plem.PCPlus4M[13] ));
 sky130_fd_sc_hd__dfxtp_1 _31520_ (.CLK(clk),
    .D(\rvcpu.dp.plde.PCPlus4E[14] ),
    .Q(\rvcpu.dp.plem.PCPlus4M[14] ));
 sky130_fd_sc_hd__dfxtp_1 _31521_ (.CLK(clk),
    .D(\rvcpu.dp.plde.PCPlus4E[15] ),
    .Q(\rvcpu.dp.plem.PCPlus4M[15] ));
 sky130_fd_sc_hd__dfxtp_1 _31522_ (.CLK(clk),
    .D(\rvcpu.dp.plde.PCPlus4E[16] ),
    .Q(\rvcpu.dp.plem.PCPlus4M[16] ));
 sky130_fd_sc_hd__dfxtp_1 _31523_ (.CLK(clk),
    .D(\rvcpu.dp.plde.PCPlus4E[17] ),
    .Q(\rvcpu.dp.plem.PCPlus4M[17] ));
 sky130_fd_sc_hd__dfxtp_1 _31524_ (.CLK(clk),
    .D(\rvcpu.dp.plde.PCPlus4E[18] ),
    .Q(\rvcpu.dp.plem.PCPlus4M[18] ));
 sky130_fd_sc_hd__dfxtp_1 _31525_ (.CLK(clk),
    .D(\rvcpu.dp.plde.PCPlus4E[19] ),
    .Q(\rvcpu.dp.plem.PCPlus4M[19] ));
 sky130_fd_sc_hd__dfxtp_1 _31526_ (.CLK(clk),
    .D(\rvcpu.dp.plde.PCPlus4E[20] ),
    .Q(\rvcpu.dp.plem.PCPlus4M[20] ));
 sky130_fd_sc_hd__dfxtp_1 _31527_ (.CLK(clk),
    .D(\rvcpu.dp.plde.PCPlus4E[21] ),
    .Q(\rvcpu.dp.plem.PCPlus4M[21] ));
 sky130_fd_sc_hd__dfxtp_1 _31528_ (.CLK(clk),
    .D(\rvcpu.dp.plde.PCPlus4E[22] ),
    .Q(\rvcpu.dp.plem.PCPlus4M[22] ));
 sky130_fd_sc_hd__dfxtp_1 _31529_ (.CLK(clk),
    .D(\rvcpu.dp.plde.PCPlus4E[23] ),
    .Q(\rvcpu.dp.plem.PCPlus4M[23] ));
 sky130_fd_sc_hd__dfxtp_1 _31530_ (.CLK(clk),
    .D(\rvcpu.dp.plde.PCPlus4E[24] ),
    .Q(\rvcpu.dp.plem.PCPlus4M[24] ));
 sky130_fd_sc_hd__dfxtp_1 _31531_ (.CLK(clk),
    .D(\rvcpu.dp.plde.PCPlus4E[25] ),
    .Q(\rvcpu.dp.plem.PCPlus4M[25] ));
 sky130_fd_sc_hd__dfxtp_1 _31532_ (.CLK(clk),
    .D(\rvcpu.dp.plde.PCPlus4E[26] ),
    .Q(\rvcpu.dp.plem.PCPlus4M[26] ));
 sky130_fd_sc_hd__dfxtp_1 _31533_ (.CLK(clk),
    .D(\rvcpu.dp.plde.PCPlus4E[27] ),
    .Q(\rvcpu.dp.plem.PCPlus4M[27] ));
 sky130_fd_sc_hd__dfxtp_1 _31534_ (.CLK(clk),
    .D(\rvcpu.dp.plde.PCPlus4E[28] ),
    .Q(\rvcpu.dp.plem.PCPlus4M[28] ));
 sky130_fd_sc_hd__dfxtp_1 _31535_ (.CLK(clk),
    .D(\rvcpu.dp.plde.PCPlus4E[29] ),
    .Q(\rvcpu.dp.plem.PCPlus4M[29] ));
 sky130_fd_sc_hd__dfxtp_1 _31536_ (.CLK(clk),
    .D(\rvcpu.dp.plde.PCPlus4E[30] ),
    .Q(\rvcpu.dp.plem.PCPlus4M[30] ));
 sky130_fd_sc_hd__dfxtp_1 _31537_ (.CLK(clk),
    .D(\rvcpu.dp.plde.PCPlus4E[31] ),
    .Q(\rvcpu.dp.plem.PCPlus4M[31] ));
 sky130_fd_sc_hd__dfxtp_1 _31538_ (.CLK(clk),
    .D(\rvcpu.dp.plde.funct3E[0] ),
    .Q(\rvcpu.dp.plem.funct3M[0] ));
 sky130_fd_sc_hd__dfxtp_1 _31539_ (.CLK(clk),
    .D(\rvcpu.dp.plde.funct3E[1] ),
    .Q(\rvcpu.dp.plem.funct3M[1] ));
 sky130_fd_sc_hd__dfxtp_1 _31540_ (.CLK(clk),
    .D(\rvcpu.dp.plde.funct3E[2] ),
    .Q(\rvcpu.dp.plem.funct3M[2] ));
 sky130_fd_sc_hd__dfxtp_1 _31541_ (.CLK(clk),
    .D(\rvcpu.dp.plde.MemWriteE ),
    .Q(\rvcpu.dp.plem.MemWriteM ));
 sky130_fd_sc_hd__dfxtp_1 _31542_ (.CLK(clk),
    .D(\rvcpu.dp.plde.RdE[0] ),
    .Q(\rvcpu.dp.plem.RdM[0] ));
 sky130_fd_sc_hd__dfxtp_1 _31543_ (.CLK(clk),
    .D(\rvcpu.dp.plde.RdE[1] ),
    .Q(\rvcpu.dp.plem.RdM[1] ));
 sky130_fd_sc_hd__dfxtp_1 _31544_ (.CLK(clk),
    .D(\rvcpu.dp.plde.RdE[2] ),
    .Q(\rvcpu.dp.plem.RdM[2] ));
 sky130_fd_sc_hd__dfxtp_1 _31545_ (.CLK(clk),
    .D(\rvcpu.dp.plde.RdE[3] ),
    .Q(\rvcpu.dp.plem.RdM[3] ));
 sky130_fd_sc_hd__dfxtp_1 _31546_ (.CLK(clk),
    .D(\rvcpu.dp.plde.RdE[4] ),
    .Q(\rvcpu.dp.plem.RdM[4] ));
 sky130_fd_sc_hd__dfxtp_1 _31547_ (.CLK(clk),
    .D(\rvcpu.dp.plde.RegWriteE ),
    .Q(\rvcpu.dp.plem.RegWriteM ));
 sky130_fd_sc_hd__dfxtp_2 _31548_ (.CLK(clk),
    .D(\rvcpu.dp.plem.ResultSrcM[0] ),
    .Q(\rvcpu.dp.plmw.ResultSrcW[0] ));
 sky130_fd_sc_hd__dfxtp_1 _31549_ (.CLK(clk),
    .D(\rvcpu.dp.plem.ResultSrcM[1] ),
    .Q(\rvcpu.dp.plmw.ResultSrcW[1] ));
 sky130_fd_sc_hd__dfxtp_1 _31550_ (.CLK(clk),
    .D(\datamem.rd_data_mem[0] ),
    .Q(\rvcpu.dp.plmw.ReadDataW[0] ));
 sky130_fd_sc_hd__dfxtp_1 _31551_ (.CLK(clk),
    .D(\datamem.rd_data_mem[1] ),
    .Q(\rvcpu.dp.plmw.ReadDataW[1] ));
 sky130_fd_sc_hd__dfxtp_1 _31552_ (.CLK(clk),
    .D(\datamem.rd_data_mem[2] ),
    .Q(\rvcpu.dp.plmw.ReadDataW[2] ));
 sky130_fd_sc_hd__dfxtp_1 _31553_ (.CLK(clk),
    .D(\datamem.rd_data_mem[3] ),
    .Q(\rvcpu.dp.plmw.ReadDataW[3] ));
 sky130_fd_sc_hd__dfxtp_1 _31554_ (.CLK(clk),
    .D(\datamem.rd_data_mem[4] ),
    .Q(\rvcpu.dp.plmw.ReadDataW[4] ));
 sky130_fd_sc_hd__dfxtp_1 _31555_ (.CLK(clk),
    .D(\datamem.rd_data_mem[5] ),
    .Q(\rvcpu.dp.plmw.ReadDataW[5] ));
 sky130_fd_sc_hd__dfxtp_1 _31556_ (.CLK(clk),
    .D(\datamem.rd_data_mem[6] ),
    .Q(\rvcpu.dp.plmw.ReadDataW[6] ));
 sky130_fd_sc_hd__dfxtp_1 _31557_ (.CLK(clk),
    .D(\datamem.rd_data_mem[7] ),
    .Q(\rvcpu.dp.plmw.ReadDataW[7] ));
 sky130_fd_sc_hd__dfxtp_1 _31558_ (.CLK(clk),
    .D(\datamem.rd_data_mem[8] ),
    .Q(\rvcpu.dp.plmw.ReadDataW[8] ));
 sky130_fd_sc_hd__dfxtp_1 _31559_ (.CLK(clk),
    .D(\datamem.rd_data_mem[9] ),
    .Q(\rvcpu.dp.plmw.ReadDataW[9] ));
 sky130_fd_sc_hd__dfxtp_1 _31560_ (.CLK(clk),
    .D(\datamem.rd_data_mem[10] ),
    .Q(\rvcpu.dp.plmw.ReadDataW[10] ));
 sky130_fd_sc_hd__dfxtp_1 _31561_ (.CLK(clk),
    .D(\datamem.rd_data_mem[11] ),
    .Q(\rvcpu.dp.plmw.ReadDataW[11] ));
 sky130_fd_sc_hd__dfxtp_1 _31562_ (.CLK(clk),
    .D(\datamem.rd_data_mem[12] ),
    .Q(\rvcpu.dp.plmw.ReadDataW[12] ));
 sky130_fd_sc_hd__dfxtp_1 _31563_ (.CLK(clk),
    .D(\datamem.rd_data_mem[13] ),
    .Q(\rvcpu.dp.plmw.ReadDataW[13] ));
 sky130_fd_sc_hd__dfxtp_1 _31564_ (.CLK(clk),
    .D(\datamem.rd_data_mem[14] ),
    .Q(\rvcpu.dp.plmw.ReadDataW[14] ));
 sky130_fd_sc_hd__dfxtp_1 _31565_ (.CLK(clk),
    .D(\datamem.rd_data_mem[15] ),
    .Q(\rvcpu.dp.plmw.ReadDataW[15] ));
 sky130_fd_sc_hd__dfxtp_1 _31566_ (.CLK(clk),
    .D(\datamem.rd_data_mem[16] ),
    .Q(\rvcpu.dp.plmw.ReadDataW[16] ));
 sky130_fd_sc_hd__dfxtp_1 _31567_ (.CLK(clk),
    .D(\datamem.rd_data_mem[17] ),
    .Q(\rvcpu.dp.plmw.ReadDataW[17] ));
 sky130_fd_sc_hd__dfxtp_1 _31568_ (.CLK(clk),
    .D(\datamem.rd_data_mem[18] ),
    .Q(\rvcpu.dp.plmw.ReadDataW[18] ));
 sky130_fd_sc_hd__dfxtp_1 _31569_ (.CLK(clk),
    .D(\datamem.rd_data_mem[19] ),
    .Q(\rvcpu.dp.plmw.ReadDataW[19] ));
 sky130_fd_sc_hd__dfxtp_1 _31570_ (.CLK(clk),
    .D(\datamem.rd_data_mem[20] ),
    .Q(\rvcpu.dp.plmw.ReadDataW[20] ));
 sky130_fd_sc_hd__dfxtp_1 _31571_ (.CLK(clk),
    .D(\datamem.rd_data_mem[21] ),
    .Q(\rvcpu.dp.plmw.ReadDataW[21] ));
 sky130_fd_sc_hd__dfxtp_1 _31572_ (.CLK(clk),
    .D(\datamem.rd_data_mem[22] ),
    .Q(\rvcpu.dp.plmw.ReadDataW[22] ));
 sky130_fd_sc_hd__dfxtp_1 _31573_ (.CLK(clk),
    .D(\datamem.rd_data_mem[23] ),
    .Q(\rvcpu.dp.plmw.ReadDataW[23] ));
 sky130_fd_sc_hd__dfxtp_1 _31574_ (.CLK(clk),
    .D(\datamem.rd_data_mem[24] ),
    .Q(\rvcpu.dp.plmw.ReadDataW[24] ));
 sky130_fd_sc_hd__dfxtp_1 _31575_ (.CLK(clk),
    .D(\datamem.rd_data_mem[25] ),
    .Q(\rvcpu.dp.plmw.ReadDataW[25] ));
 sky130_fd_sc_hd__dfxtp_1 _31576_ (.CLK(clk),
    .D(\datamem.rd_data_mem[26] ),
    .Q(\rvcpu.dp.plmw.ReadDataW[26] ));
 sky130_fd_sc_hd__dfxtp_1 _31577_ (.CLK(clk),
    .D(\datamem.rd_data_mem[27] ),
    .Q(\rvcpu.dp.plmw.ReadDataW[27] ));
 sky130_fd_sc_hd__dfxtp_1 _31578_ (.CLK(clk),
    .D(\datamem.rd_data_mem[28] ),
    .Q(\rvcpu.dp.plmw.ReadDataW[28] ));
 sky130_fd_sc_hd__dfxtp_1 _31579_ (.CLK(clk),
    .D(\datamem.rd_data_mem[29] ),
    .Q(\rvcpu.dp.plmw.ReadDataW[29] ));
 sky130_fd_sc_hd__dfxtp_1 _31580_ (.CLK(clk),
    .D(\datamem.rd_data_mem[30] ),
    .Q(\rvcpu.dp.plmw.ReadDataW[30] ));
 sky130_fd_sc_hd__dfxtp_1 _31581_ (.CLK(clk),
    .D(\datamem.rd_data_mem[31] ),
    .Q(\rvcpu.dp.plmw.ReadDataW[31] ));
 sky130_fd_sc_hd__dfxtp_1 _31582_ (.CLK(clk),
    .D(\rvcpu.dp.plem.PCPlus4M[0] ),
    .Q(\rvcpu.dp.plmw.PCPlus4W[0] ));
 sky130_fd_sc_hd__dfxtp_1 _31583_ (.CLK(clk),
    .D(\rvcpu.dp.plem.PCPlus4M[1] ),
    .Q(\rvcpu.dp.plmw.PCPlus4W[1] ));
 sky130_fd_sc_hd__dfxtp_1 _31584_ (.CLK(clk),
    .D(\rvcpu.dp.plem.PCPlus4M[2] ),
    .Q(\rvcpu.dp.plmw.PCPlus4W[2] ));
 sky130_fd_sc_hd__dfxtp_1 _31585_ (.CLK(clk),
    .D(\rvcpu.dp.plem.PCPlus4M[3] ),
    .Q(\rvcpu.dp.plmw.PCPlus4W[3] ));
 sky130_fd_sc_hd__dfxtp_1 _31586_ (.CLK(clk),
    .D(\rvcpu.dp.plem.PCPlus4M[4] ),
    .Q(\rvcpu.dp.plmw.PCPlus4W[4] ));
 sky130_fd_sc_hd__dfxtp_1 _31587_ (.CLK(clk),
    .D(\rvcpu.dp.plem.PCPlus4M[5] ),
    .Q(\rvcpu.dp.plmw.PCPlus4W[5] ));
 sky130_fd_sc_hd__dfxtp_1 _31588_ (.CLK(clk),
    .D(\rvcpu.dp.plem.PCPlus4M[6] ),
    .Q(\rvcpu.dp.plmw.PCPlus4W[6] ));
 sky130_fd_sc_hd__dfxtp_1 _31589_ (.CLK(clk),
    .D(\rvcpu.dp.plem.PCPlus4M[7] ),
    .Q(\rvcpu.dp.plmw.PCPlus4W[7] ));
 sky130_fd_sc_hd__dfxtp_1 _31590_ (.CLK(clk),
    .D(\rvcpu.dp.plem.PCPlus4M[8] ),
    .Q(\rvcpu.dp.plmw.PCPlus4W[8] ));
 sky130_fd_sc_hd__dfxtp_1 _31591_ (.CLK(clk),
    .D(\rvcpu.dp.plem.PCPlus4M[9] ),
    .Q(\rvcpu.dp.plmw.PCPlus4W[9] ));
 sky130_fd_sc_hd__dfxtp_1 _31592_ (.CLK(clk),
    .D(\rvcpu.dp.plem.PCPlus4M[10] ),
    .Q(\rvcpu.dp.plmw.PCPlus4W[10] ));
 sky130_fd_sc_hd__dfxtp_1 _31593_ (.CLK(clk),
    .D(\rvcpu.dp.plem.PCPlus4M[11] ),
    .Q(\rvcpu.dp.plmw.PCPlus4W[11] ));
 sky130_fd_sc_hd__dfxtp_1 _31594_ (.CLK(clk),
    .D(\rvcpu.dp.plem.PCPlus4M[12] ),
    .Q(\rvcpu.dp.plmw.PCPlus4W[12] ));
 sky130_fd_sc_hd__dfxtp_1 _31595_ (.CLK(clk),
    .D(\rvcpu.dp.plem.PCPlus4M[13] ),
    .Q(\rvcpu.dp.plmw.PCPlus4W[13] ));
 sky130_fd_sc_hd__dfxtp_1 _31596_ (.CLK(clk),
    .D(\rvcpu.dp.plem.PCPlus4M[14] ),
    .Q(\rvcpu.dp.plmw.PCPlus4W[14] ));
 sky130_fd_sc_hd__dfxtp_1 _31597_ (.CLK(clk),
    .D(\rvcpu.dp.plem.PCPlus4M[15] ),
    .Q(\rvcpu.dp.plmw.PCPlus4W[15] ));
 sky130_fd_sc_hd__dfxtp_1 _31598_ (.CLK(clk),
    .D(\rvcpu.dp.plem.PCPlus4M[16] ),
    .Q(\rvcpu.dp.plmw.PCPlus4W[16] ));
 sky130_fd_sc_hd__dfxtp_1 _31599_ (.CLK(clk),
    .D(\rvcpu.dp.plem.PCPlus4M[17] ),
    .Q(\rvcpu.dp.plmw.PCPlus4W[17] ));
 sky130_fd_sc_hd__dfxtp_1 _31600_ (.CLK(clk),
    .D(\rvcpu.dp.plem.PCPlus4M[18] ),
    .Q(\rvcpu.dp.plmw.PCPlus4W[18] ));
 sky130_fd_sc_hd__dfxtp_1 _31601_ (.CLK(clk),
    .D(\rvcpu.dp.plem.PCPlus4M[19] ),
    .Q(\rvcpu.dp.plmw.PCPlus4W[19] ));
 sky130_fd_sc_hd__dfxtp_1 _31602_ (.CLK(clk),
    .D(\rvcpu.dp.plem.PCPlus4M[20] ),
    .Q(\rvcpu.dp.plmw.PCPlus4W[20] ));
 sky130_fd_sc_hd__dfxtp_1 _31603_ (.CLK(clk),
    .D(\rvcpu.dp.plem.PCPlus4M[21] ),
    .Q(\rvcpu.dp.plmw.PCPlus4W[21] ));
 sky130_fd_sc_hd__dfxtp_1 _31604_ (.CLK(clk),
    .D(\rvcpu.dp.plem.PCPlus4M[22] ),
    .Q(\rvcpu.dp.plmw.PCPlus4W[22] ));
 sky130_fd_sc_hd__dfxtp_1 _31605_ (.CLK(clk),
    .D(\rvcpu.dp.plem.PCPlus4M[23] ),
    .Q(\rvcpu.dp.plmw.PCPlus4W[23] ));
 sky130_fd_sc_hd__dfxtp_1 _31606_ (.CLK(clk),
    .D(\rvcpu.dp.plem.PCPlus4M[24] ),
    .Q(\rvcpu.dp.plmw.PCPlus4W[24] ));
 sky130_fd_sc_hd__dfxtp_1 _31607_ (.CLK(clk),
    .D(\rvcpu.dp.plem.PCPlus4M[25] ),
    .Q(\rvcpu.dp.plmw.PCPlus4W[25] ));
 sky130_fd_sc_hd__dfxtp_1 _31608_ (.CLK(clk),
    .D(\rvcpu.dp.plem.PCPlus4M[26] ),
    .Q(\rvcpu.dp.plmw.PCPlus4W[26] ));
 sky130_fd_sc_hd__dfxtp_1 _31609_ (.CLK(clk),
    .D(\rvcpu.dp.plem.PCPlus4M[27] ),
    .Q(\rvcpu.dp.plmw.PCPlus4W[27] ));
 sky130_fd_sc_hd__dfxtp_1 _31610_ (.CLK(clk),
    .D(\rvcpu.dp.plem.PCPlus4M[28] ),
    .Q(\rvcpu.dp.plmw.PCPlus4W[28] ));
 sky130_fd_sc_hd__dfxtp_1 _31611_ (.CLK(clk),
    .D(\rvcpu.dp.plem.PCPlus4M[29] ),
    .Q(\rvcpu.dp.plmw.PCPlus4W[29] ));
 sky130_fd_sc_hd__dfxtp_1 _31612_ (.CLK(clk),
    .D(\rvcpu.dp.plem.PCPlus4M[30] ),
    .Q(\rvcpu.dp.plmw.PCPlus4W[30] ));
 sky130_fd_sc_hd__dfxtp_1 _31613_ (.CLK(clk),
    .D(\rvcpu.dp.plem.PCPlus4M[31] ),
    .Q(\rvcpu.dp.plmw.PCPlus4W[31] ));
 sky130_fd_sc_hd__dfxtp_2 _31614_ (.CLK(clk),
    .D(\rvcpu.dp.plem.RdM[0] ),
    .Q(\rvcpu.dp.plmw.RdW[0] ));
 sky130_fd_sc_hd__dfxtp_4 _31615_ (.CLK(clk),
    .D(\rvcpu.dp.plem.RdM[1] ),
    .Q(\rvcpu.dp.plmw.RdW[1] ));
 sky130_fd_sc_hd__dfxtp_1 _31616_ (.CLK(clk),
    .D(\rvcpu.dp.plem.RdM[2] ),
    .Q(\rvcpu.dp.plmw.RdW[2] ));
 sky130_fd_sc_hd__dfxtp_4 _31617_ (.CLK(clk),
    .D(\rvcpu.dp.plem.RdM[3] ),
    .Q(\rvcpu.dp.plmw.RdW[3] ));
 sky130_fd_sc_hd__dfxtp_1 _31618_ (.CLK(clk),
    .D(\rvcpu.dp.plem.RdM[4] ),
    .Q(\rvcpu.dp.plmw.RdW[4] ));
 sky130_fd_sc_hd__dfxtp_2 _31619_ (.CLK(clk),
    .D(\rvcpu.dp.plem.RegWriteM ),
    .Q(\rvcpu.dp.plmw.RegWriteW ));
 sky130_fd_sc_hd__dfxtp_1 _31620_ (.CLK(clk),
    .D(\rvcpu.dp.plem.lAuiPCM[0] ),
    .Q(\rvcpu.dp.plmw.lAuiPCW[0] ));
 sky130_fd_sc_hd__dfxtp_1 _31621_ (.CLK(clk),
    .D(\rvcpu.dp.plem.lAuiPCM[1] ),
    .Q(\rvcpu.dp.plmw.lAuiPCW[1] ));
 sky130_fd_sc_hd__dfxtp_1 _31622_ (.CLK(clk),
    .D(\rvcpu.dp.plem.lAuiPCM[2] ),
    .Q(\rvcpu.dp.plmw.lAuiPCW[2] ));
 sky130_fd_sc_hd__dfxtp_1 _31623_ (.CLK(clk),
    .D(\rvcpu.dp.plem.lAuiPCM[3] ),
    .Q(\rvcpu.dp.plmw.lAuiPCW[3] ));
 sky130_fd_sc_hd__dfxtp_1 _31624_ (.CLK(clk),
    .D(\rvcpu.dp.plem.lAuiPCM[4] ),
    .Q(\rvcpu.dp.plmw.lAuiPCW[4] ));
 sky130_fd_sc_hd__dfxtp_1 _31625_ (.CLK(clk),
    .D(\rvcpu.dp.plem.lAuiPCM[5] ),
    .Q(\rvcpu.dp.plmw.lAuiPCW[5] ));
 sky130_fd_sc_hd__dfxtp_1 _31626_ (.CLK(clk),
    .D(\rvcpu.dp.plem.lAuiPCM[6] ),
    .Q(\rvcpu.dp.plmw.lAuiPCW[6] ));
 sky130_fd_sc_hd__dfxtp_1 _31627_ (.CLK(clk),
    .D(\rvcpu.dp.plem.lAuiPCM[7] ),
    .Q(\rvcpu.dp.plmw.lAuiPCW[7] ));
 sky130_fd_sc_hd__dfxtp_1 _31628_ (.CLK(clk),
    .D(\rvcpu.dp.plem.lAuiPCM[8] ),
    .Q(\rvcpu.dp.plmw.lAuiPCW[8] ));
 sky130_fd_sc_hd__dfxtp_1 _31629_ (.CLK(clk),
    .D(\rvcpu.dp.plem.lAuiPCM[9] ),
    .Q(\rvcpu.dp.plmw.lAuiPCW[9] ));
 sky130_fd_sc_hd__dfxtp_1 _31630_ (.CLK(clk),
    .D(\rvcpu.dp.plem.lAuiPCM[10] ),
    .Q(\rvcpu.dp.plmw.lAuiPCW[10] ));
 sky130_fd_sc_hd__dfxtp_1 _31631_ (.CLK(clk),
    .D(\rvcpu.dp.plem.lAuiPCM[11] ),
    .Q(\rvcpu.dp.plmw.lAuiPCW[11] ));
 sky130_fd_sc_hd__dfxtp_1 _31632_ (.CLK(clk),
    .D(\rvcpu.dp.plem.lAuiPCM[12] ),
    .Q(\rvcpu.dp.plmw.lAuiPCW[12] ));
 sky130_fd_sc_hd__dfxtp_1 _31633_ (.CLK(clk),
    .D(\rvcpu.dp.plem.lAuiPCM[13] ),
    .Q(\rvcpu.dp.plmw.lAuiPCW[13] ));
 sky130_fd_sc_hd__dfxtp_1 _31634_ (.CLK(clk),
    .D(\rvcpu.dp.plem.lAuiPCM[14] ),
    .Q(\rvcpu.dp.plmw.lAuiPCW[14] ));
 sky130_fd_sc_hd__dfxtp_1 _31635_ (.CLK(clk),
    .D(\rvcpu.dp.plem.lAuiPCM[15] ),
    .Q(\rvcpu.dp.plmw.lAuiPCW[15] ));
 sky130_fd_sc_hd__dfxtp_1 _31636_ (.CLK(clk),
    .D(\rvcpu.dp.plem.lAuiPCM[16] ),
    .Q(\rvcpu.dp.plmw.lAuiPCW[16] ));
 sky130_fd_sc_hd__dfxtp_1 _31637_ (.CLK(clk),
    .D(\rvcpu.dp.plem.lAuiPCM[17] ),
    .Q(\rvcpu.dp.plmw.lAuiPCW[17] ));
 sky130_fd_sc_hd__dfxtp_1 _31638_ (.CLK(clk),
    .D(\rvcpu.dp.plem.lAuiPCM[18] ),
    .Q(\rvcpu.dp.plmw.lAuiPCW[18] ));
 sky130_fd_sc_hd__dfxtp_1 _31639_ (.CLK(clk),
    .D(\rvcpu.dp.plem.lAuiPCM[19] ),
    .Q(\rvcpu.dp.plmw.lAuiPCW[19] ));
 sky130_fd_sc_hd__dfxtp_1 _31640_ (.CLK(clk),
    .D(\rvcpu.dp.plem.lAuiPCM[20] ),
    .Q(\rvcpu.dp.plmw.lAuiPCW[20] ));
 sky130_fd_sc_hd__dfxtp_1 _31641_ (.CLK(clk),
    .D(\rvcpu.dp.plem.lAuiPCM[21] ),
    .Q(\rvcpu.dp.plmw.lAuiPCW[21] ));
 sky130_fd_sc_hd__dfxtp_1 _31642_ (.CLK(clk),
    .D(\rvcpu.dp.plem.lAuiPCM[22] ),
    .Q(\rvcpu.dp.plmw.lAuiPCW[22] ));
 sky130_fd_sc_hd__dfxtp_1 _31643_ (.CLK(clk),
    .D(\rvcpu.dp.plem.lAuiPCM[23] ),
    .Q(\rvcpu.dp.plmw.lAuiPCW[23] ));
 sky130_fd_sc_hd__dfxtp_1 _31644_ (.CLK(clk),
    .D(\rvcpu.dp.plem.lAuiPCM[24] ),
    .Q(\rvcpu.dp.plmw.lAuiPCW[24] ));
 sky130_fd_sc_hd__dfxtp_1 _31645_ (.CLK(clk),
    .D(\rvcpu.dp.plem.lAuiPCM[25] ),
    .Q(\rvcpu.dp.plmw.lAuiPCW[25] ));
 sky130_fd_sc_hd__dfxtp_1 _31646_ (.CLK(clk),
    .D(\rvcpu.dp.plem.lAuiPCM[26] ),
    .Q(\rvcpu.dp.plmw.lAuiPCW[26] ));
 sky130_fd_sc_hd__dfxtp_1 _31647_ (.CLK(clk),
    .D(\rvcpu.dp.plem.lAuiPCM[27] ),
    .Q(\rvcpu.dp.plmw.lAuiPCW[27] ));
 sky130_fd_sc_hd__dfxtp_1 _31648_ (.CLK(clk),
    .D(\rvcpu.dp.plem.lAuiPCM[28] ),
    .Q(\rvcpu.dp.plmw.lAuiPCW[28] ));
 sky130_fd_sc_hd__dfxtp_1 _31649_ (.CLK(clk),
    .D(\rvcpu.dp.plem.lAuiPCM[29] ),
    .Q(\rvcpu.dp.plmw.lAuiPCW[29] ));
 sky130_fd_sc_hd__dfxtp_1 _31650_ (.CLK(clk),
    .D(\rvcpu.dp.plem.lAuiPCM[30] ),
    .Q(\rvcpu.dp.plmw.lAuiPCW[30] ));
 sky130_fd_sc_hd__dfxtp_1 _31651_ (.CLK(clk),
    .D(\rvcpu.dp.plem.lAuiPCM[31] ),
    .Q(\rvcpu.dp.plmw.lAuiPCW[31] ));
 sky130_fd_sc_hd__dfxtp_1 _31652_ (.CLK(clk),
    .D(\rvcpu.dp.plem.ALUResultM[0] ),
    .Q(\rvcpu.dp.plmw.ALUResultW[0] ));
 sky130_fd_sc_hd__dfxtp_1 _31653_ (.CLK(clk),
    .D(\rvcpu.dp.plem.ALUResultM[1] ),
    .Q(\rvcpu.dp.plmw.ALUResultW[1] ));
 sky130_fd_sc_hd__dfxtp_1 _31654_ (.CLK(clk),
    .D(\rvcpu.dp.plem.ALUResultM[2] ),
    .Q(\rvcpu.dp.plmw.ALUResultW[2] ));
 sky130_fd_sc_hd__dfxtp_1 _31655_ (.CLK(clk),
    .D(\rvcpu.dp.plem.ALUResultM[3] ),
    .Q(\rvcpu.dp.plmw.ALUResultW[3] ));
 sky130_fd_sc_hd__dfxtp_1 _31656_ (.CLK(clk),
    .D(\rvcpu.dp.plem.ALUResultM[4] ),
    .Q(\rvcpu.dp.plmw.ALUResultW[4] ));
 sky130_fd_sc_hd__dfxtp_1 _31657_ (.CLK(clk),
    .D(\rvcpu.dp.plem.ALUResultM[5] ),
    .Q(\rvcpu.dp.plmw.ALUResultW[5] ));
 sky130_fd_sc_hd__dfxtp_1 _31658_ (.CLK(clk),
    .D(\rvcpu.dp.plem.ALUResultM[6] ),
    .Q(\rvcpu.dp.plmw.ALUResultW[6] ));
 sky130_fd_sc_hd__dfxtp_1 _31659_ (.CLK(clk),
    .D(\rvcpu.dp.plem.ALUResultM[7] ),
    .Q(\rvcpu.dp.plmw.ALUResultW[7] ));
 sky130_fd_sc_hd__dfxtp_1 _31660_ (.CLK(clk),
    .D(\rvcpu.dp.plem.ALUResultM[8] ),
    .Q(\rvcpu.dp.plmw.ALUResultW[8] ));
 sky130_fd_sc_hd__dfxtp_1 _31661_ (.CLK(clk),
    .D(\rvcpu.dp.plem.ALUResultM[9] ),
    .Q(\rvcpu.dp.plmw.ALUResultW[9] ));
 sky130_fd_sc_hd__dfxtp_1 _31662_ (.CLK(clk),
    .D(\rvcpu.dp.plem.ALUResultM[10] ),
    .Q(\rvcpu.dp.plmw.ALUResultW[10] ));
 sky130_fd_sc_hd__dfxtp_1 _31663_ (.CLK(clk),
    .D(\rvcpu.dp.plem.ALUResultM[11] ),
    .Q(\rvcpu.dp.plmw.ALUResultW[11] ));
 sky130_fd_sc_hd__dfxtp_1 _31664_ (.CLK(clk),
    .D(\rvcpu.dp.plem.ALUResultM[12] ),
    .Q(\rvcpu.dp.plmw.ALUResultW[12] ));
 sky130_fd_sc_hd__dfxtp_1 _31665_ (.CLK(clk),
    .D(\rvcpu.dp.plem.ALUResultM[13] ),
    .Q(\rvcpu.dp.plmw.ALUResultW[13] ));
 sky130_fd_sc_hd__dfxtp_1 _31666_ (.CLK(clk),
    .D(\rvcpu.dp.plem.ALUResultM[14] ),
    .Q(\rvcpu.dp.plmw.ALUResultW[14] ));
 sky130_fd_sc_hd__dfxtp_1 _31667_ (.CLK(clk),
    .D(\rvcpu.dp.plem.ALUResultM[15] ),
    .Q(\rvcpu.dp.plmw.ALUResultW[15] ));
 sky130_fd_sc_hd__dfxtp_1 _31668_ (.CLK(clk),
    .D(\rvcpu.dp.plem.ALUResultM[16] ),
    .Q(\rvcpu.dp.plmw.ALUResultW[16] ));
 sky130_fd_sc_hd__dfxtp_1 _31669_ (.CLK(clk),
    .D(\rvcpu.dp.plem.ALUResultM[17] ),
    .Q(\rvcpu.dp.plmw.ALUResultW[17] ));
 sky130_fd_sc_hd__dfxtp_1 _31670_ (.CLK(clk),
    .D(\rvcpu.dp.plem.ALUResultM[18] ),
    .Q(\rvcpu.dp.plmw.ALUResultW[18] ));
 sky130_fd_sc_hd__dfxtp_1 _31671_ (.CLK(clk),
    .D(\rvcpu.dp.plem.ALUResultM[19] ),
    .Q(\rvcpu.dp.plmw.ALUResultW[19] ));
 sky130_fd_sc_hd__dfxtp_1 _31672_ (.CLK(clk),
    .D(\rvcpu.dp.plem.ALUResultM[20] ),
    .Q(\rvcpu.dp.plmw.ALUResultW[20] ));
 sky130_fd_sc_hd__dfxtp_1 _31673_ (.CLK(clk),
    .D(\rvcpu.dp.plem.ALUResultM[21] ),
    .Q(\rvcpu.dp.plmw.ALUResultW[21] ));
 sky130_fd_sc_hd__dfxtp_1 _31674_ (.CLK(clk),
    .D(\rvcpu.dp.plem.ALUResultM[22] ),
    .Q(\rvcpu.dp.plmw.ALUResultW[22] ));
 sky130_fd_sc_hd__dfxtp_1 _31675_ (.CLK(clk),
    .D(\rvcpu.dp.plem.ALUResultM[23] ),
    .Q(\rvcpu.dp.plmw.ALUResultW[23] ));
 sky130_fd_sc_hd__dfxtp_1 _31676_ (.CLK(clk),
    .D(\rvcpu.dp.plem.ALUResultM[24] ),
    .Q(\rvcpu.dp.plmw.ALUResultW[24] ));
 sky130_fd_sc_hd__dfxtp_1 _31677_ (.CLK(clk),
    .D(\rvcpu.dp.plem.ALUResultM[25] ),
    .Q(\rvcpu.dp.plmw.ALUResultW[25] ));
 sky130_fd_sc_hd__dfxtp_1 _31678_ (.CLK(clk),
    .D(\rvcpu.dp.plem.ALUResultM[26] ),
    .Q(\rvcpu.dp.plmw.ALUResultW[26] ));
 sky130_fd_sc_hd__dfxtp_1 _31679_ (.CLK(clk),
    .D(\rvcpu.dp.plem.ALUResultM[27] ),
    .Q(\rvcpu.dp.plmw.ALUResultW[27] ));
 sky130_fd_sc_hd__dfxtp_1 _31680_ (.CLK(clk),
    .D(\rvcpu.dp.plem.ALUResultM[28] ),
    .Q(\rvcpu.dp.plmw.ALUResultW[28] ));
 sky130_fd_sc_hd__dfxtp_1 _31681_ (.CLK(clk),
    .D(\rvcpu.dp.plem.ALUResultM[29] ),
    .Q(\rvcpu.dp.plmw.ALUResultW[29] ));
 sky130_fd_sc_hd__dfxtp_1 _31682_ (.CLK(clk),
    .D(\rvcpu.dp.plem.ALUResultM[30] ),
    .Q(\rvcpu.dp.plmw.ALUResultW[30] ));
 sky130_fd_sc_hd__dfxtp_1 _31683_ (.CLK(clk),
    .D(\rvcpu.dp.plem.ALUResultM[31] ),
    .Q(\rvcpu.dp.plmw.ALUResultW[31] ));
 sky130_fd_sc_hd__dfxtp_2 _31684_ (.CLK(clk),
    .D(_03142_),
    .Q(\rvcpu.dp.pcreg.q[2] ));
 sky130_fd_sc_hd__dfxtp_4 _31685_ (.CLK(clk),
    .D(_03143_),
    .Q(\rvcpu.dp.pcreg.q[3] ));
 sky130_fd_sc_hd__dfxtp_2 _31686_ (.CLK(clk),
    .D(_03144_),
    .Q(\rvcpu.dp.pcreg.q[4] ));
 sky130_fd_sc_hd__dfxtp_4 _31687_ (.CLK(clk),
    .D(_03145_),
    .Q(\rvcpu.dp.pcreg.q[5] ));
 sky130_fd_sc_hd__dfxtp_2 _31688_ (.CLK(clk),
    .D(_03146_),
    .Q(\rvcpu.dp.pcreg.q[6] ));
 sky130_fd_sc_hd__dfxtp_1 _31689_ (.CLK(clk),
    .D(_03147_),
    .Q(\rvcpu.dp.pcreg.q[7] ));
 sky130_fd_sc_hd__dfxtp_2 _31690_ (.CLK(clk),
    .D(_03148_),
    .Q(\rvcpu.dp.pcreg.q[8] ));
 sky130_fd_sc_hd__dfxtp_4 _31691_ (.CLK(clk),
    .D(_03149_),
    .Q(\rvcpu.dp.pcreg.q[9] ));
 sky130_fd_sc_hd__dfxtp_1 _31692_ (.CLK(clk),
    .D(_03150_),
    .Q(\rvcpu.dp.pcreg.q[10] ));
 sky130_fd_sc_hd__dfxtp_1 _31693_ (.CLK(clk),
    .D(_03151_),
    .Q(\rvcpu.dp.pcreg.q[11] ));
 sky130_fd_sc_hd__dfxtp_1 _31694_ (.CLK(clk),
    .D(_03152_),
    .Q(\rvcpu.dp.pcreg.q[12] ));
 sky130_fd_sc_hd__dfxtp_1 _31695_ (.CLK(clk),
    .D(_03153_),
    .Q(\rvcpu.dp.pcreg.q[13] ));
 sky130_fd_sc_hd__dfxtp_1 _31696_ (.CLK(clk),
    .D(_03154_),
    .Q(\rvcpu.dp.pcreg.q[14] ));
 sky130_fd_sc_hd__dfxtp_1 _31697_ (.CLK(clk),
    .D(_03155_),
    .Q(\rvcpu.dp.pcreg.q[15] ));
 sky130_fd_sc_hd__dfxtp_1 _31698_ (.CLK(clk),
    .D(_03156_),
    .Q(\rvcpu.dp.pcreg.q[16] ));
 sky130_fd_sc_hd__dfxtp_1 _31699_ (.CLK(clk),
    .D(_03157_),
    .Q(\rvcpu.dp.pcreg.q[17] ));
 sky130_fd_sc_hd__dfxtp_1 _31700_ (.CLK(clk),
    .D(_03158_),
    .Q(\rvcpu.dp.pcreg.q[18] ));
 sky130_fd_sc_hd__dfxtp_1 _31701_ (.CLK(clk),
    .D(_03159_),
    .Q(\rvcpu.dp.pcreg.q[19] ));
 sky130_fd_sc_hd__dfxtp_1 _31702_ (.CLK(clk),
    .D(_03160_),
    .Q(\rvcpu.dp.pcreg.q[20] ));
 sky130_fd_sc_hd__dfxtp_1 _31703_ (.CLK(clk),
    .D(_03161_),
    .Q(\rvcpu.dp.pcreg.q[21] ));
 sky130_fd_sc_hd__dfxtp_1 _31704_ (.CLK(clk),
    .D(_03162_),
    .Q(\rvcpu.dp.pcreg.q[22] ));
 sky130_fd_sc_hd__dfxtp_1 _31705_ (.CLK(clk),
    .D(_03163_),
    .Q(\rvcpu.dp.pcreg.q[23] ));
 sky130_fd_sc_hd__dfxtp_1 _31706_ (.CLK(clk),
    .D(_03164_),
    .Q(\rvcpu.dp.pcreg.q[24] ));
 sky130_fd_sc_hd__dfxtp_1 _31707_ (.CLK(clk),
    .D(_03165_),
    .Q(\rvcpu.dp.pcreg.q[25] ));
 sky130_fd_sc_hd__dfxtp_1 _31708_ (.CLK(clk),
    .D(_03166_),
    .Q(\rvcpu.dp.pcreg.q[26] ));
 sky130_fd_sc_hd__dfxtp_1 _31709_ (.CLK(clk),
    .D(_03167_),
    .Q(\rvcpu.dp.pcreg.q[27] ));
 sky130_fd_sc_hd__dfxtp_1 _31710_ (.CLK(clk),
    .D(_03168_),
    .Q(\rvcpu.dp.pcreg.q[28] ));
 sky130_fd_sc_hd__dfxtp_1 _31711_ (.CLK(clk),
    .D(_03169_),
    .Q(\rvcpu.dp.pcreg.q[29] ));
 sky130_fd_sc_hd__dfxtp_1 _31712_ (.CLK(clk),
    .D(_03170_),
    .Q(\rvcpu.dp.pcreg.q[30] ));
 sky130_fd_sc_hd__dfxtp_1 _31713_ (.CLK(clk),
    .D(_03171_),
    .Q(\rvcpu.dp.pcreg.q[31] ));
 sky130_fd_sc_hd__dfxtp_1 _31714_ (.CLK(_00996_),
    .D(_03172_),
    .Q(\rvcpu.dp.rf.reg_file_arr[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _31715_ (.CLK(_00997_),
    .D(_03173_),
    .Q(\rvcpu.dp.rf.reg_file_arr[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _31716_ (.CLK(_00998_),
    .D(_03174_),
    .Q(\rvcpu.dp.rf.reg_file_arr[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _31717_ (.CLK(_00999_),
    .D(_03175_),
    .Q(\rvcpu.dp.rf.reg_file_arr[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _31718_ (.CLK(_01000_),
    .D(_03176_),
    .Q(\rvcpu.dp.rf.reg_file_arr[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _31719_ (.CLK(_01001_),
    .D(_03177_),
    .Q(\rvcpu.dp.rf.reg_file_arr[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _31720_ (.CLK(_01002_),
    .D(_03178_),
    .Q(\rvcpu.dp.rf.reg_file_arr[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _31721_ (.CLK(_01003_),
    .D(_03179_),
    .Q(\rvcpu.dp.rf.reg_file_arr[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _31722_ (.CLK(_01004_),
    .D(_03180_),
    .Q(\rvcpu.dp.rf.reg_file_arr[9][8] ));
 sky130_fd_sc_hd__dfxtp_1 _31723_ (.CLK(_01005_),
    .D(_03181_),
    .Q(\rvcpu.dp.rf.reg_file_arr[9][9] ));
 sky130_fd_sc_hd__dfxtp_1 _31724_ (.CLK(_01006_),
    .D(_03182_),
    .Q(\rvcpu.dp.rf.reg_file_arr[9][10] ));
 sky130_fd_sc_hd__dfxtp_1 _31725_ (.CLK(_01007_),
    .D(_03183_),
    .Q(\rvcpu.dp.rf.reg_file_arr[9][11] ));
 sky130_fd_sc_hd__dfxtp_1 _31726_ (.CLK(_01008_),
    .D(_03184_),
    .Q(\rvcpu.dp.rf.reg_file_arr[9][12] ));
 sky130_fd_sc_hd__dfxtp_1 _31727_ (.CLK(_01009_),
    .D(_03185_),
    .Q(\rvcpu.dp.rf.reg_file_arr[9][13] ));
 sky130_fd_sc_hd__dfxtp_1 _31728_ (.CLK(_01010_),
    .D(_03186_),
    .Q(\rvcpu.dp.rf.reg_file_arr[9][14] ));
 sky130_fd_sc_hd__dfxtp_1 _31729_ (.CLK(_01011_),
    .D(_03187_),
    .Q(\rvcpu.dp.rf.reg_file_arr[9][15] ));
 sky130_fd_sc_hd__dfxtp_1 _31730_ (.CLK(_01012_),
    .D(_03188_),
    .Q(\rvcpu.dp.rf.reg_file_arr[9][16] ));
 sky130_fd_sc_hd__dfxtp_1 _31731_ (.CLK(_01013_),
    .D(_03189_),
    .Q(\rvcpu.dp.rf.reg_file_arr[9][17] ));
 sky130_fd_sc_hd__dfxtp_1 _31732_ (.CLK(_01014_),
    .D(_03190_),
    .Q(\rvcpu.dp.rf.reg_file_arr[9][18] ));
 sky130_fd_sc_hd__dfxtp_1 _31733_ (.CLK(_01015_),
    .D(_03191_),
    .Q(\rvcpu.dp.rf.reg_file_arr[9][19] ));
 sky130_fd_sc_hd__dfxtp_1 _31734_ (.CLK(_01016_),
    .D(_03192_),
    .Q(\rvcpu.dp.rf.reg_file_arr[9][20] ));
 sky130_fd_sc_hd__dfxtp_1 _31735_ (.CLK(_01017_),
    .D(_03193_),
    .Q(\rvcpu.dp.rf.reg_file_arr[9][21] ));
 sky130_fd_sc_hd__dfxtp_1 _31736_ (.CLK(_01018_),
    .D(_03194_),
    .Q(\rvcpu.dp.rf.reg_file_arr[9][22] ));
 sky130_fd_sc_hd__dfxtp_1 _31737_ (.CLK(_01019_),
    .D(_03195_),
    .Q(\rvcpu.dp.rf.reg_file_arr[9][23] ));
 sky130_fd_sc_hd__dfxtp_1 _31738_ (.CLK(_01020_),
    .D(_03196_),
    .Q(\rvcpu.dp.rf.reg_file_arr[9][24] ));
 sky130_fd_sc_hd__dfxtp_1 _31739_ (.CLK(_01021_),
    .D(_03197_),
    .Q(\rvcpu.dp.rf.reg_file_arr[9][25] ));
 sky130_fd_sc_hd__dfxtp_1 _31740_ (.CLK(_01022_),
    .D(_03198_),
    .Q(\rvcpu.dp.rf.reg_file_arr[9][26] ));
 sky130_fd_sc_hd__dfxtp_1 _31741_ (.CLK(_01023_),
    .D(_03199_),
    .Q(\rvcpu.dp.rf.reg_file_arr[9][27] ));
 sky130_fd_sc_hd__dfxtp_1 _31742_ (.CLK(_01024_),
    .D(_03200_),
    .Q(\rvcpu.dp.rf.reg_file_arr[9][28] ));
 sky130_fd_sc_hd__dfxtp_1 _31743_ (.CLK(_01025_),
    .D(_03201_),
    .Q(\rvcpu.dp.rf.reg_file_arr[9][29] ));
 sky130_fd_sc_hd__dfxtp_1 _31744_ (.CLK(_01026_),
    .D(_03202_),
    .Q(\rvcpu.dp.rf.reg_file_arr[9][30] ));
 sky130_fd_sc_hd__dfxtp_1 _31745_ (.CLK(_01027_),
    .D(_03203_),
    .Q(\rvcpu.dp.rf.reg_file_arr[9][31] ));
 sky130_fd_sc_hd__dlxtn_1 _31746_ (.D(_04447_),
    .GATE_N(net123),
    .Q(\rvcpu.ALUControl[0] ));
 sky130_fd_sc_hd__dlxtn_1 _31747_ (.D(_04448_),
    .GATE_N(net124),
    .Q(\rvcpu.ALUControl[1] ));
 sky130_fd_sc_hd__dlxtn_1 _31748_ (.D(_04449_),
    .GATE_N(net125),
    .Q(\rvcpu.ALUControl[2] ));
 sky130_fd_sc_hd__dlxtn_1 _31749_ (.D(_04450_),
    .GATE_N(net126),
    .Q(\rvcpu.ALUControl[3] ));
 sky130_fd_sc_hd__dfxtp_1 _31750_ (.CLK(clk),
    .D(_03204_),
    .Q(\datamem.data_ram[45][0] ));
 sky130_fd_sc_hd__dfxtp_1 _31751_ (.CLK(clk),
    .D(_03205_),
    .Q(\datamem.data_ram[45][1] ));
 sky130_fd_sc_hd__dfxtp_1 _31752_ (.CLK(clk),
    .D(_03206_),
    .Q(\datamem.data_ram[45][2] ));
 sky130_fd_sc_hd__dfxtp_1 _31753_ (.CLK(clk),
    .D(_03207_),
    .Q(\datamem.data_ram[45][3] ));
 sky130_fd_sc_hd__dfxtp_1 _31754_ (.CLK(clk),
    .D(_03208_),
    .Q(\datamem.data_ram[45][4] ));
 sky130_fd_sc_hd__dfxtp_1 _31755_ (.CLK(clk),
    .D(_03209_),
    .Q(\datamem.data_ram[45][5] ));
 sky130_fd_sc_hd__dfxtp_1 _31756_ (.CLK(clk),
    .D(_03210_),
    .Q(\datamem.data_ram[45][6] ));
 sky130_fd_sc_hd__dfxtp_1 _31757_ (.CLK(clk),
    .D(_03211_),
    .Q(\datamem.data_ram[45][7] ));
 sky130_fd_sc_hd__dfxtp_2 _31758_ (.CLK(clk),
    .D(_03212_),
    .Q(\rvcpu.dp.plde.ALUSrcE ));
 sky130_fd_sc_hd__dfxtp_1 _31759_ (.CLK(clk),
    .D(_03213_),
    .Q(\datamem.data_ram[18][0] ));
 sky130_fd_sc_hd__dfxtp_1 _31760_ (.CLK(clk),
    .D(_03214_),
    .Q(\datamem.data_ram[18][1] ));
 sky130_fd_sc_hd__dfxtp_1 _31761_ (.CLK(clk),
    .D(_03215_),
    .Q(\datamem.data_ram[18][2] ));
 sky130_fd_sc_hd__dfxtp_1 _31762_ (.CLK(clk),
    .D(_03216_),
    .Q(\datamem.data_ram[18][3] ));
 sky130_fd_sc_hd__dfxtp_1 _31763_ (.CLK(clk),
    .D(_03217_),
    .Q(\datamem.data_ram[18][4] ));
 sky130_fd_sc_hd__dfxtp_1 _31764_ (.CLK(clk),
    .D(_03218_),
    .Q(\datamem.data_ram[18][5] ));
 sky130_fd_sc_hd__dfxtp_1 _31765_ (.CLK(clk),
    .D(_03219_),
    .Q(\datamem.data_ram[18][6] ));
 sky130_fd_sc_hd__dfxtp_1 _31766_ (.CLK(clk),
    .D(_03220_),
    .Q(\datamem.data_ram[18][7] ));
 sky130_fd_sc_hd__dfxtp_1 _31767_ (.CLK(clk),
    .D(_03221_),
    .Q(\datamem.data_ram[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _31768_ (.CLK(clk),
    .D(_03222_),
    .Q(\datamem.data_ram[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _31769_ (.CLK(clk),
    .D(_03223_),
    .Q(\datamem.data_ram[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _31770_ (.CLK(clk),
    .D(_03224_),
    .Q(\datamem.data_ram[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _31771_ (.CLK(clk),
    .D(_03225_),
    .Q(\datamem.data_ram[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _31772_ (.CLK(clk),
    .D(_03226_),
    .Q(\datamem.data_ram[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _31773_ (.CLK(clk),
    .D(_03227_),
    .Q(\datamem.data_ram[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _31774_ (.CLK(clk),
    .D(_03228_),
    .Q(\datamem.data_ram[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _31775_ (.CLK(clk),
    .D(_03229_),
    .Q(\datamem.data_ram[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _31776_ (.CLK(clk),
    .D(_03230_),
    .Q(\datamem.data_ram[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _31777_ (.CLK(clk),
    .D(_03231_),
    .Q(\datamem.data_ram[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _31778_ (.CLK(clk),
    .D(_03232_),
    .Q(\datamem.data_ram[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _31779_ (.CLK(clk),
    .D(_03233_),
    .Q(\datamem.data_ram[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _31780_ (.CLK(clk),
    .D(_03234_),
    .Q(\datamem.data_ram[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _31781_ (.CLK(clk),
    .D(_03235_),
    .Q(\datamem.data_ram[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _31782_ (.CLK(clk),
    .D(_03236_),
    .Q(\datamem.data_ram[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _31783_ (.CLK(clk),
    .D(_03237_),
    .Q(\datamem.data_ram[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _31784_ (.CLK(clk),
    .D(_03238_),
    .Q(\datamem.data_ram[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _31785_ (.CLK(clk),
    .D(_03239_),
    .Q(\datamem.data_ram[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _31786_ (.CLK(clk),
    .D(_03240_),
    .Q(\datamem.data_ram[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _31787_ (.CLK(clk),
    .D(_03241_),
    .Q(\datamem.data_ram[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _31788_ (.CLK(clk),
    .D(_03242_),
    .Q(\datamem.data_ram[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _31789_ (.CLK(clk),
    .D(_03243_),
    .Q(\datamem.data_ram[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _31790_ (.CLK(clk),
    .D(_03244_),
    .Q(\datamem.data_ram[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _31791_ (.CLK(clk),
    .D(_03245_),
    .Q(\datamem.data_ram[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _31792_ (.CLK(clk),
    .D(_03246_),
    .Q(\datamem.data_ram[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _31793_ (.CLK(clk),
    .D(_03247_),
    .Q(\datamem.data_ram[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _31794_ (.CLK(clk),
    .D(_03248_),
    .Q(\datamem.data_ram[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _31795_ (.CLK(clk),
    .D(_03249_),
    .Q(\datamem.data_ram[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _31796_ (.CLK(clk),
    .D(_03250_),
    .Q(\datamem.data_ram[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _31797_ (.CLK(clk),
    .D(_03251_),
    .Q(\datamem.data_ram[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _31798_ (.CLK(clk),
    .D(_03252_),
    .Q(\datamem.data_ram[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _31799_ (.CLK(clk),
    .D(_03253_),
    .Q(\datamem.data_ram[46][0] ));
 sky130_fd_sc_hd__dfxtp_1 _31800_ (.CLK(clk),
    .D(_03254_),
    .Q(\datamem.data_ram[46][1] ));
 sky130_fd_sc_hd__dfxtp_1 _31801_ (.CLK(clk),
    .D(_03255_),
    .Q(\datamem.data_ram[46][2] ));
 sky130_fd_sc_hd__dfxtp_1 _31802_ (.CLK(clk),
    .D(_03256_),
    .Q(\datamem.data_ram[46][3] ));
 sky130_fd_sc_hd__dfxtp_1 _31803_ (.CLK(clk),
    .D(_03257_),
    .Q(\datamem.data_ram[46][4] ));
 sky130_fd_sc_hd__dfxtp_1 _31804_ (.CLK(clk),
    .D(_03258_),
    .Q(\datamem.data_ram[46][5] ));
 sky130_fd_sc_hd__dfxtp_1 _31805_ (.CLK(clk),
    .D(_03259_),
    .Q(\datamem.data_ram[46][6] ));
 sky130_fd_sc_hd__dfxtp_1 _31806_ (.CLK(clk),
    .D(_03260_),
    .Q(\datamem.data_ram[46][7] ));
 sky130_fd_sc_hd__dfxtp_1 _31807_ (.CLK(clk),
    .D(_03261_),
    .Q(\datamem.data_ram[17][0] ));
 sky130_fd_sc_hd__dfxtp_1 _31808_ (.CLK(clk),
    .D(_03262_),
    .Q(\datamem.data_ram[17][1] ));
 sky130_fd_sc_hd__dfxtp_1 _31809_ (.CLK(clk),
    .D(_03263_),
    .Q(\datamem.data_ram[17][2] ));
 sky130_fd_sc_hd__dfxtp_1 _31810_ (.CLK(clk),
    .D(_03264_),
    .Q(\datamem.data_ram[17][3] ));
 sky130_fd_sc_hd__dfxtp_1 _31811_ (.CLK(clk),
    .D(_03265_),
    .Q(\datamem.data_ram[17][4] ));
 sky130_fd_sc_hd__dfxtp_1 _31812_ (.CLK(clk),
    .D(_03266_),
    .Q(\datamem.data_ram[17][5] ));
 sky130_fd_sc_hd__dfxtp_1 _31813_ (.CLK(clk),
    .D(_03267_),
    .Q(\datamem.data_ram[17][6] ));
 sky130_fd_sc_hd__dfxtp_1 _31814_ (.CLK(clk),
    .D(_03268_),
    .Q(\datamem.data_ram[17][7] ));
 sky130_fd_sc_hd__dfxtp_1 _31815_ (.CLK(clk),
    .D(_03269_),
    .Q(\datamem.data_ram[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _31816_ (.CLK(clk),
    .D(_03270_),
    .Q(\datamem.data_ram[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _31817_ (.CLK(clk),
    .D(_03271_),
    .Q(\datamem.data_ram[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _31818_ (.CLK(clk),
    .D(_03272_),
    .Q(\datamem.data_ram[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _31819_ (.CLK(clk),
    .D(_03273_),
    .Q(\datamem.data_ram[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _31820_ (.CLK(clk),
    .D(_03274_),
    .Q(\datamem.data_ram[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _31821_ (.CLK(clk),
    .D(_03275_),
    .Q(\datamem.data_ram[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _31822_ (.CLK(clk),
    .D(_03276_),
    .Q(\datamem.data_ram[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _31823_ (.CLK(clk),
    .D(_03277_),
    .Q(\datamem.data_ram[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 _31824_ (.CLK(clk),
    .D(_03278_),
    .Q(\datamem.data_ram[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 _31825_ (.CLK(clk),
    .D(_03279_),
    .Q(\datamem.data_ram[16][2] ));
 sky130_fd_sc_hd__dfxtp_1 _31826_ (.CLK(clk),
    .D(_03280_),
    .Q(\datamem.data_ram[16][3] ));
 sky130_fd_sc_hd__dfxtp_1 _31827_ (.CLK(clk),
    .D(_03281_),
    .Q(\datamem.data_ram[16][4] ));
 sky130_fd_sc_hd__dfxtp_1 _31828_ (.CLK(clk),
    .D(_03282_),
    .Q(\datamem.data_ram[16][5] ));
 sky130_fd_sc_hd__dfxtp_1 _31829_ (.CLK(clk),
    .D(_03283_),
    .Q(\datamem.data_ram[16][6] ));
 sky130_fd_sc_hd__dfxtp_1 _31830_ (.CLK(clk),
    .D(_03284_),
    .Q(\datamem.data_ram[16][7] ));
 sky130_fd_sc_hd__dfxtp_1 _31831_ (.CLK(clk),
    .D(_03285_),
    .Q(\datamem.data_ram[3][24] ));
 sky130_fd_sc_hd__dfxtp_1 _31832_ (.CLK(clk),
    .D(_03286_),
    .Q(\datamem.data_ram[3][25] ));
 sky130_fd_sc_hd__dfxtp_1 _31833_ (.CLK(clk),
    .D(_03287_),
    .Q(\datamem.data_ram[3][26] ));
 sky130_fd_sc_hd__dfxtp_1 _31834_ (.CLK(clk),
    .D(_03288_),
    .Q(\datamem.data_ram[3][27] ));
 sky130_fd_sc_hd__dfxtp_1 _31835_ (.CLK(clk),
    .D(_03289_),
    .Q(\datamem.data_ram[3][28] ));
 sky130_fd_sc_hd__dfxtp_1 _31836_ (.CLK(clk),
    .D(_03290_),
    .Q(\datamem.data_ram[3][29] ));
 sky130_fd_sc_hd__dfxtp_1 _31837_ (.CLK(clk),
    .D(_03291_),
    .Q(\datamem.data_ram[3][30] ));
 sky130_fd_sc_hd__dfxtp_1 _31838_ (.CLK(clk),
    .D(_03292_),
    .Q(\datamem.data_ram[3][31] ));
 sky130_fd_sc_hd__dfxtp_1 _31839_ (.CLK(clk),
    .D(_03293_),
    .Q(\datamem.data_ram[8][16] ));
 sky130_fd_sc_hd__dfxtp_1 _31840_ (.CLK(clk),
    .D(_03294_),
    .Q(\datamem.data_ram[8][17] ));
 sky130_fd_sc_hd__dfxtp_1 _31841_ (.CLK(clk),
    .D(_03295_),
    .Q(\datamem.data_ram[8][18] ));
 sky130_fd_sc_hd__dfxtp_1 _31842_ (.CLK(clk),
    .D(_03296_),
    .Q(\datamem.data_ram[8][19] ));
 sky130_fd_sc_hd__dfxtp_1 _31843_ (.CLK(clk),
    .D(_03297_),
    .Q(\datamem.data_ram[8][20] ));
 sky130_fd_sc_hd__dfxtp_1 _31844_ (.CLK(clk),
    .D(_03298_),
    .Q(\datamem.data_ram[8][21] ));
 sky130_fd_sc_hd__dfxtp_1 _31845_ (.CLK(clk),
    .D(_03299_),
    .Q(\datamem.data_ram[8][22] ));
 sky130_fd_sc_hd__dfxtp_1 _31846_ (.CLK(clk),
    .D(_03300_),
    .Q(\datamem.data_ram[8][23] ));
 sky130_fd_sc_hd__dfxtp_1 _31847_ (.CLK(clk),
    .D(_03301_),
    .Q(\datamem.data_ram[61][0] ));
 sky130_fd_sc_hd__dfxtp_1 _31848_ (.CLK(clk),
    .D(_03302_),
    .Q(\datamem.data_ram[61][1] ));
 sky130_fd_sc_hd__dfxtp_1 _31849_ (.CLK(clk),
    .D(_03303_),
    .Q(\datamem.data_ram[61][2] ));
 sky130_fd_sc_hd__dfxtp_1 _31850_ (.CLK(clk),
    .D(_03304_),
    .Q(\datamem.data_ram[61][3] ));
 sky130_fd_sc_hd__dfxtp_1 _31851_ (.CLK(clk),
    .D(_03305_),
    .Q(\datamem.data_ram[61][4] ));
 sky130_fd_sc_hd__dfxtp_1 _31852_ (.CLK(clk),
    .D(_03306_),
    .Q(\datamem.data_ram[61][5] ));
 sky130_fd_sc_hd__dfxtp_1 _31853_ (.CLK(clk),
    .D(_03307_),
    .Q(\datamem.data_ram[61][6] ));
 sky130_fd_sc_hd__dfxtp_1 _31854_ (.CLK(clk),
    .D(_03308_),
    .Q(\datamem.data_ram[61][7] ));
 sky130_fd_sc_hd__dfxtp_1 _31855_ (.CLK(clk),
    .D(_03309_),
    .Q(\datamem.data_ram[62][0] ));
 sky130_fd_sc_hd__dfxtp_1 _31856_ (.CLK(clk),
    .D(_03310_),
    .Q(\datamem.data_ram[62][1] ));
 sky130_fd_sc_hd__dfxtp_1 _31857_ (.CLK(clk),
    .D(_03311_),
    .Q(\datamem.data_ram[62][2] ));
 sky130_fd_sc_hd__dfxtp_1 _31858_ (.CLK(clk),
    .D(_03312_),
    .Q(\datamem.data_ram[62][3] ));
 sky130_fd_sc_hd__dfxtp_1 _31859_ (.CLK(clk),
    .D(_03313_),
    .Q(\datamem.data_ram[62][4] ));
 sky130_fd_sc_hd__dfxtp_1 _31860_ (.CLK(clk),
    .D(_03314_),
    .Q(\datamem.data_ram[62][5] ));
 sky130_fd_sc_hd__dfxtp_1 _31861_ (.CLK(clk),
    .D(_03315_),
    .Q(\datamem.data_ram[62][6] ));
 sky130_fd_sc_hd__dfxtp_1 _31862_ (.CLK(clk),
    .D(_03316_),
    .Q(\datamem.data_ram[62][7] ));
 sky130_fd_sc_hd__dfxtp_1 _31863_ (.CLK(clk),
    .D(_03317_),
    .Q(\datamem.data_ram[63][0] ));
 sky130_fd_sc_hd__dfxtp_1 _31864_ (.CLK(clk),
    .D(_03318_),
    .Q(\datamem.data_ram[63][1] ));
 sky130_fd_sc_hd__dfxtp_1 _31865_ (.CLK(clk),
    .D(_03319_),
    .Q(\datamem.data_ram[63][2] ));
 sky130_fd_sc_hd__dfxtp_1 _31866_ (.CLK(clk),
    .D(_03320_),
    .Q(\datamem.data_ram[63][3] ));
 sky130_fd_sc_hd__dfxtp_1 _31867_ (.CLK(clk),
    .D(_03321_),
    .Q(\datamem.data_ram[63][4] ));
 sky130_fd_sc_hd__dfxtp_1 _31868_ (.CLK(clk),
    .D(_03322_),
    .Q(\datamem.data_ram[63][5] ));
 sky130_fd_sc_hd__dfxtp_1 _31869_ (.CLK(clk),
    .D(_03323_),
    .Q(\datamem.data_ram[63][6] ));
 sky130_fd_sc_hd__dfxtp_1 _31870_ (.CLK(clk),
    .D(_03324_),
    .Q(\datamem.data_ram[63][7] ));
 sky130_fd_sc_hd__dfxtp_1 _31871_ (.CLK(clk),
    .D(_03325_),
    .Q(\datamem.data_ram[56][0] ));
 sky130_fd_sc_hd__dfxtp_1 _31872_ (.CLK(clk),
    .D(_03326_),
    .Q(\datamem.data_ram[56][1] ));
 sky130_fd_sc_hd__dfxtp_1 _31873_ (.CLK(clk),
    .D(_03327_),
    .Q(\datamem.data_ram[56][2] ));
 sky130_fd_sc_hd__dfxtp_1 _31874_ (.CLK(clk),
    .D(_03328_),
    .Q(\datamem.data_ram[56][3] ));
 sky130_fd_sc_hd__dfxtp_1 _31875_ (.CLK(clk),
    .D(_03329_),
    .Q(\datamem.data_ram[56][4] ));
 sky130_fd_sc_hd__dfxtp_1 _31876_ (.CLK(clk),
    .D(_03330_),
    .Q(\datamem.data_ram[56][5] ));
 sky130_fd_sc_hd__dfxtp_1 _31877_ (.CLK(clk),
    .D(_03331_),
    .Q(\datamem.data_ram[56][6] ));
 sky130_fd_sc_hd__dfxtp_1 _31878_ (.CLK(clk),
    .D(_03332_),
    .Q(\datamem.data_ram[56][7] ));
 sky130_fd_sc_hd__dfxtp_1 _31879_ (.CLK(clk),
    .D(_03333_),
    .Q(\datamem.data_ram[57][0] ));
 sky130_fd_sc_hd__dfxtp_1 _31880_ (.CLK(clk),
    .D(_03334_),
    .Q(\datamem.data_ram[57][1] ));
 sky130_fd_sc_hd__dfxtp_1 _31881_ (.CLK(clk),
    .D(_03335_),
    .Q(\datamem.data_ram[57][2] ));
 sky130_fd_sc_hd__dfxtp_1 _31882_ (.CLK(clk),
    .D(_03336_),
    .Q(\datamem.data_ram[57][3] ));
 sky130_fd_sc_hd__dfxtp_1 _31883_ (.CLK(clk),
    .D(_03337_),
    .Q(\datamem.data_ram[57][4] ));
 sky130_fd_sc_hd__dfxtp_1 _31884_ (.CLK(clk),
    .D(_03338_),
    .Q(\datamem.data_ram[57][5] ));
 sky130_fd_sc_hd__dfxtp_1 _31885_ (.CLK(clk),
    .D(_03339_),
    .Q(\datamem.data_ram[57][6] ));
 sky130_fd_sc_hd__dfxtp_1 _31886_ (.CLK(clk),
    .D(_03340_),
    .Q(\datamem.data_ram[57][7] ));
 sky130_fd_sc_hd__dfxtp_1 _31887_ (.CLK(clk),
    .D(_03341_),
    .Q(\datamem.data_ram[36][0] ));
 sky130_fd_sc_hd__dfxtp_1 _31888_ (.CLK(clk),
    .D(_03342_),
    .Q(\datamem.data_ram[36][1] ));
 sky130_fd_sc_hd__dfxtp_1 _31889_ (.CLK(clk),
    .D(_03343_),
    .Q(\datamem.data_ram[36][2] ));
 sky130_fd_sc_hd__dfxtp_1 _31890_ (.CLK(clk),
    .D(_03344_),
    .Q(\datamem.data_ram[36][3] ));
 sky130_fd_sc_hd__dfxtp_1 _31891_ (.CLK(clk),
    .D(_03345_),
    .Q(\datamem.data_ram[36][4] ));
 sky130_fd_sc_hd__dfxtp_1 _31892_ (.CLK(clk),
    .D(_03346_),
    .Q(\datamem.data_ram[36][5] ));
 sky130_fd_sc_hd__dfxtp_1 _31893_ (.CLK(clk),
    .D(_03347_),
    .Q(\datamem.data_ram[36][6] ));
 sky130_fd_sc_hd__dfxtp_1 _31894_ (.CLK(clk),
    .D(_03348_),
    .Q(\datamem.data_ram[36][7] ));
 sky130_fd_sc_hd__dlxtn_1 _31895_ (.D(_04415_),
    .GATE_N(net118),
    .Q(\datamem.rd_data_mem[0] ));
 sky130_fd_sc_hd__dlxtn_1 _31896_ (.D(_04426_),
    .GATE_N(net120),
    .Q(\datamem.rd_data_mem[1] ));
 sky130_fd_sc_hd__dlxtn_1 _31897_ (.D(_04437_),
    .GATE_N(net120),
    .Q(\datamem.rd_data_mem[2] ));
 sky130_fd_sc_hd__dlxtn_1 _31898_ (.D(_04440_),
    .GATE_N(net120),
    .Q(\datamem.rd_data_mem[3] ));
 sky130_fd_sc_hd__dlxtn_1 _31899_ (.D(_04441_),
    .GATE_N(net118),
    .Q(\datamem.rd_data_mem[4] ));
 sky130_fd_sc_hd__dlxtn_1 _31900_ (.D(_04442_),
    .GATE_N(net121),
    .Q(\datamem.rd_data_mem[5] ));
 sky130_fd_sc_hd__dlxtn_1 _31901_ (.D(_04443_),
    .GATE_N(net121),
    .Q(\datamem.rd_data_mem[6] ));
 sky130_fd_sc_hd__dlxtn_1 _31902_ (.D(_04444_),
    .GATE_N(net121),
    .Q(\datamem.rd_data_mem[7] ));
 sky130_fd_sc_hd__dlxtn_1 _31903_ (.D(_04445_),
    .GATE_N(net118),
    .Q(\datamem.rd_data_mem[8] ));
 sky130_fd_sc_hd__dlxtn_1 _31904_ (.D(_04446_),
    .GATE_N(net119),
    .Q(\datamem.rd_data_mem[9] ));
 sky130_fd_sc_hd__dlxtn_1 _31905_ (.D(_04416_),
    .GATE_N(net120),
    .Q(\datamem.rd_data_mem[10] ));
 sky130_fd_sc_hd__dlxtn_1 _31906_ (.D(_04417_),
    .GATE_N(net120),
    .Q(\datamem.rd_data_mem[11] ));
 sky130_fd_sc_hd__dlxtn_1 _31907_ (.D(_04418_),
    .GATE_N(net119),
    .Q(\datamem.rd_data_mem[12] ));
 sky130_fd_sc_hd__dlxtn_1 _31908_ (.D(_04419_),
    .GATE_N(net118),
    .Q(\datamem.rd_data_mem[13] ));
 sky130_fd_sc_hd__dlxtn_1 _31909_ (.D(_04420_),
    .GATE_N(net121),
    .Q(\datamem.rd_data_mem[14] ));
 sky130_fd_sc_hd__dlxtn_1 _31910_ (.D(_04421_),
    .GATE_N(net118),
    .Q(\datamem.rd_data_mem[15] ));
 sky130_fd_sc_hd__dlxtn_1 _31911_ (.D(_04422_),
    .GATE_N(net121),
    .Q(\datamem.rd_data_mem[16] ));
 sky130_fd_sc_hd__dlxtn_1 _31912_ (.D(_04423_),
    .GATE_N(net120),
    .Q(\datamem.rd_data_mem[17] ));
 sky130_fd_sc_hd__dlxtn_1 _31913_ (.D(_04424_),
    .GATE_N(net121),
    .Q(\datamem.rd_data_mem[18] ));
 sky130_fd_sc_hd__dlxtn_1 _31914_ (.D(_04425_),
    .GATE_N(net120),
    .Q(\datamem.rd_data_mem[19] ));
 sky130_fd_sc_hd__dlxtn_1 _31915_ (.D(_04427_),
    .GATE_N(net120),
    .Q(\datamem.rd_data_mem[20] ));
 sky130_fd_sc_hd__dlxtn_1 _31916_ (.D(_04428_),
    .GATE_N(net120),
    .Q(\datamem.rd_data_mem[21] ));
 sky130_fd_sc_hd__dlxtn_1 _31917_ (.D(_04429_),
    .GATE_N(net120),
    .Q(\datamem.rd_data_mem[22] ));
 sky130_fd_sc_hd__dlxtn_1 _31918_ (.D(_04430_),
    .GATE_N(net119),
    .Q(\datamem.rd_data_mem[23] ));
 sky130_fd_sc_hd__dlxtn_1 _31919_ (.D(_04431_),
    .GATE_N(net119),
    .Q(\datamem.rd_data_mem[24] ));
 sky130_fd_sc_hd__dlxtn_1 _31920_ (.D(_04432_),
    .GATE_N(net119),
    .Q(\datamem.rd_data_mem[25] ));
 sky130_fd_sc_hd__dlxtn_1 _31921_ (.D(_04433_),
    .GATE_N(net119),
    .Q(\datamem.rd_data_mem[26] ));
 sky130_fd_sc_hd__dlxtn_1 _31922_ (.D(_04434_),
    .GATE_N(net118),
    .Q(\datamem.rd_data_mem[27] ));
 sky130_fd_sc_hd__dlxtn_1 _31923_ (.D(_04435_),
    .GATE_N(net118),
    .Q(\datamem.rd_data_mem[28] ));
 sky130_fd_sc_hd__dlxtn_1 _31924_ (.D(_04436_),
    .GATE_N(net118),
    .Q(\datamem.rd_data_mem[29] ));
 sky130_fd_sc_hd__dlxtn_1 _31925_ (.D(_04438_),
    .GATE_N(net118),
    .Q(\datamem.rd_data_mem[30] ));
 sky130_fd_sc_hd__dlxtn_1 _31926_ (.D(_04439_),
    .GATE_N(net119),
    .Q(\datamem.rd_data_mem[31] ));
 sky130_fd_sc_hd__dfxtp_1 _31927_ (.CLK(clk),
    .D(_03349_),
    .Q(\datamem.data_ram[60][0] ));
 sky130_fd_sc_hd__dfxtp_1 _31928_ (.CLK(clk),
    .D(_03350_),
    .Q(\datamem.data_ram[60][1] ));
 sky130_fd_sc_hd__dfxtp_1 _31929_ (.CLK(clk),
    .D(_03351_),
    .Q(\datamem.data_ram[60][2] ));
 sky130_fd_sc_hd__dfxtp_1 _31930_ (.CLK(clk),
    .D(_03352_),
    .Q(\datamem.data_ram[60][3] ));
 sky130_fd_sc_hd__dfxtp_1 _31931_ (.CLK(clk),
    .D(_03353_),
    .Q(\datamem.data_ram[60][4] ));
 sky130_fd_sc_hd__dfxtp_1 _31932_ (.CLK(clk),
    .D(_03354_),
    .Q(\datamem.data_ram[60][5] ));
 sky130_fd_sc_hd__dfxtp_1 _31933_ (.CLK(clk),
    .D(_03355_),
    .Q(\datamem.data_ram[60][6] ));
 sky130_fd_sc_hd__dfxtp_1 _31934_ (.CLK(clk),
    .D(_03356_),
    .Q(\datamem.data_ram[60][7] ));
 sky130_fd_sc_hd__dfxtp_1 _31935_ (.CLK(clk),
    .D(_03357_),
    .Q(\datamem.data_ram[59][0] ));
 sky130_fd_sc_hd__dfxtp_1 _31936_ (.CLK(clk),
    .D(_03358_),
    .Q(\datamem.data_ram[59][1] ));
 sky130_fd_sc_hd__dfxtp_1 _31937_ (.CLK(clk),
    .D(_03359_),
    .Q(\datamem.data_ram[59][2] ));
 sky130_fd_sc_hd__dfxtp_1 _31938_ (.CLK(clk),
    .D(_03360_),
    .Q(\datamem.data_ram[59][3] ));
 sky130_fd_sc_hd__dfxtp_1 _31939_ (.CLK(clk),
    .D(_03361_),
    .Q(\datamem.data_ram[59][4] ));
 sky130_fd_sc_hd__dfxtp_1 _31940_ (.CLK(clk),
    .D(_03362_),
    .Q(\datamem.data_ram[59][5] ));
 sky130_fd_sc_hd__dfxtp_1 _31941_ (.CLK(clk),
    .D(_03363_),
    .Q(\datamem.data_ram[59][6] ));
 sky130_fd_sc_hd__dfxtp_1 _31942_ (.CLK(clk),
    .D(_03364_),
    .Q(\datamem.data_ram[59][7] ));
 sky130_fd_sc_hd__dfxtp_1 _31943_ (.CLK(clk),
    .D(_03365_),
    .Q(\datamem.data_ram[32][0] ));
 sky130_fd_sc_hd__dfxtp_1 _31944_ (.CLK(clk),
    .D(_03366_),
    .Q(\datamem.data_ram[32][1] ));
 sky130_fd_sc_hd__dfxtp_1 _31945_ (.CLK(clk),
    .D(_03367_),
    .Q(\datamem.data_ram[32][2] ));
 sky130_fd_sc_hd__dfxtp_1 _31946_ (.CLK(clk),
    .D(_03368_),
    .Q(\datamem.data_ram[32][3] ));
 sky130_fd_sc_hd__dfxtp_1 _31947_ (.CLK(clk),
    .D(_03369_),
    .Q(\datamem.data_ram[32][4] ));
 sky130_fd_sc_hd__dfxtp_1 _31948_ (.CLK(clk),
    .D(_03370_),
    .Q(\datamem.data_ram[32][5] ));
 sky130_fd_sc_hd__dfxtp_1 _31949_ (.CLK(clk),
    .D(_03371_),
    .Q(\datamem.data_ram[32][6] ));
 sky130_fd_sc_hd__dfxtp_1 _31950_ (.CLK(clk),
    .D(_03372_),
    .Q(\datamem.data_ram[32][7] ));
 sky130_fd_sc_hd__dfxtp_1 _31951_ (.CLK(clk),
    .D(_03373_),
    .Q(\datamem.data_ram[55][0] ));
 sky130_fd_sc_hd__dfxtp_1 _31952_ (.CLK(clk),
    .D(_03374_),
    .Q(\datamem.data_ram[55][1] ));
 sky130_fd_sc_hd__dfxtp_1 _31953_ (.CLK(clk),
    .D(_03375_),
    .Q(\datamem.data_ram[55][2] ));
 sky130_fd_sc_hd__dfxtp_1 _31954_ (.CLK(clk),
    .D(_03376_),
    .Q(\datamem.data_ram[55][3] ));
 sky130_fd_sc_hd__dfxtp_1 _31955_ (.CLK(clk),
    .D(_03377_),
    .Q(\datamem.data_ram[55][4] ));
 sky130_fd_sc_hd__dfxtp_1 _31956_ (.CLK(clk),
    .D(_03378_),
    .Q(\datamem.data_ram[55][5] ));
 sky130_fd_sc_hd__dfxtp_1 _31957_ (.CLK(clk),
    .D(_03379_),
    .Q(\datamem.data_ram[55][6] ));
 sky130_fd_sc_hd__dfxtp_1 _31958_ (.CLK(clk),
    .D(_03380_),
    .Q(\datamem.data_ram[55][7] ));
 sky130_fd_sc_hd__dfxtp_1 _31959_ (.CLK(clk),
    .D(_03381_),
    .Q(\datamem.data_ram[28][0] ));
 sky130_fd_sc_hd__dfxtp_1 _31960_ (.CLK(clk),
    .D(_03382_),
    .Q(\datamem.data_ram[28][1] ));
 sky130_fd_sc_hd__dfxtp_1 _31961_ (.CLK(clk),
    .D(_03383_),
    .Q(\datamem.data_ram[28][2] ));
 sky130_fd_sc_hd__dfxtp_1 _31962_ (.CLK(clk),
    .D(_03384_),
    .Q(\datamem.data_ram[28][3] ));
 sky130_fd_sc_hd__dfxtp_1 _31963_ (.CLK(clk),
    .D(_03385_),
    .Q(\datamem.data_ram[28][4] ));
 sky130_fd_sc_hd__dfxtp_1 _31964_ (.CLK(clk),
    .D(_03386_),
    .Q(\datamem.data_ram[28][5] ));
 sky130_fd_sc_hd__dfxtp_1 _31965_ (.CLK(clk),
    .D(_03387_),
    .Q(\datamem.data_ram[28][6] ));
 sky130_fd_sc_hd__dfxtp_1 _31966_ (.CLK(clk),
    .D(_03388_),
    .Q(\datamem.data_ram[28][7] ));
 sky130_fd_sc_hd__dfxtp_1 _31967_ (.CLK(clk),
    .D(_03389_),
    .Q(\datamem.data_ram[54][0] ));
 sky130_fd_sc_hd__dfxtp_1 _31968_ (.CLK(clk),
    .D(_03390_),
    .Q(\datamem.data_ram[54][1] ));
 sky130_fd_sc_hd__dfxtp_1 _31969_ (.CLK(clk),
    .D(_03391_),
    .Q(\datamem.data_ram[54][2] ));
 sky130_fd_sc_hd__dfxtp_1 _31970_ (.CLK(clk),
    .D(_03392_),
    .Q(\datamem.data_ram[54][3] ));
 sky130_fd_sc_hd__dfxtp_1 _31971_ (.CLK(clk),
    .D(_03393_),
    .Q(\datamem.data_ram[54][4] ));
 sky130_fd_sc_hd__dfxtp_1 _31972_ (.CLK(clk),
    .D(_03394_),
    .Q(\datamem.data_ram[54][5] ));
 sky130_fd_sc_hd__dfxtp_1 _31973_ (.CLK(clk),
    .D(_03395_),
    .Q(\datamem.data_ram[54][6] ));
 sky130_fd_sc_hd__dfxtp_1 _31974_ (.CLK(clk),
    .D(_03396_),
    .Q(\datamem.data_ram[54][7] ));
 sky130_fd_sc_hd__dfxtp_1 _31975_ (.CLK(clk),
    .D(_03397_),
    .Q(\datamem.data_ram[53][16] ));
 sky130_fd_sc_hd__dfxtp_1 _31976_ (.CLK(clk),
    .D(_03398_),
    .Q(\datamem.data_ram[53][17] ));
 sky130_fd_sc_hd__dfxtp_1 _31977_ (.CLK(clk),
    .D(_03399_),
    .Q(\datamem.data_ram[53][18] ));
 sky130_fd_sc_hd__dfxtp_1 _31978_ (.CLK(clk),
    .D(_03400_),
    .Q(\datamem.data_ram[53][19] ));
 sky130_fd_sc_hd__dfxtp_1 _31979_ (.CLK(clk),
    .D(_03401_),
    .Q(\datamem.data_ram[53][20] ));
 sky130_fd_sc_hd__dfxtp_1 _31980_ (.CLK(clk),
    .D(_03402_),
    .Q(\datamem.data_ram[53][21] ));
 sky130_fd_sc_hd__dfxtp_1 _31981_ (.CLK(clk),
    .D(_03403_),
    .Q(\datamem.data_ram[53][22] ));
 sky130_fd_sc_hd__dfxtp_1 _31982_ (.CLK(clk),
    .D(_03404_),
    .Q(\datamem.data_ram[53][23] ));
 sky130_fd_sc_hd__dfxtp_1 _31983_ (.CLK(clk),
    .D(_03405_),
    .Q(\datamem.data_ram[37][0] ));
 sky130_fd_sc_hd__dfxtp_1 _31984_ (.CLK(clk),
    .D(_03406_),
    .Q(\datamem.data_ram[37][1] ));
 sky130_fd_sc_hd__dfxtp_1 _31985_ (.CLK(clk),
    .D(_03407_),
    .Q(\datamem.data_ram[37][2] ));
 sky130_fd_sc_hd__dfxtp_1 _31986_ (.CLK(clk),
    .D(_03408_),
    .Q(\datamem.data_ram[37][3] ));
 sky130_fd_sc_hd__dfxtp_1 _31987_ (.CLK(clk),
    .D(_03409_),
    .Q(\datamem.data_ram[37][4] ));
 sky130_fd_sc_hd__dfxtp_1 _31988_ (.CLK(clk),
    .D(_03410_),
    .Q(\datamem.data_ram[37][5] ));
 sky130_fd_sc_hd__dfxtp_1 _31989_ (.CLK(clk),
    .D(_03411_),
    .Q(\datamem.data_ram[37][6] ));
 sky130_fd_sc_hd__dfxtp_1 _31990_ (.CLK(clk),
    .D(_03412_),
    .Q(\datamem.data_ram[37][7] ));
 sky130_fd_sc_hd__dfxtp_1 _31991_ (.CLK(clk),
    .D(_03413_),
    .Q(\datamem.data_ram[31][0] ));
 sky130_fd_sc_hd__dfxtp_1 _31992_ (.CLK(clk),
    .D(_03414_),
    .Q(\datamem.data_ram[31][1] ));
 sky130_fd_sc_hd__dfxtp_1 _31993_ (.CLK(clk),
    .D(_03415_),
    .Q(\datamem.data_ram[31][2] ));
 sky130_fd_sc_hd__dfxtp_1 _31994_ (.CLK(clk),
    .D(_03416_),
    .Q(\datamem.data_ram[31][3] ));
 sky130_fd_sc_hd__dfxtp_1 _31995_ (.CLK(clk),
    .D(_03417_),
    .Q(\datamem.data_ram[31][4] ));
 sky130_fd_sc_hd__dfxtp_1 _31996_ (.CLK(clk),
    .D(_03418_),
    .Q(\datamem.data_ram[31][5] ));
 sky130_fd_sc_hd__dfxtp_1 _31997_ (.CLK(clk),
    .D(_03419_),
    .Q(\datamem.data_ram[31][6] ));
 sky130_fd_sc_hd__dfxtp_1 _31998_ (.CLK(clk),
    .D(_03420_),
    .Q(\datamem.data_ram[31][7] ));
 sky130_fd_sc_hd__dfxtp_1 _31999_ (.CLK(clk),
    .D(_03421_),
    .Q(\datamem.data_ram[52][0] ));
 sky130_fd_sc_hd__dfxtp_1 _32000_ (.CLK(clk),
    .D(_03422_),
    .Q(\datamem.data_ram[52][1] ));
 sky130_fd_sc_hd__dfxtp_1 _32001_ (.CLK(clk),
    .D(_03423_),
    .Q(\datamem.data_ram[52][2] ));
 sky130_fd_sc_hd__dfxtp_2 _32002_ (.CLK(clk),
    .D(_03424_),
    .Q(\datamem.data_ram[52][3] ));
 sky130_fd_sc_hd__dfxtp_1 _32003_ (.CLK(clk),
    .D(_03425_),
    .Q(\datamem.data_ram[52][4] ));
 sky130_fd_sc_hd__dfxtp_1 _32004_ (.CLK(clk),
    .D(_03426_),
    .Q(\datamem.data_ram[52][5] ));
 sky130_fd_sc_hd__dfxtp_1 _32005_ (.CLK(clk),
    .D(_03427_),
    .Q(\datamem.data_ram[52][6] ));
 sky130_fd_sc_hd__dfxtp_2 _32006_ (.CLK(clk),
    .D(_03428_),
    .Q(\datamem.data_ram[52][7] ));
 sky130_fd_sc_hd__dfxtp_1 _32007_ (.CLK(clk),
    .D(_03429_),
    .Q(\datamem.data_ram[27][0] ));
 sky130_fd_sc_hd__dfxtp_1 _32008_ (.CLK(clk),
    .D(_03430_),
    .Q(\datamem.data_ram[27][1] ));
 sky130_fd_sc_hd__dfxtp_1 _32009_ (.CLK(clk),
    .D(_03431_),
    .Q(\datamem.data_ram[27][2] ));
 sky130_fd_sc_hd__dfxtp_1 _32010_ (.CLK(clk),
    .D(_03432_),
    .Q(\datamem.data_ram[27][3] ));
 sky130_fd_sc_hd__dfxtp_1 _32011_ (.CLK(clk),
    .D(_03433_),
    .Q(\datamem.data_ram[27][4] ));
 sky130_fd_sc_hd__dfxtp_1 _32012_ (.CLK(clk),
    .D(_03434_),
    .Q(\datamem.data_ram[27][5] ));
 sky130_fd_sc_hd__dfxtp_1 _32013_ (.CLK(clk),
    .D(_03435_),
    .Q(\datamem.data_ram[27][6] ));
 sky130_fd_sc_hd__dfxtp_1 _32014_ (.CLK(clk),
    .D(_03436_),
    .Q(\datamem.data_ram[27][7] ));
 sky130_fd_sc_hd__dfxtp_1 _32015_ (.CLK(clk),
    .D(_03437_),
    .Q(\rvcpu.dp.pcreg.q[0] ));
 sky130_fd_sc_hd__dfxtp_1 _32016_ (.CLK(clk),
    .D(_03438_),
    .Q(\rvcpu.dp.pcreg.q[1] ));
 sky130_fd_sc_hd__dfxtp_1 _32017_ (.CLK(clk),
    .D(_03439_),
    .Q(\datamem.data_ram[51][0] ));
 sky130_fd_sc_hd__dfxtp_1 _32018_ (.CLK(clk),
    .D(_03440_),
    .Q(\datamem.data_ram[51][1] ));
 sky130_fd_sc_hd__dfxtp_1 _32019_ (.CLK(clk),
    .D(_03441_),
    .Q(\datamem.data_ram[51][2] ));
 sky130_fd_sc_hd__dfxtp_1 _32020_ (.CLK(clk),
    .D(_03442_),
    .Q(\datamem.data_ram[51][3] ));
 sky130_fd_sc_hd__dfxtp_1 _32021_ (.CLK(clk),
    .D(_03443_),
    .Q(\datamem.data_ram[51][4] ));
 sky130_fd_sc_hd__dfxtp_1 _32022_ (.CLK(clk),
    .D(_03444_),
    .Q(\datamem.data_ram[51][5] ));
 sky130_fd_sc_hd__dfxtp_1 _32023_ (.CLK(clk),
    .D(_03445_),
    .Q(\datamem.data_ram[51][6] ));
 sky130_fd_sc_hd__dfxtp_1 _32024_ (.CLK(clk),
    .D(_03446_),
    .Q(\datamem.data_ram[51][7] ));
 sky130_fd_sc_hd__dfxtp_1 _32025_ (.CLK(clk),
    .D(_03447_),
    .Q(\datamem.data_ram[26][0] ));
 sky130_fd_sc_hd__dfxtp_1 _32026_ (.CLK(clk),
    .D(_03448_),
    .Q(\datamem.data_ram[26][1] ));
 sky130_fd_sc_hd__dfxtp_1 _32027_ (.CLK(clk),
    .D(_03449_),
    .Q(\datamem.data_ram[26][2] ));
 sky130_fd_sc_hd__dfxtp_1 _32028_ (.CLK(clk),
    .D(_03450_),
    .Q(\datamem.data_ram[26][3] ));
 sky130_fd_sc_hd__dfxtp_1 _32029_ (.CLK(clk),
    .D(_03451_),
    .Q(\datamem.data_ram[26][4] ));
 sky130_fd_sc_hd__dfxtp_1 _32030_ (.CLK(clk),
    .D(_03452_),
    .Q(\datamem.data_ram[26][5] ));
 sky130_fd_sc_hd__dfxtp_1 _32031_ (.CLK(clk),
    .D(_03453_),
    .Q(\datamem.data_ram[26][6] ));
 sky130_fd_sc_hd__dfxtp_1 _32032_ (.CLK(clk),
    .D(_03454_),
    .Q(\datamem.data_ram[26][7] ));
 sky130_fd_sc_hd__dfxtp_1 _32033_ (.CLK(clk),
    .D(_03455_),
    .Q(\datamem.data_ram[50][0] ));
 sky130_fd_sc_hd__dfxtp_1 _32034_ (.CLK(clk),
    .D(_03456_),
    .Q(\datamem.data_ram[50][1] ));
 sky130_fd_sc_hd__dfxtp_1 _32035_ (.CLK(clk),
    .D(_03457_),
    .Q(\datamem.data_ram[50][2] ));
 sky130_fd_sc_hd__dfxtp_1 _32036_ (.CLK(clk),
    .D(_03458_),
    .Q(\datamem.data_ram[50][3] ));
 sky130_fd_sc_hd__dfxtp_1 _32037_ (.CLK(clk),
    .D(_03459_),
    .Q(\datamem.data_ram[50][4] ));
 sky130_fd_sc_hd__dfxtp_1 _32038_ (.CLK(clk),
    .D(_03460_),
    .Q(\datamem.data_ram[50][5] ));
 sky130_fd_sc_hd__dfxtp_1 _32039_ (.CLK(clk),
    .D(_03461_),
    .Q(\datamem.data_ram[50][6] ));
 sky130_fd_sc_hd__dfxtp_1 _32040_ (.CLK(clk),
    .D(_03462_),
    .Q(\datamem.data_ram[50][7] ));
 sky130_fd_sc_hd__dfxtp_1 _32041_ (.CLK(clk),
    .D(_03463_),
    .Q(\datamem.data_ram[49][0] ));
 sky130_fd_sc_hd__dfxtp_1 _32042_ (.CLK(clk),
    .D(_03464_),
    .Q(\datamem.data_ram[49][1] ));
 sky130_fd_sc_hd__dfxtp_1 _32043_ (.CLK(clk),
    .D(_03465_),
    .Q(\datamem.data_ram[49][2] ));
 sky130_fd_sc_hd__dfxtp_1 _32044_ (.CLK(clk),
    .D(_03466_),
    .Q(\datamem.data_ram[49][3] ));
 sky130_fd_sc_hd__dfxtp_1 _32045_ (.CLK(clk),
    .D(_03467_),
    .Q(\datamem.data_ram[49][4] ));
 sky130_fd_sc_hd__dfxtp_1 _32046_ (.CLK(clk),
    .D(_03468_),
    .Q(\datamem.data_ram[49][5] ));
 sky130_fd_sc_hd__dfxtp_1 _32047_ (.CLK(clk),
    .D(_03469_),
    .Q(\datamem.data_ram[49][6] ));
 sky130_fd_sc_hd__dfxtp_1 _32048_ (.CLK(clk),
    .D(_03470_),
    .Q(\datamem.data_ram[49][7] ));
 sky130_fd_sc_hd__dfxtp_1 _32049_ (.CLK(clk),
    .D(_03471_),
    .Q(\datamem.data_ram[30][0] ));
 sky130_fd_sc_hd__dfxtp_1 _32050_ (.CLK(clk),
    .D(_03472_),
    .Q(\datamem.data_ram[30][1] ));
 sky130_fd_sc_hd__dfxtp_1 _32051_ (.CLK(clk),
    .D(_03473_),
    .Q(\datamem.data_ram[30][2] ));
 sky130_fd_sc_hd__dfxtp_1 _32052_ (.CLK(clk),
    .D(_03474_),
    .Q(\datamem.data_ram[30][3] ));
 sky130_fd_sc_hd__dfxtp_1 _32053_ (.CLK(clk),
    .D(_03475_),
    .Q(\datamem.data_ram[30][4] ));
 sky130_fd_sc_hd__dfxtp_1 _32054_ (.CLK(clk),
    .D(_03476_),
    .Q(\datamem.data_ram[30][5] ));
 sky130_fd_sc_hd__dfxtp_1 _32055_ (.CLK(clk),
    .D(_03477_),
    .Q(\datamem.data_ram[30][6] ));
 sky130_fd_sc_hd__dfxtp_1 _32056_ (.CLK(clk),
    .D(_03478_),
    .Q(\datamem.data_ram[30][7] ));
 sky130_fd_sc_hd__dfxtp_1 _32057_ (.CLK(clk),
    .D(_03479_),
    .Q(\datamem.data_ram[48][0] ));
 sky130_fd_sc_hd__dfxtp_1 _32058_ (.CLK(clk),
    .D(_03480_),
    .Q(\datamem.data_ram[48][1] ));
 sky130_fd_sc_hd__dfxtp_1 _32059_ (.CLK(clk),
    .D(_03481_),
    .Q(\datamem.data_ram[48][2] ));
 sky130_fd_sc_hd__dfxtp_1 _32060_ (.CLK(clk),
    .D(_03482_),
    .Q(\datamem.data_ram[48][3] ));
 sky130_fd_sc_hd__dfxtp_1 _32061_ (.CLK(clk),
    .D(_03483_),
    .Q(\datamem.data_ram[48][4] ));
 sky130_fd_sc_hd__dfxtp_1 _32062_ (.CLK(clk),
    .D(_03484_),
    .Q(\datamem.data_ram[48][5] ));
 sky130_fd_sc_hd__dfxtp_1 _32063_ (.CLK(clk),
    .D(_03485_),
    .Q(\datamem.data_ram[48][6] ));
 sky130_fd_sc_hd__dfxtp_1 _32064_ (.CLK(clk),
    .D(_03486_),
    .Q(\datamem.data_ram[48][7] ));
 sky130_fd_sc_hd__dfxtp_1 _32065_ (.CLK(clk),
    .D(_03487_),
    .Q(\datamem.data_ram[29][0] ));
 sky130_fd_sc_hd__dfxtp_1 _32066_ (.CLK(clk),
    .D(_03488_),
    .Q(\datamem.data_ram[29][1] ));
 sky130_fd_sc_hd__dfxtp_1 _32067_ (.CLK(clk),
    .D(_03489_),
    .Q(\datamem.data_ram[29][2] ));
 sky130_fd_sc_hd__dfxtp_1 _32068_ (.CLK(clk),
    .D(_03490_),
    .Q(\datamem.data_ram[29][3] ));
 sky130_fd_sc_hd__dfxtp_1 _32069_ (.CLK(clk),
    .D(_03491_),
    .Q(\datamem.data_ram[29][4] ));
 sky130_fd_sc_hd__dfxtp_1 _32070_ (.CLK(clk),
    .D(_03492_),
    .Q(\datamem.data_ram[29][5] ));
 sky130_fd_sc_hd__dfxtp_1 _32071_ (.CLK(clk),
    .D(_03493_),
    .Q(\datamem.data_ram[29][6] ));
 sky130_fd_sc_hd__dfxtp_1 _32072_ (.CLK(clk),
    .D(_03494_),
    .Q(\datamem.data_ram[29][7] ));
 sky130_fd_sc_hd__dfxtp_1 _32073_ (.CLK(clk),
    .D(_03495_),
    .Q(\datamem.data_ram[33][0] ));
 sky130_fd_sc_hd__dfxtp_1 _32074_ (.CLK(clk),
    .D(_03496_),
    .Q(\datamem.data_ram[33][1] ));
 sky130_fd_sc_hd__dfxtp_1 _32075_ (.CLK(clk),
    .D(_03497_),
    .Q(\datamem.data_ram[33][2] ));
 sky130_fd_sc_hd__dfxtp_1 _32076_ (.CLK(clk),
    .D(_03498_),
    .Q(\datamem.data_ram[33][3] ));
 sky130_fd_sc_hd__dfxtp_1 _32077_ (.CLK(clk),
    .D(_03499_),
    .Q(\datamem.data_ram[33][4] ));
 sky130_fd_sc_hd__dfxtp_1 _32078_ (.CLK(clk),
    .D(_03500_),
    .Q(\datamem.data_ram[33][5] ));
 sky130_fd_sc_hd__dfxtp_1 _32079_ (.CLK(clk),
    .D(_03501_),
    .Q(\datamem.data_ram[33][6] ));
 sky130_fd_sc_hd__dfxtp_1 _32080_ (.CLK(clk),
    .D(_03502_),
    .Q(\datamem.data_ram[33][7] ));
 sky130_fd_sc_hd__dfxtp_1 _32081_ (.CLK(clk),
    .D(_03503_),
    .Q(\datamem.data_ram[47][0] ));
 sky130_fd_sc_hd__dfxtp_1 _32082_ (.CLK(clk),
    .D(_03504_),
    .Q(\datamem.data_ram[47][1] ));
 sky130_fd_sc_hd__dfxtp_1 _32083_ (.CLK(clk),
    .D(_03505_),
    .Q(\datamem.data_ram[47][2] ));
 sky130_fd_sc_hd__dfxtp_1 _32084_ (.CLK(clk),
    .D(_03506_),
    .Q(\datamem.data_ram[47][3] ));
 sky130_fd_sc_hd__dfxtp_1 _32085_ (.CLK(clk),
    .D(_03507_),
    .Q(\datamem.data_ram[47][4] ));
 sky130_fd_sc_hd__dfxtp_1 _32086_ (.CLK(clk),
    .D(_03508_),
    .Q(\datamem.data_ram[47][5] ));
 sky130_fd_sc_hd__dfxtp_1 _32087_ (.CLK(clk),
    .D(_03509_),
    .Q(\datamem.data_ram[47][6] ));
 sky130_fd_sc_hd__dfxtp_1 _32088_ (.CLK(clk),
    .D(_03510_),
    .Q(\datamem.data_ram[47][7] ));
 sky130_fd_sc_hd__dfxtp_1 _32089_ (.CLK(clk),
    .D(_03511_),
    .Q(\datamem.data_ram[8][24] ));
 sky130_fd_sc_hd__dfxtp_1 _32090_ (.CLK(clk),
    .D(_03512_),
    .Q(\datamem.data_ram[8][25] ));
 sky130_fd_sc_hd__dfxtp_1 _32091_ (.CLK(clk),
    .D(_03513_),
    .Q(\datamem.data_ram[8][26] ));
 sky130_fd_sc_hd__dfxtp_1 _32092_ (.CLK(clk),
    .D(_03514_),
    .Q(\datamem.data_ram[8][27] ));
 sky130_fd_sc_hd__dfxtp_1 _32093_ (.CLK(clk),
    .D(_03515_),
    .Q(\datamem.data_ram[8][28] ));
 sky130_fd_sc_hd__dfxtp_1 _32094_ (.CLK(clk),
    .D(_03516_),
    .Q(\datamem.data_ram[8][29] ));
 sky130_fd_sc_hd__dfxtp_1 _32095_ (.CLK(clk),
    .D(_03517_),
    .Q(\datamem.data_ram[8][30] ));
 sky130_fd_sc_hd__dfxtp_1 _32096_ (.CLK(clk),
    .D(_03518_),
    .Q(\datamem.data_ram[8][31] ));
 sky130_fd_sc_hd__dfxtp_1 _32097_ (.CLK(clk),
    .D(_03519_),
    .Q(\datamem.data_ram[23][0] ));
 sky130_fd_sc_hd__dfxtp_1 _32098_ (.CLK(clk),
    .D(_03520_),
    .Q(\datamem.data_ram[23][1] ));
 sky130_fd_sc_hd__dfxtp_1 _32099_ (.CLK(clk),
    .D(_03521_),
    .Q(\datamem.data_ram[23][2] ));
 sky130_fd_sc_hd__dfxtp_1 _32100_ (.CLK(clk),
    .D(_03522_),
    .Q(\datamem.data_ram[23][3] ));
 sky130_fd_sc_hd__dfxtp_1 _32101_ (.CLK(clk),
    .D(_03523_),
    .Q(\datamem.data_ram[23][4] ));
 sky130_fd_sc_hd__dfxtp_1 _32102_ (.CLK(clk),
    .D(_03524_),
    .Q(\datamem.data_ram[23][5] ));
 sky130_fd_sc_hd__dfxtp_1 _32103_ (.CLK(clk),
    .D(_03525_),
    .Q(\datamem.data_ram[23][6] ));
 sky130_fd_sc_hd__dfxtp_1 _32104_ (.CLK(clk),
    .D(_03526_),
    .Q(\datamem.data_ram[23][7] ));
 sky130_fd_sc_hd__dfxtp_1 _32105_ (.CLK(clk),
    .D(_03527_),
    .Q(\datamem.data_ram[58][0] ));
 sky130_fd_sc_hd__dfxtp_1 _32106_ (.CLK(clk),
    .D(_03528_),
    .Q(\datamem.data_ram[58][1] ));
 sky130_fd_sc_hd__dfxtp_1 _32107_ (.CLK(clk),
    .D(_03529_),
    .Q(\datamem.data_ram[58][2] ));
 sky130_fd_sc_hd__dfxtp_1 _32108_ (.CLK(clk),
    .D(_03530_),
    .Q(\datamem.data_ram[58][3] ));
 sky130_fd_sc_hd__dfxtp_1 _32109_ (.CLK(clk),
    .D(_03531_),
    .Q(\datamem.data_ram[58][4] ));
 sky130_fd_sc_hd__dfxtp_1 _32110_ (.CLK(clk),
    .D(_03532_),
    .Q(\datamem.data_ram[58][5] ));
 sky130_fd_sc_hd__dfxtp_1 _32111_ (.CLK(clk),
    .D(_03533_),
    .Q(\datamem.data_ram[58][6] ));
 sky130_fd_sc_hd__dfxtp_1 _32112_ (.CLK(clk),
    .D(_03534_),
    .Q(\datamem.data_ram[58][7] ));
 sky130_fd_sc_hd__dfxtp_1 _32113_ (.CLK(clk),
    .D(_03535_),
    .Q(\datamem.data_ram[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _32114_ (.CLK(clk),
    .D(_03536_),
    .Q(\datamem.data_ram[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _32115_ (.CLK(clk),
    .D(_03537_),
    .Q(\datamem.data_ram[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _32116_ (.CLK(clk),
    .D(_03538_),
    .Q(\datamem.data_ram[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _32117_ (.CLK(clk),
    .D(_03539_),
    .Q(\datamem.data_ram[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _32118_ (.CLK(clk),
    .D(_03540_),
    .Q(\datamem.data_ram[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _32119_ (.CLK(clk),
    .D(_03541_),
    .Q(\datamem.data_ram[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _32120_ (.CLK(clk),
    .D(_03542_),
    .Q(\datamem.data_ram[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _32121_ (.CLK(clk),
    .D(_03543_),
    .Q(\datamem.data_ram[7][24] ));
 sky130_fd_sc_hd__dfxtp_1 _32122_ (.CLK(clk),
    .D(_03544_),
    .Q(\datamem.data_ram[7][25] ));
 sky130_fd_sc_hd__dfxtp_1 _32123_ (.CLK(clk),
    .D(_03545_),
    .Q(\datamem.data_ram[7][26] ));
 sky130_fd_sc_hd__dfxtp_1 _32124_ (.CLK(clk),
    .D(_03546_),
    .Q(\datamem.data_ram[7][27] ));
 sky130_fd_sc_hd__dfxtp_1 _32125_ (.CLK(clk),
    .D(_03547_),
    .Q(\datamem.data_ram[7][28] ));
 sky130_fd_sc_hd__dfxtp_1 _32126_ (.CLK(clk),
    .D(_03548_),
    .Q(\datamem.data_ram[7][29] ));
 sky130_fd_sc_hd__dfxtp_1 _32127_ (.CLK(clk),
    .D(_03549_),
    .Q(\datamem.data_ram[7][30] ));
 sky130_fd_sc_hd__dfxtp_1 _32128_ (.CLK(clk),
    .D(_03550_),
    .Q(\datamem.data_ram[7][31] ));
 sky130_fd_sc_hd__dfxtp_1 _32129_ (.CLK(clk),
    .D(_03551_),
    .Q(\datamem.data_ram[10][24] ));
 sky130_fd_sc_hd__dfxtp_1 _32130_ (.CLK(clk),
    .D(_03552_),
    .Q(\datamem.data_ram[10][25] ));
 sky130_fd_sc_hd__dfxtp_1 _32131_ (.CLK(clk),
    .D(_03553_),
    .Q(\datamem.data_ram[10][26] ));
 sky130_fd_sc_hd__dfxtp_1 _32132_ (.CLK(clk),
    .D(_03554_),
    .Q(\datamem.data_ram[10][27] ));
 sky130_fd_sc_hd__dfxtp_1 _32133_ (.CLK(clk),
    .D(_03555_),
    .Q(\datamem.data_ram[10][28] ));
 sky130_fd_sc_hd__dfxtp_1 _32134_ (.CLK(clk),
    .D(_03556_),
    .Q(\datamem.data_ram[10][29] ));
 sky130_fd_sc_hd__dfxtp_1 _32135_ (.CLK(clk),
    .D(_03557_),
    .Q(\datamem.data_ram[10][30] ));
 sky130_fd_sc_hd__dfxtp_1 _32136_ (.CLK(clk),
    .D(_03558_),
    .Q(\datamem.data_ram[10][31] ));
 sky130_fd_sc_hd__dfxtp_1 _32137_ (.CLK(clk),
    .D(_03559_),
    .Q(\datamem.data_ram[39][8] ));
 sky130_fd_sc_hd__dfxtp_1 _32138_ (.CLK(clk),
    .D(_03560_),
    .Q(\datamem.data_ram[39][9] ));
 sky130_fd_sc_hd__dfxtp_1 _32139_ (.CLK(clk),
    .D(_03561_),
    .Q(\datamem.data_ram[39][10] ));
 sky130_fd_sc_hd__dfxtp_1 _32140_ (.CLK(clk),
    .D(_03562_),
    .Q(\datamem.data_ram[39][11] ));
 sky130_fd_sc_hd__dfxtp_1 _32141_ (.CLK(clk),
    .D(_03563_),
    .Q(\datamem.data_ram[39][12] ));
 sky130_fd_sc_hd__dfxtp_1 _32142_ (.CLK(clk),
    .D(_03564_),
    .Q(\datamem.data_ram[39][13] ));
 sky130_fd_sc_hd__dfxtp_1 _32143_ (.CLK(clk),
    .D(_03565_),
    .Q(\datamem.data_ram[39][14] ));
 sky130_fd_sc_hd__dfxtp_1 _32144_ (.CLK(clk),
    .D(_03566_),
    .Q(\datamem.data_ram[39][15] ));
 sky130_fd_sc_hd__dfxtp_1 _32145_ (.CLK(clk),
    .D(_03567_),
    .Q(\datamem.data_ram[38][24] ));
 sky130_fd_sc_hd__dfxtp_1 _32146_ (.CLK(clk),
    .D(_03568_),
    .Q(\datamem.data_ram[38][25] ));
 sky130_fd_sc_hd__dfxtp_1 _32147_ (.CLK(clk),
    .D(_03569_),
    .Q(\datamem.data_ram[38][26] ));
 sky130_fd_sc_hd__dfxtp_1 _32148_ (.CLK(clk),
    .D(_03570_),
    .Q(\datamem.data_ram[38][27] ));
 sky130_fd_sc_hd__dfxtp_1 _32149_ (.CLK(clk),
    .D(_03571_),
    .Q(\datamem.data_ram[38][28] ));
 sky130_fd_sc_hd__dfxtp_1 _32150_ (.CLK(clk),
    .D(_03572_),
    .Q(\datamem.data_ram[38][29] ));
 sky130_fd_sc_hd__dfxtp_1 _32151_ (.CLK(clk),
    .D(_03573_),
    .Q(\datamem.data_ram[38][30] ));
 sky130_fd_sc_hd__dfxtp_1 _32152_ (.CLK(clk),
    .D(_03574_),
    .Q(\datamem.data_ram[38][31] ));
 sky130_fd_sc_hd__dfxtp_1 _32153_ (.CLK(clk),
    .D(_03575_),
    .Q(\datamem.data_ram[38][16] ));
 sky130_fd_sc_hd__dfxtp_1 _32154_ (.CLK(clk),
    .D(_03576_),
    .Q(\datamem.data_ram[38][17] ));
 sky130_fd_sc_hd__dfxtp_1 _32155_ (.CLK(clk),
    .D(_03577_),
    .Q(\datamem.data_ram[38][18] ));
 sky130_fd_sc_hd__dfxtp_1 _32156_ (.CLK(clk),
    .D(_03578_),
    .Q(\datamem.data_ram[38][19] ));
 sky130_fd_sc_hd__dfxtp_1 _32157_ (.CLK(clk),
    .D(_03579_),
    .Q(\datamem.data_ram[38][20] ));
 sky130_fd_sc_hd__dfxtp_1 _32158_ (.CLK(clk),
    .D(_03580_),
    .Q(\datamem.data_ram[38][21] ));
 sky130_fd_sc_hd__dfxtp_1 _32159_ (.CLK(clk),
    .D(_03581_),
    .Q(\datamem.data_ram[38][22] ));
 sky130_fd_sc_hd__dfxtp_1 _32160_ (.CLK(clk),
    .D(_03582_),
    .Q(\datamem.data_ram[38][23] ));
 sky130_fd_sc_hd__dfxtp_1 _32161_ (.CLK(clk),
    .D(_03583_),
    .Q(\datamem.data_ram[38][8] ));
 sky130_fd_sc_hd__dfxtp_1 _32162_ (.CLK(clk),
    .D(_03584_),
    .Q(\datamem.data_ram[38][9] ));
 sky130_fd_sc_hd__dfxtp_1 _32163_ (.CLK(clk),
    .D(_03585_),
    .Q(\datamem.data_ram[38][10] ));
 sky130_fd_sc_hd__dfxtp_1 _32164_ (.CLK(clk),
    .D(_03586_),
    .Q(\datamem.data_ram[38][11] ));
 sky130_fd_sc_hd__dfxtp_1 _32165_ (.CLK(clk),
    .D(_03587_),
    .Q(\datamem.data_ram[38][12] ));
 sky130_fd_sc_hd__dfxtp_1 _32166_ (.CLK(clk),
    .D(_03588_),
    .Q(\datamem.data_ram[38][13] ));
 sky130_fd_sc_hd__dfxtp_1 _32167_ (.CLK(clk),
    .D(_03589_),
    .Q(\datamem.data_ram[38][14] ));
 sky130_fd_sc_hd__dfxtp_1 _32168_ (.CLK(clk),
    .D(_03590_),
    .Q(\datamem.data_ram[38][15] ));
 sky130_fd_sc_hd__dfxtp_1 _32169_ (.CLK(clk),
    .D(_03591_),
    .Q(\datamem.data_ram[37][24] ));
 sky130_fd_sc_hd__dfxtp_1 _32170_ (.CLK(clk),
    .D(_03592_),
    .Q(\datamem.data_ram[37][25] ));
 sky130_fd_sc_hd__dfxtp_1 _32171_ (.CLK(clk),
    .D(_03593_),
    .Q(\datamem.data_ram[37][26] ));
 sky130_fd_sc_hd__dfxtp_1 _32172_ (.CLK(clk),
    .D(_03594_),
    .Q(\datamem.data_ram[37][27] ));
 sky130_fd_sc_hd__dfxtp_1 _32173_ (.CLK(clk),
    .D(_03595_),
    .Q(\datamem.data_ram[37][28] ));
 sky130_fd_sc_hd__dfxtp_1 _32174_ (.CLK(clk),
    .D(_03596_),
    .Q(\datamem.data_ram[37][29] ));
 sky130_fd_sc_hd__dfxtp_1 _32175_ (.CLK(clk),
    .D(_03597_),
    .Q(\datamem.data_ram[37][30] ));
 sky130_fd_sc_hd__dfxtp_1 _32176_ (.CLK(clk),
    .D(_03598_),
    .Q(\datamem.data_ram[37][31] ));
 sky130_fd_sc_hd__dfxtp_1 _32177_ (.CLK(clk),
    .D(_03599_),
    .Q(\datamem.data_ram[37][16] ));
 sky130_fd_sc_hd__dfxtp_1 _32178_ (.CLK(clk),
    .D(_03600_),
    .Q(\datamem.data_ram[37][17] ));
 sky130_fd_sc_hd__dfxtp_1 _32179_ (.CLK(clk),
    .D(_03601_),
    .Q(\datamem.data_ram[37][18] ));
 sky130_fd_sc_hd__dfxtp_1 _32180_ (.CLK(clk),
    .D(_03602_),
    .Q(\datamem.data_ram[37][19] ));
 sky130_fd_sc_hd__dfxtp_1 _32181_ (.CLK(clk),
    .D(_03603_),
    .Q(\datamem.data_ram[37][20] ));
 sky130_fd_sc_hd__dfxtp_1 _32182_ (.CLK(clk),
    .D(_03604_),
    .Q(\datamem.data_ram[37][21] ));
 sky130_fd_sc_hd__dfxtp_1 _32183_ (.CLK(clk),
    .D(_03605_),
    .Q(\datamem.data_ram[37][22] ));
 sky130_fd_sc_hd__dfxtp_1 _32184_ (.CLK(clk),
    .D(_03606_),
    .Q(\datamem.data_ram[37][23] ));
 sky130_fd_sc_hd__dfxtp_1 _32185_ (.CLK(clk),
    .D(_03607_),
    .Q(\datamem.data_ram[37][8] ));
 sky130_fd_sc_hd__dfxtp_1 _32186_ (.CLK(clk),
    .D(_03608_),
    .Q(\datamem.data_ram[37][9] ));
 sky130_fd_sc_hd__dfxtp_1 _32187_ (.CLK(clk),
    .D(_03609_),
    .Q(\datamem.data_ram[37][10] ));
 sky130_fd_sc_hd__dfxtp_1 _32188_ (.CLK(clk),
    .D(_03610_),
    .Q(\datamem.data_ram[37][11] ));
 sky130_fd_sc_hd__dfxtp_1 _32189_ (.CLK(clk),
    .D(_03611_),
    .Q(\datamem.data_ram[37][12] ));
 sky130_fd_sc_hd__dfxtp_1 _32190_ (.CLK(clk),
    .D(_03612_),
    .Q(\datamem.data_ram[37][13] ));
 sky130_fd_sc_hd__dfxtp_1 _32191_ (.CLK(clk),
    .D(_03613_),
    .Q(\datamem.data_ram[37][14] ));
 sky130_fd_sc_hd__dfxtp_1 _32192_ (.CLK(clk),
    .D(_03614_),
    .Q(\datamem.data_ram[37][15] ));
 sky130_fd_sc_hd__dfxtp_1 _32193_ (.CLK(clk),
    .D(_03615_),
    .Q(\datamem.data_ram[36][24] ));
 sky130_fd_sc_hd__dfxtp_1 _32194_ (.CLK(clk),
    .D(_03616_),
    .Q(\datamem.data_ram[36][25] ));
 sky130_fd_sc_hd__dfxtp_1 _32195_ (.CLK(clk),
    .D(_03617_),
    .Q(\datamem.data_ram[36][26] ));
 sky130_fd_sc_hd__dfxtp_1 _32196_ (.CLK(clk),
    .D(_03618_),
    .Q(\datamem.data_ram[36][27] ));
 sky130_fd_sc_hd__dfxtp_1 _32197_ (.CLK(clk),
    .D(_03619_),
    .Q(\datamem.data_ram[36][28] ));
 sky130_fd_sc_hd__dfxtp_1 _32198_ (.CLK(clk),
    .D(_03620_),
    .Q(\datamem.data_ram[36][29] ));
 sky130_fd_sc_hd__dfxtp_1 _32199_ (.CLK(clk),
    .D(_03621_),
    .Q(\datamem.data_ram[36][30] ));
 sky130_fd_sc_hd__dfxtp_1 _32200_ (.CLK(clk),
    .D(_03622_),
    .Q(\datamem.data_ram[36][31] ));
 sky130_fd_sc_hd__dfxtp_1 _32201_ (.CLK(clk),
    .D(_03623_),
    .Q(\datamem.data_ram[36][16] ));
 sky130_fd_sc_hd__dfxtp_1 _32202_ (.CLK(clk),
    .D(_03624_),
    .Q(\datamem.data_ram[36][17] ));
 sky130_fd_sc_hd__dfxtp_1 _32203_ (.CLK(clk),
    .D(_03625_),
    .Q(\datamem.data_ram[36][18] ));
 sky130_fd_sc_hd__dfxtp_1 _32204_ (.CLK(clk),
    .D(_03626_),
    .Q(\datamem.data_ram[36][19] ));
 sky130_fd_sc_hd__dfxtp_1 _32205_ (.CLK(clk),
    .D(_03627_),
    .Q(\datamem.data_ram[36][20] ));
 sky130_fd_sc_hd__dfxtp_1 _32206_ (.CLK(clk),
    .D(_03628_),
    .Q(\datamem.data_ram[36][21] ));
 sky130_fd_sc_hd__dfxtp_1 _32207_ (.CLK(clk),
    .D(_03629_),
    .Q(\datamem.data_ram[36][22] ));
 sky130_fd_sc_hd__dfxtp_1 _32208_ (.CLK(clk),
    .D(_03630_),
    .Q(\datamem.data_ram[36][23] ));
 sky130_fd_sc_hd__dfxtp_1 _32209_ (.CLK(clk),
    .D(_03631_),
    .Q(\datamem.data_ram[36][8] ));
 sky130_fd_sc_hd__dfxtp_1 _32210_ (.CLK(clk),
    .D(_03632_),
    .Q(\datamem.data_ram[36][9] ));
 sky130_fd_sc_hd__dfxtp_1 _32211_ (.CLK(clk),
    .D(_03633_),
    .Q(\datamem.data_ram[36][10] ));
 sky130_fd_sc_hd__dfxtp_1 _32212_ (.CLK(clk),
    .D(_03634_),
    .Q(\datamem.data_ram[36][11] ));
 sky130_fd_sc_hd__dfxtp_1 _32213_ (.CLK(clk),
    .D(_03635_),
    .Q(\datamem.data_ram[36][12] ));
 sky130_fd_sc_hd__dfxtp_1 _32214_ (.CLK(clk),
    .D(_03636_),
    .Q(\datamem.data_ram[36][13] ));
 sky130_fd_sc_hd__dfxtp_1 _32215_ (.CLK(clk),
    .D(_03637_),
    .Q(\datamem.data_ram[36][14] ));
 sky130_fd_sc_hd__dfxtp_1 _32216_ (.CLK(clk),
    .D(_03638_),
    .Q(\datamem.data_ram[36][15] ));
 sky130_fd_sc_hd__dfxtp_1 _32217_ (.CLK(clk),
    .D(_03639_),
    .Q(\datamem.data_ram[35][24] ));
 sky130_fd_sc_hd__dfxtp_1 _32218_ (.CLK(clk),
    .D(_03640_),
    .Q(\datamem.data_ram[35][25] ));
 sky130_fd_sc_hd__dfxtp_1 _32219_ (.CLK(clk),
    .D(_03641_),
    .Q(\datamem.data_ram[35][26] ));
 sky130_fd_sc_hd__dfxtp_1 _32220_ (.CLK(clk),
    .D(_03642_),
    .Q(\datamem.data_ram[35][27] ));
 sky130_fd_sc_hd__dfxtp_1 _32221_ (.CLK(clk),
    .D(_03643_),
    .Q(\datamem.data_ram[35][28] ));
 sky130_fd_sc_hd__dfxtp_1 _32222_ (.CLK(clk),
    .D(_03644_),
    .Q(\datamem.data_ram[35][29] ));
 sky130_fd_sc_hd__dfxtp_1 _32223_ (.CLK(clk),
    .D(_03645_),
    .Q(\datamem.data_ram[35][30] ));
 sky130_fd_sc_hd__dfxtp_1 _32224_ (.CLK(clk),
    .D(_03646_),
    .Q(\datamem.data_ram[35][31] ));
 sky130_fd_sc_hd__dfxtp_1 _32225_ (.CLK(clk),
    .D(_03647_),
    .Q(\datamem.data_ram[35][16] ));
 sky130_fd_sc_hd__dfxtp_1 _32226_ (.CLK(clk),
    .D(_03648_),
    .Q(\datamem.data_ram[35][17] ));
 sky130_fd_sc_hd__dfxtp_1 _32227_ (.CLK(clk),
    .D(_03649_),
    .Q(\datamem.data_ram[35][18] ));
 sky130_fd_sc_hd__dfxtp_1 _32228_ (.CLK(clk),
    .D(_03650_),
    .Q(\datamem.data_ram[35][19] ));
 sky130_fd_sc_hd__dfxtp_1 _32229_ (.CLK(clk),
    .D(_03651_),
    .Q(\datamem.data_ram[35][20] ));
 sky130_fd_sc_hd__dfxtp_1 _32230_ (.CLK(clk),
    .D(_03652_),
    .Q(\datamem.data_ram[35][21] ));
 sky130_fd_sc_hd__dfxtp_1 _32231_ (.CLK(clk),
    .D(_03653_),
    .Q(\datamem.data_ram[35][22] ));
 sky130_fd_sc_hd__dfxtp_1 _32232_ (.CLK(clk),
    .D(_03654_),
    .Q(\datamem.data_ram[35][23] ));
 sky130_fd_sc_hd__dfxtp_1 _32233_ (.CLK(clk),
    .D(_03655_),
    .Q(\datamem.data_ram[35][8] ));
 sky130_fd_sc_hd__dfxtp_1 _32234_ (.CLK(clk),
    .D(_03656_),
    .Q(\datamem.data_ram[35][9] ));
 sky130_fd_sc_hd__dfxtp_1 _32235_ (.CLK(clk),
    .D(_03657_),
    .Q(\datamem.data_ram[35][10] ));
 sky130_fd_sc_hd__dfxtp_1 _32236_ (.CLK(clk),
    .D(_03658_),
    .Q(\datamem.data_ram[35][11] ));
 sky130_fd_sc_hd__dfxtp_1 _32237_ (.CLK(clk),
    .D(_03659_),
    .Q(\datamem.data_ram[35][12] ));
 sky130_fd_sc_hd__dfxtp_1 _32238_ (.CLK(clk),
    .D(_03660_),
    .Q(\datamem.data_ram[35][13] ));
 sky130_fd_sc_hd__dfxtp_1 _32239_ (.CLK(clk),
    .D(_03661_),
    .Q(\datamem.data_ram[35][14] ));
 sky130_fd_sc_hd__dfxtp_1 _32240_ (.CLK(clk),
    .D(_03662_),
    .Q(\datamem.data_ram[35][15] ));
 sky130_fd_sc_hd__dfxtp_1 _32241_ (.CLK(clk),
    .D(_03663_),
    .Q(\datamem.data_ram[34][24] ));
 sky130_fd_sc_hd__dfxtp_1 _32242_ (.CLK(clk),
    .D(_03664_),
    .Q(\datamem.data_ram[34][25] ));
 sky130_fd_sc_hd__dfxtp_1 _32243_ (.CLK(clk),
    .D(_03665_),
    .Q(\datamem.data_ram[34][26] ));
 sky130_fd_sc_hd__dfxtp_1 _32244_ (.CLK(clk),
    .D(_03666_),
    .Q(\datamem.data_ram[34][27] ));
 sky130_fd_sc_hd__dfxtp_1 _32245_ (.CLK(clk),
    .D(_03667_),
    .Q(\datamem.data_ram[34][28] ));
 sky130_fd_sc_hd__dfxtp_1 _32246_ (.CLK(clk),
    .D(_03668_),
    .Q(\datamem.data_ram[34][29] ));
 sky130_fd_sc_hd__dfxtp_1 _32247_ (.CLK(clk),
    .D(_03669_),
    .Q(\datamem.data_ram[34][30] ));
 sky130_fd_sc_hd__dfxtp_1 _32248_ (.CLK(clk),
    .D(_03670_),
    .Q(\datamem.data_ram[34][31] ));
 sky130_fd_sc_hd__dfxtp_1 _32249_ (.CLK(clk),
    .D(_03671_),
    .Q(\datamem.data_ram[34][16] ));
 sky130_fd_sc_hd__dfxtp_1 _32250_ (.CLK(clk),
    .D(_03672_),
    .Q(\datamem.data_ram[34][17] ));
 sky130_fd_sc_hd__dfxtp_1 _32251_ (.CLK(clk),
    .D(_03673_),
    .Q(\datamem.data_ram[34][18] ));
 sky130_fd_sc_hd__dfxtp_1 _32252_ (.CLK(clk),
    .D(_03674_),
    .Q(\datamem.data_ram[34][19] ));
 sky130_fd_sc_hd__dfxtp_1 _32253_ (.CLK(clk),
    .D(_03675_),
    .Q(\datamem.data_ram[34][20] ));
 sky130_fd_sc_hd__dfxtp_1 _32254_ (.CLK(clk),
    .D(_03676_),
    .Q(\datamem.data_ram[34][21] ));
 sky130_fd_sc_hd__dfxtp_1 _32255_ (.CLK(clk),
    .D(_03677_),
    .Q(\datamem.data_ram[34][22] ));
 sky130_fd_sc_hd__dfxtp_1 _32256_ (.CLK(clk),
    .D(_03678_),
    .Q(\datamem.data_ram[34][23] ));
 sky130_fd_sc_hd__dfxtp_1 _32257_ (.CLK(clk),
    .D(_03679_),
    .Q(\datamem.data_ram[34][8] ));
 sky130_fd_sc_hd__dfxtp_1 _32258_ (.CLK(clk),
    .D(_03680_),
    .Q(\datamem.data_ram[34][9] ));
 sky130_fd_sc_hd__dfxtp_1 _32259_ (.CLK(clk),
    .D(_03681_),
    .Q(\datamem.data_ram[34][10] ));
 sky130_fd_sc_hd__dfxtp_1 _32260_ (.CLK(clk),
    .D(_03682_),
    .Q(\datamem.data_ram[34][11] ));
 sky130_fd_sc_hd__dfxtp_1 _32261_ (.CLK(clk),
    .D(_03683_),
    .Q(\datamem.data_ram[34][12] ));
 sky130_fd_sc_hd__dfxtp_1 _32262_ (.CLK(clk),
    .D(_03684_),
    .Q(\datamem.data_ram[34][13] ));
 sky130_fd_sc_hd__dfxtp_1 _32263_ (.CLK(clk),
    .D(_03685_),
    .Q(\datamem.data_ram[34][14] ));
 sky130_fd_sc_hd__dfxtp_1 _32264_ (.CLK(clk),
    .D(_03686_),
    .Q(\datamem.data_ram[34][15] ));
 sky130_fd_sc_hd__dfxtp_1 _32265_ (.CLK(clk),
    .D(_03687_),
    .Q(\datamem.data_ram[33][24] ));
 sky130_fd_sc_hd__dfxtp_1 _32266_ (.CLK(clk),
    .D(_03688_),
    .Q(\datamem.data_ram[33][25] ));
 sky130_fd_sc_hd__dfxtp_1 _32267_ (.CLK(clk),
    .D(_03689_),
    .Q(\datamem.data_ram[33][26] ));
 sky130_fd_sc_hd__dfxtp_1 _32268_ (.CLK(clk),
    .D(_03690_),
    .Q(\datamem.data_ram[33][27] ));
 sky130_fd_sc_hd__dfxtp_1 _32269_ (.CLK(clk),
    .D(_03691_),
    .Q(\datamem.data_ram[33][28] ));
 sky130_fd_sc_hd__dfxtp_1 _32270_ (.CLK(clk),
    .D(_03692_),
    .Q(\datamem.data_ram[33][29] ));
 sky130_fd_sc_hd__dfxtp_1 _32271_ (.CLK(clk),
    .D(_03693_),
    .Q(\datamem.data_ram[33][30] ));
 sky130_fd_sc_hd__dfxtp_1 _32272_ (.CLK(clk),
    .D(_03694_),
    .Q(\datamem.data_ram[33][31] ));
 sky130_fd_sc_hd__dfxtp_1 _32273_ (.CLK(clk),
    .D(_03695_),
    .Q(\datamem.data_ram[33][16] ));
 sky130_fd_sc_hd__dfxtp_1 _32274_ (.CLK(clk),
    .D(_03696_),
    .Q(\datamem.data_ram[33][17] ));
 sky130_fd_sc_hd__dfxtp_1 _32275_ (.CLK(clk),
    .D(_03697_),
    .Q(\datamem.data_ram[33][18] ));
 sky130_fd_sc_hd__dfxtp_1 _32276_ (.CLK(clk),
    .D(_03698_),
    .Q(\datamem.data_ram[33][19] ));
 sky130_fd_sc_hd__dfxtp_1 _32277_ (.CLK(clk),
    .D(_03699_),
    .Q(\datamem.data_ram[33][20] ));
 sky130_fd_sc_hd__dfxtp_1 _32278_ (.CLK(clk),
    .D(_03700_),
    .Q(\datamem.data_ram[33][21] ));
 sky130_fd_sc_hd__dfxtp_1 _32279_ (.CLK(clk),
    .D(_03701_),
    .Q(\datamem.data_ram[33][22] ));
 sky130_fd_sc_hd__dfxtp_1 _32280_ (.CLK(clk),
    .D(_03702_),
    .Q(\datamem.data_ram[33][23] ));
 sky130_fd_sc_hd__dfxtp_1 _32281_ (.CLK(clk),
    .D(_03703_),
    .Q(\datamem.data_ram[33][8] ));
 sky130_fd_sc_hd__dfxtp_1 _32282_ (.CLK(clk),
    .D(_03704_),
    .Q(\datamem.data_ram[33][9] ));
 sky130_fd_sc_hd__dfxtp_1 _32283_ (.CLK(clk),
    .D(_03705_),
    .Q(\datamem.data_ram[33][10] ));
 sky130_fd_sc_hd__dfxtp_1 _32284_ (.CLK(clk),
    .D(_03706_),
    .Q(\datamem.data_ram[33][11] ));
 sky130_fd_sc_hd__dfxtp_1 _32285_ (.CLK(clk),
    .D(_03707_),
    .Q(\datamem.data_ram[33][12] ));
 sky130_fd_sc_hd__dfxtp_1 _32286_ (.CLK(clk),
    .D(_03708_),
    .Q(\datamem.data_ram[33][13] ));
 sky130_fd_sc_hd__dfxtp_1 _32287_ (.CLK(clk),
    .D(_03709_),
    .Q(\datamem.data_ram[33][14] ));
 sky130_fd_sc_hd__dfxtp_1 _32288_ (.CLK(clk),
    .D(_03710_),
    .Q(\datamem.data_ram[33][15] ));
 sky130_fd_sc_hd__dfxtp_1 _32289_ (.CLK(clk),
    .D(_03711_),
    .Q(\datamem.data_ram[32][24] ));
 sky130_fd_sc_hd__dfxtp_1 _32290_ (.CLK(clk),
    .D(_03712_),
    .Q(\datamem.data_ram[32][25] ));
 sky130_fd_sc_hd__dfxtp_1 _32291_ (.CLK(clk),
    .D(_03713_),
    .Q(\datamem.data_ram[32][26] ));
 sky130_fd_sc_hd__dfxtp_1 _32292_ (.CLK(clk),
    .D(_03714_),
    .Q(\datamem.data_ram[32][27] ));
 sky130_fd_sc_hd__dfxtp_1 _32293_ (.CLK(clk),
    .D(_03715_),
    .Q(\datamem.data_ram[32][28] ));
 sky130_fd_sc_hd__dfxtp_1 _32294_ (.CLK(clk),
    .D(_03716_),
    .Q(\datamem.data_ram[32][29] ));
 sky130_fd_sc_hd__dfxtp_1 _32295_ (.CLK(clk),
    .D(_03717_),
    .Q(\datamem.data_ram[32][30] ));
 sky130_fd_sc_hd__dfxtp_1 _32296_ (.CLK(clk),
    .D(_03718_),
    .Q(\datamem.data_ram[32][31] ));
 sky130_fd_sc_hd__dfxtp_1 _32297_ (.CLK(clk),
    .D(_03719_),
    .Q(\datamem.data_ram[32][16] ));
 sky130_fd_sc_hd__dfxtp_1 _32298_ (.CLK(clk),
    .D(_03720_),
    .Q(\datamem.data_ram[32][17] ));
 sky130_fd_sc_hd__dfxtp_1 _32299_ (.CLK(clk),
    .D(_03721_),
    .Q(\datamem.data_ram[32][18] ));
 sky130_fd_sc_hd__dfxtp_1 _32300_ (.CLK(clk),
    .D(_03722_),
    .Q(\datamem.data_ram[32][19] ));
 sky130_fd_sc_hd__dfxtp_1 _32301_ (.CLK(clk),
    .D(_03723_),
    .Q(\datamem.data_ram[32][20] ));
 sky130_fd_sc_hd__dfxtp_1 _32302_ (.CLK(clk),
    .D(_03724_),
    .Q(\datamem.data_ram[32][21] ));
 sky130_fd_sc_hd__dfxtp_1 _32303_ (.CLK(clk),
    .D(_03725_),
    .Q(\datamem.data_ram[32][22] ));
 sky130_fd_sc_hd__dfxtp_1 _32304_ (.CLK(clk),
    .D(_03726_),
    .Q(\datamem.data_ram[32][23] ));
 sky130_fd_sc_hd__dfxtp_1 _32305_ (.CLK(clk),
    .D(_03727_),
    .Q(\datamem.data_ram[32][8] ));
 sky130_fd_sc_hd__dfxtp_1 _32306_ (.CLK(clk),
    .D(_03728_),
    .Q(\datamem.data_ram[32][9] ));
 sky130_fd_sc_hd__dfxtp_1 _32307_ (.CLK(clk),
    .D(_03729_),
    .Q(\datamem.data_ram[32][10] ));
 sky130_fd_sc_hd__dfxtp_1 _32308_ (.CLK(clk),
    .D(_03730_),
    .Q(\datamem.data_ram[32][11] ));
 sky130_fd_sc_hd__dfxtp_1 _32309_ (.CLK(clk),
    .D(_03731_),
    .Q(\datamem.data_ram[32][12] ));
 sky130_fd_sc_hd__dfxtp_1 _32310_ (.CLK(clk),
    .D(_03732_),
    .Q(\datamem.data_ram[32][13] ));
 sky130_fd_sc_hd__dfxtp_1 _32311_ (.CLK(clk),
    .D(_03733_),
    .Q(\datamem.data_ram[32][14] ));
 sky130_fd_sc_hd__dfxtp_1 _32312_ (.CLK(clk),
    .D(_03734_),
    .Q(\datamem.data_ram[32][15] ));
 sky130_fd_sc_hd__dfxtp_1 _32313_ (.CLK(clk),
    .D(_03735_),
    .Q(\datamem.data_ram[31][24] ));
 sky130_fd_sc_hd__dfxtp_1 _32314_ (.CLK(clk),
    .D(_03736_),
    .Q(\datamem.data_ram[31][25] ));
 sky130_fd_sc_hd__dfxtp_1 _32315_ (.CLK(clk),
    .D(_03737_),
    .Q(\datamem.data_ram[31][26] ));
 sky130_fd_sc_hd__dfxtp_1 _32316_ (.CLK(clk),
    .D(_03738_),
    .Q(\datamem.data_ram[31][27] ));
 sky130_fd_sc_hd__dfxtp_1 _32317_ (.CLK(clk),
    .D(_03739_),
    .Q(\datamem.data_ram[31][28] ));
 sky130_fd_sc_hd__dfxtp_1 _32318_ (.CLK(clk),
    .D(_03740_),
    .Q(\datamem.data_ram[31][29] ));
 sky130_fd_sc_hd__dfxtp_1 _32319_ (.CLK(clk),
    .D(_03741_),
    .Q(\datamem.data_ram[31][30] ));
 sky130_fd_sc_hd__dfxtp_1 _32320_ (.CLK(clk),
    .D(_03742_),
    .Q(\datamem.data_ram[31][31] ));
 sky130_fd_sc_hd__dfxtp_1 _32321_ (.CLK(clk),
    .D(_03743_),
    .Q(\datamem.data_ram[31][16] ));
 sky130_fd_sc_hd__dfxtp_1 _32322_ (.CLK(clk),
    .D(_03744_),
    .Q(\datamem.data_ram[31][17] ));
 sky130_fd_sc_hd__dfxtp_1 _32323_ (.CLK(clk),
    .D(_03745_),
    .Q(\datamem.data_ram[31][18] ));
 sky130_fd_sc_hd__dfxtp_1 _32324_ (.CLK(clk),
    .D(_03746_),
    .Q(\datamem.data_ram[31][19] ));
 sky130_fd_sc_hd__dfxtp_1 _32325_ (.CLK(clk),
    .D(_03747_),
    .Q(\datamem.data_ram[31][20] ));
 sky130_fd_sc_hd__dfxtp_1 _32326_ (.CLK(clk),
    .D(_03748_),
    .Q(\datamem.data_ram[31][21] ));
 sky130_fd_sc_hd__dfxtp_1 _32327_ (.CLK(clk),
    .D(_03749_),
    .Q(\datamem.data_ram[31][22] ));
 sky130_fd_sc_hd__dfxtp_1 _32328_ (.CLK(clk),
    .D(_03750_),
    .Q(\datamem.data_ram[31][23] ));
 sky130_fd_sc_hd__dfxtp_1 _32329_ (.CLK(clk),
    .D(_03751_),
    .Q(\datamem.data_ram[31][8] ));
 sky130_fd_sc_hd__dfxtp_1 _32330_ (.CLK(clk),
    .D(_03752_),
    .Q(\datamem.data_ram[31][9] ));
 sky130_fd_sc_hd__dfxtp_1 _32331_ (.CLK(clk),
    .D(_03753_),
    .Q(\datamem.data_ram[31][10] ));
 sky130_fd_sc_hd__dfxtp_1 _32332_ (.CLK(clk),
    .D(_03754_),
    .Q(\datamem.data_ram[31][11] ));
 sky130_fd_sc_hd__dfxtp_1 _32333_ (.CLK(clk),
    .D(_03755_),
    .Q(\datamem.data_ram[31][12] ));
 sky130_fd_sc_hd__dfxtp_1 _32334_ (.CLK(clk),
    .D(_03756_),
    .Q(\datamem.data_ram[31][13] ));
 sky130_fd_sc_hd__dfxtp_1 _32335_ (.CLK(clk),
    .D(_03757_),
    .Q(\datamem.data_ram[31][14] ));
 sky130_fd_sc_hd__dfxtp_1 _32336_ (.CLK(clk),
    .D(_03758_),
    .Q(\datamem.data_ram[31][15] ));
 sky130_fd_sc_hd__dfxtp_1 _32337_ (.CLK(clk),
    .D(_03759_),
    .Q(\datamem.data_ram[30][24] ));
 sky130_fd_sc_hd__dfxtp_1 _32338_ (.CLK(clk),
    .D(_03760_),
    .Q(\datamem.data_ram[30][25] ));
 sky130_fd_sc_hd__dfxtp_1 _32339_ (.CLK(clk),
    .D(_03761_),
    .Q(\datamem.data_ram[30][26] ));
 sky130_fd_sc_hd__dfxtp_1 _32340_ (.CLK(clk),
    .D(_03762_),
    .Q(\datamem.data_ram[30][27] ));
 sky130_fd_sc_hd__dfxtp_1 _32341_ (.CLK(clk),
    .D(_03763_),
    .Q(\datamem.data_ram[30][28] ));
 sky130_fd_sc_hd__dfxtp_1 _32342_ (.CLK(clk),
    .D(_03764_),
    .Q(\datamem.data_ram[30][29] ));
 sky130_fd_sc_hd__dfxtp_1 _32343_ (.CLK(clk),
    .D(_03765_),
    .Q(\datamem.data_ram[30][30] ));
 sky130_fd_sc_hd__dfxtp_1 _32344_ (.CLK(clk),
    .D(_03766_),
    .Q(\datamem.data_ram[30][31] ));
 sky130_fd_sc_hd__dfxtp_1 _32345_ (.CLK(clk),
    .D(_03767_),
    .Q(\datamem.data_ram[30][16] ));
 sky130_fd_sc_hd__dfxtp_1 _32346_ (.CLK(clk),
    .D(_03768_),
    .Q(\datamem.data_ram[30][17] ));
 sky130_fd_sc_hd__dfxtp_1 _32347_ (.CLK(clk),
    .D(_03769_),
    .Q(\datamem.data_ram[30][18] ));
 sky130_fd_sc_hd__dfxtp_1 _32348_ (.CLK(clk),
    .D(_03770_),
    .Q(\datamem.data_ram[30][19] ));
 sky130_fd_sc_hd__dfxtp_1 _32349_ (.CLK(clk),
    .D(_03771_),
    .Q(\datamem.data_ram[30][20] ));
 sky130_fd_sc_hd__dfxtp_1 _32350_ (.CLK(clk),
    .D(_03772_),
    .Q(\datamem.data_ram[30][21] ));
 sky130_fd_sc_hd__dfxtp_1 _32351_ (.CLK(clk),
    .D(_03773_),
    .Q(\datamem.data_ram[30][22] ));
 sky130_fd_sc_hd__dfxtp_1 _32352_ (.CLK(clk),
    .D(_03774_),
    .Q(\datamem.data_ram[30][23] ));
 sky130_fd_sc_hd__dfxtp_1 _32353_ (.CLK(clk),
    .D(_03775_),
    .Q(\datamem.data_ram[30][8] ));
 sky130_fd_sc_hd__dfxtp_1 _32354_ (.CLK(clk),
    .D(_03776_),
    .Q(\datamem.data_ram[30][9] ));
 sky130_fd_sc_hd__dfxtp_1 _32355_ (.CLK(clk),
    .D(_03777_),
    .Q(\datamem.data_ram[30][10] ));
 sky130_fd_sc_hd__dfxtp_1 _32356_ (.CLK(clk),
    .D(_03778_),
    .Q(\datamem.data_ram[30][11] ));
 sky130_fd_sc_hd__dfxtp_1 _32357_ (.CLK(clk),
    .D(_03779_),
    .Q(\datamem.data_ram[30][12] ));
 sky130_fd_sc_hd__dfxtp_1 _32358_ (.CLK(clk),
    .D(_03780_),
    .Q(\datamem.data_ram[30][13] ));
 sky130_fd_sc_hd__dfxtp_1 _32359_ (.CLK(clk),
    .D(_03781_),
    .Q(\datamem.data_ram[30][14] ));
 sky130_fd_sc_hd__dfxtp_1 _32360_ (.CLK(clk),
    .D(_03782_),
    .Q(\datamem.data_ram[30][15] ));
 sky130_fd_sc_hd__dfxtp_1 _32361_ (.CLK(clk),
    .D(_03783_),
    .Q(\datamem.data_ram[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _32362_ (.CLK(clk),
    .D(_03784_),
    .Q(\datamem.data_ram[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _32363_ (.CLK(clk),
    .D(_03785_),
    .Q(\datamem.data_ram[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _32364_ (.CLK(clk),
    .D(_03786_),
    .Q(\datamem.data_ram[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _32365_ (.CLK(clk),
    .D(_03787_),
    .Q(\datamem.data_ram[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _32366_ (.CLK(clk),
    .D(_03788_),
    .Q(\datamem.data_ram[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _32367_ (.CLK(clk),
    .D(_03789_),
    .Q(\datamem.data_ram[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _32368_ (.CLK(clk),
    .D(_03790_),
    .Q(\datamem.data_ram[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _32369_ (.CLK(clk),
    .D(_03791_),
    .Q(\datamem.data_ram[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _32370_ (.CLK(clk),
    .D(_03792_),
    .Q(\datamem.data_ram[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _32371_ (.CLK(clk),
    .D(_03793_),
    .Q(\datamem.data_ram[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _32372_ (.CLK(clk),
    .D(_03794_),
    .Q(\datamem.data_ram[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _32373_ (.CLK(clk),
    .D(_03795_),
    .Q(\datamem.data_ram[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _32374_ (.CLK(clk),
    .D(_03796_),
    .Q(\datamem.data_ram[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _32375_ (.CLK(clk),
    .D(_03797_),
    .Q(\datamem.data_ram[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _32376_ (.CLK(clk),
    .D(_03798_),
    .Q(\datamem.data_ram[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _32377_ (.CLK(clk),
    .D(_03799_),
    .Q(\datamem.data_ram[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _32378_ (.CLK(clk),
    .D(_03800_),
    .Q(\datamem.data_ram[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _32379_ (.CLK(clk),
    .D(_03801_),
    .Q(\datamem.data_ram[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _32380_ (.CLK(clk),
    .D(_03802_),
    .Q(\datamem.data_ram[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _32381_ (.CLK(clk),
    .D(_03803_),
    .Q(\datamem.data_ram[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _32382_ (.CLK(clk),
    .D(_03804_),
    .Q(\datamem.data_ram[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _32383_ (.CLK(clk),
    .D(_03805_),
    .Q(\datamem.data_ram[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _32384_ (.CLK(clk),
    .D(_03806_),
    .Q(\datamem.data_ram[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _32385_ (.CLK(clk),
    .D(_03807_),
    .Q(\datamem.data_ram[29][24] ));
 sky130_fd_sc_hd__dfxtp_1 _32386_ (.CLK(clk),
    .D(_03808_),
    .Q(\datamem.data_ram[29][25] ));
 sky130_fd_sc_hd__dfxtp_1 _32387_ (.CLK(clk),
    .D(_03809_),
    .Q(\datamem.data_ram[29][26] ));
 sky130_fd_sc_hd__dfxtp_1 _32388_ (.CLK(clk),
    .D(_03810_),
    .Q(\datamem.data_ram[29][27] ));
 sky130_fd_sc_hd__dfxtp_1 _32389_ (.CLK(clk),
    .D(_03811_),
    .Q(\datamem.data_ram[29][28] ));
 sky130_fd_sc_hd__dfxtp_1 _32390_ (.CLK(clk),
    .D(_03812_),
    .Q(\datamem.data_ram[29][29] ));
 sky130_fd_sc_hd__dfxtp_1 _32391_ (.CLK(clk),
    .D(_03813_),
    .Q(\datamem.data_ram[29][30] ));
 sky130_fd_sc_hd__dfxtp_1 _32392_ (.CLK(clk),
    .D(_03814_),
    .Q(\datamem.data_ram[29][31] ));
 sky130_fd_sc_hd__dfxtp_1 _32393_ (.CLK(clk),
    .D(_03815_),
    .Q(\datamem.data_ram[29][16] ));
 sky130_fd_sc_hd__dfxtp_1 _32394_ (.CLK(clk),
    .D(_03816_),
    .Q(\datamem.data_ram[29][17] ));
 sky130_fd_sc_hd__dfxtp_1 _32395_ (.CLK(clk),
    .D(_03817_),
    .Q(\datamem.data_ram[29][18] ));
 sky130_fd_sc_hd__dfxtp_1 _32396_ (.CLK(clk),
    .D(_03818_),
    .Q(\datamem.data_ram[29][19] ));
 sky130_fd_sc_hd__dfxtp_1 _32397_ (.CLK(clk),
    .D(_03819_),
    .Q(\datamem.data_ram[29][20] ));
 sky130_fd_sc_hd__dfxtp_1 _32398_ (.CLK(clk),
    .D(_03820_),
    .Q(\datamem.data_ram[29][21] ));
 sky130_fd_sc_hd__dfxtp_1 _32399_ (.CLK(clk),
    .D(_03821_),
    .Q(\datamem.data_ram[29][22] ));
 sky130_fd_sc_hd__dfxtp_1 _32400_ (.CLK(clk),
    .D(_03822_),
    .Q(\datamem.data_ram[29][23] ));
 sky130_fd_sc_hd__dfxtp_1 _32401_ (.CLK(clk),
    .D(_03823_),
    .Q(\datamem.data_ram[29][8] ));
 sky130_fd_sc_hd__dfxtp_1 _32402_ (.CLK(clk),
    .D(_03824_),
    .Q(\datamem.data_ram[29][9] ));
 sky130_fd_sc_hd__dfxtp_1 _32403_ (.CLK(clk),
    .D(_03825_),
    .Q(\datamem.data_ram[29][10] ));
 sky130_fd_sc_hd__dfxtp_1 _32404_ (.CLK(clk),
    .D(_03826_),
    .Q(\datamem.data_ram[29][11] ));
 sky130_fd_sc_hd__dfxtp_1 _32405_ (.CLK(clk),
    .D(_03827_),
    .Q(\datamem.data_ram[29][12] ));
 sky130_fd_sc_hd__dfxtp_1 _32406_ (.CLK(clk),
    .D(_03828_),
    .Q(\datamem.data_ram[29][13] ));
 sky130_fd_sc_hd__dfxtp_1 _32407_ (.CLK(clk),
    .D(_03829_),
    .Q(\datamem.data_ram[29][14] ));
 sky130_fd_sc_hd__dfxtp_1 _32408_ (.CLK(clk),
    .D(_03830_),
    .Q(\datamem.data_ram[29][15] ));
 sky130_fd_sc_hd__dfxtp_1 _32409_ (.CLK(clk),
    .D(_03831_),
    .Q(\datamem.data_ram[28][24] ));
 sky130_fd_sc_hd__dfxtp_1 _32410_ (.CLK(clk),
    .D(_03832_),
    .Q(\datamem.data_ram[28][25] ));
 sky130_fd_sc_hd__dfxtp_1 _32411_ (.CLK(clk),
    .D(_03833_),
    .Q(\datamem.data_ram[28][26] ));
 sky130_fd_sc_hd__dfxtp_1 _32412_ (.CLK(clk),
    .D(_03834_),
    .Q(\datamem.data_ram[28][27] ));
 sky130_fd_sc_hd__dfxtp_1 _32413_ (.CLK(clk),
    .D(_03835_),
    .Q(\datamem.data_ram[28][28] ));
 sky130_fd_sc_hd__dfxtp_1 _32414_ (.CLK(clk),
    .D(_03836_),
    .Q(\datamem.data_ram[28][29] ));
 sky130_fd_sc_hd__dfxtp_1 _32415_ (.CLK(clk),
    .D(_03837_),
    .Q(\datamem.data_ram[28][30] ));
 sky130_fd_sc_hd__dfxtp_1 _32416_ (.CLK(clk),
    .D(_03838_),
    .Q(\datamem.data_ram[28][31] ));
 sky130_fd_sc_hd__dfxtp_1 _32417_ (.CLK(clk),
    .D(_03839_),
    .Q(\datamem.data_ram[28][16] ));
 sky130_fd_sc_hd__dfxtp_1 _32418_ (.CLK(clk),
    .D(_03840_),
    .Q(\datamem.data_ram[28][17] ));
 sky130_fd_sc_hd__dfxtp_1 _32419_ (.CLK(clk),
    .D(_03841_),
    .Q(\datamem.data_ram[28][18] ));
 sky130_fd_sc_hd__dfxtp_1 _32420_ (.CLK(clk),
    .D(_03842_),
    .Q(\datamem.data_ram[28][19] ));
 sky130_fd_sc_hd__dfxtp_1 _32421_ (.CLK(clk),
    .D(_03843_),
    .Q(\datamem.data_ram[28][20] ));
 sky130_fd_sc_hd__dfxtp_1 _32422_ (.CLK(clk),
    .D(_03844_),
    .Q(\datamem.data_ram[28][21] ));
 sky130_fd_sc_hd__dfxtp_1 _32423_ (.CLK(clk),
    .D(_03845_),
    .Q(\datamem.data_ram[28][22] ));
 sky130_fd_sc_hd__dfxtp_1 _32424_ (.CLK(clk),
    .D(_03846_),
    .Q(\datamem.data_ram[28][23] ));
 sky130_fd_sc_hd__dfxtp_1 _32425_ (.CLK(clk),
    .D(_03847_),
    .Q(\datamem.data_ram[28][8] ));
 sky130_fd_sc_hd__dfxtp_1 _32426_ (.CLK(clk),
    .D(_03848_),
    .Q(\datamem.data_ram[28][9] ));
 sky130_fd_sc_hd__dfxtp_1 _32427_ (.CLK(clk),
    .D(_03849_),
    .Q(\datamem.data_ram[28][10] ));
 sky130_fd_sc_hd__dfxtp_1 _32428_ (.CLK(clk),
    .D(_03850_),
    .Q(\datamem.data_ram[28][11] ));
 sky130_fd_sc_hd__dfxtp_1 _32429_ (.CLK(clk),
    .D(_03851_),
    .Q(\datamem.data_ram[28][12] ));
 sky130_fd_sc_hd__dfxtp_1 _32430_ (.CLK(clk),
    .D(_03852_),
    .Q(\datamem.data_ram[28][13] ));
 sky130_fd_sc_hd__dfxtp_1 _32431_ (.CLK(clk),
    .D(_03853_),
    .Q(\datamem.data_ram[28][14] ));
 sky130_fd_sc_hd__dfxtp_1 _32432_ (.CLK(clk),
    .D(_03854_),
    .Q(\datamem.data_ram[28][15] ));
 sky130_fd_sc_hd__dfxtp_1 _32433_ (.CLK(clk),
    .D(_03855_),
    .Q(\datamem.data_ram[27][24] ));
 sky130_fd_sc_hd__dfxtp_1 _32434_ (.CLK(clk),
    .D(_03856_),
    .Q(\datamem.data_ram[27][25] ));
 sky130_fd_sc_hd__dfxtp_1 _32435_ (.CLK(clk),
    .D(_03857_),
    .Q(\datamem.data_ram[27][26] ));
 sky130_fd_sc_hd__dfxtp_1 _32436_ (.CLK(clk),
    .D(_03858_),
    .Q(\datamem.data_ram[27][27] ));
 sky130_fd_sc_hd__dfxtp_1 _32437_ (.CLK(clk),
    .D(_03859_),
    .Q(\datamem.data_ram[27][28] ));
 sky130_fd_sc_hd__dfxtp_1 _32438_ (.CLK(clk),
    .D(_03860_),
    .Q(\datamem.data_ram[27][29] ));
 sky130_fd_sc_hd__dfxtp_1 _32439_ (.CLK(clk),
    .D(_03861_),
    .Q(\datamem.data_ram[27][30] ));
 sky130_fd_sc_hd__dfxtp_1 _32440_ (.CLK(clk),
    .D(_03862_),
    .Q(\datamem.data_ram[27][31] ));
 sky130_fd_sc_hd__dfxtp_1 _32441_ (.CLK(clk),
    .D(_03863_),
    .Q(\datamem.data_ram[27][16] ));
 sky130_fd_sc_hd__dfxtp_1 _32442_ (.CLK(clk),
    .D(_03864_),
    .Q(\datamem.data_ram[27][17] ));
 sky130_fd_sc_hd__dfxtp_1 _32443_ (.CLK(clk),
    .D(_03865_),
    .Q(\datamem.data_ram[27][18] ));
 sky130_fd_sc_hd__dfxtp_1 _32444_ (.CLK(clk),
    .D(_03866_),
    .Q(\datamem.data_ram[27][19] ));
 sky130_fd_sc_hd__dfxtp_1 _32445_ (.CLK(clk),
    .D(_03867_),
    .Q(\datamem.data_ram[27][20] ));
 sky130_fd_sc_hd__dfxtp_1 _32446_ (.CLK(clk),
    .D(_03868_),
    .Q(\datamem.data_ram[27][21] ));
 sky130_fd_sc_hd__dfxtp_1 _32447_ (.CLK(clk),
    .D(_03869_),
    .Q(\datamem.data_ram[27][22] ));
 sky130_fd_sc_hd__dfxtp_1 _32448_ (.CLK(clk),
    .D(_03870_),
    .Q(\datamem.data_ram[27][23] ));
 sky130_fd_sc_hd__dfxtp_1 _32449_ (.CLK(clk),
    .D(_03871_),
    .Q(\datamem.data_ram[27][8] ));
 sky130_fd_sc_hd__dfxtp_1 _32450_ (.CLK(clk),
    .D(_03872_),
    .Q(\datamem.data_ram[27][9] ));
 sky130_fd_sc_hd__dfxtp_1 _32451_ (.CLK(clk),
    .D(_03873_),
    .Q(\datamem.data_ram[27][10] ));
 sky130_fd_sc_hd__dfxtp_1 _32452_ (.CLK(clk),
    .D(_03874_),
    .Q(\datamem.data_ram[27][11] ));
 sky130_fd_sc_hd__dfxtp_1 _32453_ (.CLK(clk),
    .D(_03875_),
    .Q(\datamem.data_ram[27][12] ));
 sky130_fd_sc_hd__dfxtp_1 _32454_ (.CLK(clk),
    .D(_03876_),
    .Q(\datamem.data_ram[27][13] ));
 sky130_fd_sc_hd__dfxtp_1 _32455_ (.CLK(clk),
    .D(_03877_),
    .Q(\datamem.data_ram[27][14] ));
 sky130_fd_sc_hd__dfxtp_1 _32456_ (.CLK(clk),
    .D(_03878_),
    .Q(\datamem.data_ram[27][15] ));
 sky130_fd_sc_hd__dfxtp_1 _32457_ (.CLK(clk),
    .D(_03879_),
    .Q(\datamem.data_ram[26][24] ));
 sky130_fd_sc_hd__dfxtp_1 _32458_ (.CLK(clk),
    .D(_03880_),
    .Q(\datamem.data_ram[26][25] ));
 sky130_fd_sc_hd__dfxtp_1 _32459_ (.CLK(clk),
    .D(_03881_),
    .Q(\datamem.data_ram[26][26] ));
 sky130_fd_sc_hd__dfxtp_1 _32460_ (.CLK(clk),
    .D(_03882_),
    .Q(\datamem.data_ram[26][27] ));
 sky130_fd_sc_hd__dfxtp_1 _32461_ (.CLK(clk),
    .D(_03883_),
    .Q(\datamem.data_ram[26][28] ));
 sky130_fd_sc_hd__dfxtp_1 _32462_ (.CLK(clk),
    .D(_03884_),
    .Q(\datamem.data_ram[26][29] ));
 sky130_fd_sc_hd__dfxtp_1 _32463_ (.CLK(clk),
    .D(_03885_),
    .Q(\datamem.data_ram[26][30] ));
 sky130_fd_sc_hd__dfxtp_1 _32464_ (.CLK(clk),
    .D(_03886_),
    .Q(\datamem.data_ram[26][31] ));
 sky130_fd_sc_hd__dfxtp_1 _32465_ (.CLK(clk),
    .D(_03887_),
    .Q(\datamem.data_ram[26][16] ));
 sky130_fd_sc_hd__dfxtp_1 _32466_ (.CLK(clk),
    .D(_03888_),
    .Q(\datamem.data_ram[26][17] ));
 sky130_fd_sc_hd__dfxtp_1 _32467_ (.CLK(clk),
    .D(_03889_),
    .Q(\datamem.data_ram[26][18] ));
 sky130_fd_sc_hd__dfxtp_1 _32468_ (.CLK(clk),
    .D(_03890_),
    .Q(\datamem.data_ram[26][19] ));
 sky130_fd_sc_hd__dfxtp_1 _32469_ (.CLK(clk),
    .D(_03891_),
    .Q(\datamem.data_ram[26][20] ));
 sky130_fd_sc_hd__dfxtp_1 _32470_ (.CLK(clk),
    .D(_03892_),
    .Q(\datamem.data_ram[26][21] ));
 sky130_fd_sc_hd__dfxtp_1 _32471_ (.CLK(clk),
    .D(_03893_),
    .Q(\datamem.data_ram[26][22] ));
 sky130_fd_sc_hd__dfxtp_1 _32472_ (.CLK(clk),
    .D(_03894_),
    .Q(\datamem.data_ram[26][23] ));
 sky130_fd_sc_hd__dfxtp_1 _32473_ (.CLK(clk),
    .D(_03895_),
    .Q(\datamem.data_ram[26][8] ));
 sky130_fd_sc_hd__dfxtp_1 _32474_ (.CLK(clk),
    .D(_03896_),
    .Q(\datamem.data_ram[26][9] ));
 sky130_fd_sc_hd__dfxtp_1 _32475_ (.CLK(clk),
    .D(_03897_),
    .Q(\datamem.data_ram[26][10] ));
 sky130_fd_sc_hd__dfxtp_1 _32476_ (.CLK(clk),
    .D(_03898_),
    .Q(\datamem.data_ram[26][11] ));
 sky130_fd_sc_hd__dfxtp_1 _32477_ (.CLK(clk),
    .D(_03899_),
    .Q(\datamem.data_ram[26][12] ));
 sky130_fd_sc_hd__dfxtp_1 _32478_ (.CLK(clk),
    .D(_03900_),
    .Q(\datamem.data_ram[26][13] ));
 sky130_fd_sc_hd__dfxtp_1 _32479_ (.CLK(clk),
    .D(_03901_),
    .Q(\datamem.data_ram[26][14] ));
 sky130_fd_sc_hd__dfxtp_1 _32480_ (.CLK(clk),
    .D(_03902_),
    .Q(\datamem.data_ram[26][15] ));
 sky130_fd_sc_hd__dfxtp_1 _32481_ (.CLK(clk),
    .D(_03903_),
    .Q(\datamem.data_ram[25][24] ));
 sky130_fd_sc_hd__dfxtp_1 _32482_ (.CLK(clk),
    .D(_03904_),
    .Q(\datamem.data_ram[25][25] ));
 sky130_fd_sc_hd__dfxtp_1 _32483_ (.CLK(clk),
    .D(_03905_),
    .Q(\datamem.data_ram[25][26] ));
 sky130_fd_sc_hd__dfxtp_1 _32484_ (.CLK(clk),
    .D(_03906_),
    .Q(\datamem.data_ram[25][27] ));
 sky130_fd_sc_hd__dfxtp_1 _32485_ (.CLK(clk),
    .D(_03907_),
    .Q(\datamem.data_ram[25][28] ));
 sky130_fd_sc_hd__dfxtp_1 _32486_ (.CLK(clk),
    .D(_03908_),
    .Q(\datamem.data_ram[25][29] ));
 sky130_fd_sc_hd__dfxtp_1 _32487_ (.CLK(clk),
    .D(_03909_),
    .Q(\datamem.data_ram[25][30] ));
 sky130_fd_sc_hd__dfxtp_1 _32488_ (.CLK(clk),
    .D(_03910_),
    .Q(\datamem.data_ram[25][31] ));
 sky130_fd_sc_hd__dfxtp_1 _32489_ (.CLK(clk),
    .D(_03911_),
    .Q(\datamem.data_ram[25][16] ));
 sky130_fd_sc_hd__dfxtp_1 _32490_ (.CLK(clk),
    .D(_03912_),
    .Q(\datamem.data_ram[25][17] ));
 sky130_fd_sc_hd__dfxtp_1 _32491_ (.CLK(clk),
    .D(_03913_),
    .Q(\datamem.data_ram[25][18] ));
 sky130_fd_sc_hd__dfxtp_1 _32492_ (.CLK(clk),
    .D(_03914_),
    .Q(\datamem.data_ram[25][19] ));
 sky130_fd_sc_hd__dfxtp_1 _32493_ (.CLK(clk),
    .D(_03915_),
    .Q(\datamem.data_ram[25][20] ));
 sky130_fd_sc_hd__dfxtp_1 _32494_ (.CLK(clk),
    .D(_03916_),
    .Q(\datamem.data_ram[25][21] ));
 sky130_fd_sc_hd__dfxtp_1 _32495_ (.CLK(clk),
    .D(_03917_),
    .Q(\datamem.data_ram[25][22] ));
 sky130_fd_sc_hd__dfxtp_1 _32496_ (.CLK(clk),
    .D(_03918_),
    .Q(\datamem.data_ram[25][23] ));
 sky130_fd_sc_hd__dfxtp_1 _32497_ (.CLK(clk),
    .D(_03919_),
    .Q(\datamem.data_ram[25][8] ));
 sky130_fd_sc_hd__dfxtp_1 _32498_ (.CLK(clk),
    .D(_03920_),
    .Q(\datamem.data_ram[25][9] ));
 sky130_fd_sc_hd__dfxtp_1 _32499_ (.CLK(clk),
    .D(_03921_),
    .Q(\datamem.data_ram[25][10] ));
 sky130_fd_sc_hd__dfxtp_1 _32500_ (.CLK(clk),
    .D(_03922_),
    .Q(\datamem.data_ram[25][11] ));
 sky130_fd_sc_hd__dfxtp_1 _32501_ (.CLK(clk),
    .D(_03923_),
    .Q(\datamem.data_ram[25][12] ));
 sky130_fd_sc_hd__dfxtp_1 _32502_ (.CLK(clk),
    .D(_03924_),
    .Q(\datamem.data_ram[25][13] ));
 sky130_fd_sc_hd__dfxtp_1 _32503_ (.CLK(clk),
    .D(_03925_),
    .Q(\datamem.data_ram[25][14] ));
 sky130_fd_sc_hd__dfxtp_1 _32504_ (.CLK(clk),
    .D(_03926_),
    .Q(\datamem.data_ram[25][15] ));
 sky130_fd_sc_hd__dfxtp_1 _32505_ (.CLK(clk),
    .D(_03927_),
    .Q(\datamem.data_ram[24][24] ));
 sky130_fd_sc_hd__dfxtp_1 _32506_ (.CLK(clk),
    .D(_03928_),
    .Q(\datamem.data_ram[24][25] ));
 sky130_fd_sc_hd__dfxtp_1 _32507_ (.CLK(clk),
    .D(_03929_),
    .Q(\datamem.data_ram[24][26] ));
 sky130_fd_sc_hd__dfxtp_1 _32508_ (.CLK(clk),
    .D(_03930_),
    .Q(\datamem.data_ram[24][27] ));
 sky130_fd_sc_hd__dfxtp_1 _32509_ (.CLK(clk),
    .D(_03931_),
    .Q(\datamem.data_ram[24][28] ));
 sky130_fd_sc_hd__dfxtp_1 _32510_ (.CLK(clk),
    .D(_03932_),
    .Q(\datamem.data_ram[24][29] ));
 sky130_fd_sc_hd__dfxtp_1 _32511_ (.CLK(clk),
    .D(_03933_),
    .Q(\datamem.data_ram[24][30] ));
 sky130_fd_sc_hd__dfxtp_1 _32512_ (.CLK(clk),
    .D(_03934_),
    .Q(\datamem.data_ram[24][31] ));
 sky130_fd_sc_hd__dfxtp_1 _32513_ (.CLK(clk),
    .D(_03935_),
    .Q(\datamem.data_ram[24][16] ));
 sky130_fd_sc_hd__dfxtp_1 _32514_ (.CLK(clk),
    .D(_03936_),
    .Q(\datamem.data_ram[24][17] ));
 sky130_fd_sc_hd__dfxtp_1 _32515_ (.CLK(clk),
    .D(_03937_),
    .Q(\datamem.data_ram[24][18] ));
 sky130_fd_sc_hd__dfxtp_1 _32516_ (.CLK(clk),
    .D(_03938_),
    .Q(\datamem.data_ram[24][19] ));
 sky130_fd_sc_hd__dfxtp_1 _32517_ (.CLK(clk),
    .D(_03939_),
    .Q(\datamem.data_ram[24][20] ));
 sky130_fd_sc_hd__dfxtp_1 _32518_ (.CLK(clk),
    .D(_03940_),
    .Q(\datamem.data_ram[24][21] ));
 sky130_fd_sc_hd__dfxtp_1 _32519_ (.CLK(clk),
    .D(_03941_),
    .Q(\datamem.data_ram[24][22] ));
 sky130_fd_sc_hd__dfxtp_1 _32520_ (.CLK(clk),
    .D(_03942_),
    .Q(\datamem.data_ram[24][23] ));
 sky130_fd_sc_hd__dfxtp_1 _32521_ (.CLK(clk),
    .D(_03943_),
    .Q(\datamem.data_ram[24][8] ));
 sky130_fd_sc_hd__dfxtp_1 _32522_ (.CLK(clk),
    .D(_03944_),
    .Q(\datamem.data_ram[24][9] ));
 sky130_fd_sc_hd__dfxtp_1 _32523_ (.CLK(clk),
    .D(_03945_),
    .Q(\datamem.data_ram[24][10] ));
 sky130_fd_sc_hd__dfxtp_1 _32524_ (.CLK(clk),
    .D(_03946_),
    .Q(\datamem.data_ram[24][11] ));
 sky130_fd_sc_hd__dfxtp_1 _32525_ (.CLK(clk),
    .D(_03947_),
    .Q(\datamem.data_ram[24][12] ));
 sky130_fd_sc_hd__dfxtp_1 _32526_ (.CLK(clk),
    .D(_03948_),
    .Q(\datamem.data_ram[24][13] ));
 sky130_fd_sc_hd__dfxtp_1 _32527_ (.CLK(clk),
    .D(_03949_),
    .Q(\datamem.data_ram[24][14] ));
 sky130_fd_sc_hd__dfxtp_1 _32528_ (.CLK(clk),
    .D(_03950_),
    .Q(\datamem.data_ram[24][15] ));
 sky130_fd_sc_hd__dfxtp_1 _32529_ (.CLK(clk),
    .D(_03951_),
    .Q(\datamem.data_ram[23][24] ));
 sky130_fd_sc_hd__dfxtp_1 _32530_ (.CLK(clk),
    .D(_03952_),
    .Q(\datamem.data_ram[23][25] ));
 sky130_fd_sc_hd__dfxtp_1 _32531_ (.CLK(clk),
    .D(_03953_),
    .Q(\datamem.data_ram[23][26] ));
 sky130_fd_sc_hd__dfxtp_1 _32532_ (.CLK(clk),
    .D(_03954_),
    .Q(\datamem.data_ram[23][27] ));
 sky130_fd_sc_hd__dfxtp_1 _32533_ (.CLK(clk),
    .D(_03955_),
    .Q(\datamem.data_ram[23][28] ));
 sky130_fd_sc_hd__dfxtp_1 _32534_ (.CLK(clk),
    .D(_03956_),
    .Q(\datamem.data_ram[23][29] ));
 sky130_fd_sc_hd__dfxtp_1 _32535_ (.CLK(clk),
    .D(_03957_),
    .Q(\datamem.data_ram[23][30] ));
 sky130_fd_sc_hd__dfxtp_1 _32536_ (.CLK(clk),
    .D(_03958_),
    .Q(\datamem.data_ram[23][31] ));
 sky130_fd_sc_hd__dfxtp_1 _32537_ (.CLK(clk),
    .D(_03959_),
    .Q(\datamem.data_ram[23][16] ));
 sky130_fd_sc_hd__dfxtp_1 _32538_ (.CLK(clk),
    .D(_03960_),
    .Q(\datamem.data_ram[23][17] ));
 sky130_fd_sc_hd__dfxtp_1 _32539_ (.CLK(clk),
    .D(_03961_),
    .Q(\datamem.data_ram[23][18] ));
 sky130_fd_sc_hd__dfxtp_1 _32540_ (.CLK(clk),
    .D(_03962_),
    .Q(\datamem.data_ram[23][19] ));
 sky130_fd_sc_hd__dfxtp_1 _32541_ (.CLK(clk),
    .D(_03963_),
    .Q(\datamem.data_ram[23][20] ));
 sky130_fd_sc_hd__dfxtp_1 _32542_ (.CLK(clk),
    .D(_03964_),
    .Q(\datamem.data_ram[23][21] ));
 sky130_fd_sc_hd__dfxtp_1 _32543_ (.CLK(clk),
    .D(_03965_),
    .Q(\datamem.data_ram[23][22] ));
 sky130_fd_sc_hd__dfxtp_1 _32544_ (.CLK(clk),
    .D(_03966_),
    .Q(\datamem.data_ram[23][23] ));
 sky130_fd_sc_hd__dfxtp_1 _32545_ (.CLK(clk),
    .D(_03967_),
    .Q(\datamem.data_ram[23][8] ));
 sky130_fd_sc_hd__dfxtp_1 _32546_ (.CLK(clk),
    .D(_03968_),
    .Q(\datamem.data_ram[23][9] ));
 sky130_fd_sc_hd__dfxtp_1 _32547_ (.CLK(clk),
    .D(_03969_),
    .Q(\datamem.data_ram[23][10] ));
 sky130_fd_sc_hd__dfxtp_1 _32548_ (.CLK(clk),
    .D(_03970_),
    .Q(\datamem.data_ram[23][11] ));
 sky130_fd_sc_hd__dfxtp_1 _32549_ (.CLK(clk),
    .D(_03971_),
    .Q(\datamem.data_ram[23][12] ));
 sky130_fd_sc_hd__dfxtp_1 _32550_ (.CLK(clk),
    .D(_03972_),
    .Q(\datamem.data_ram[23][13] ));
 sky130_fd_sc_hd__dfxtp_1 _32551_ (.CLK(clk),
    .D(_03973_),
    .Q(\datamem.data_ram[23][14] ));
 sky130_fd_sc_hd__dfxtp_1 _32552_ (.CLK(clk),
    .D(_03974_),
    .Q(\datamem.data_ram[23][15] ));
 sky130_fd_sc_hd__dfxtp_1 _32553_ (.CLK(clk),
    .D(_03975_),
    .Q(\datamem.data_ram[22][24] ));
 sky130_fd_sc_hd__dfxtp_1 _32554_ (.CLK(clk),
    .D(_03976_),
    .Q(\datamem.data_ram[22][25] ));
 sky130_fd_sc_hd__dfxtp_1 _32555_ (.CLK(clk),
    .D(_03977_),
    .Q(\datamem.data_ram[22][26] ));
 sky130_fd_sc_hd__dfxtp_1 _32556_ (.CLK(clk),
    .D(_03978_),
    .Q(\datamem.data_ram[22][27] ));
 sky130_fd_sc_hd__dfxtp_1 _32557_ (.CLK(clk),
    .D(_03979_),
    .Q(\datamem.data_ram[22][28] ));
 sky130_fd_sc_hd__dfxtp_1 _32558_ (.CLK(clk),
    .D(_03980_),
    .Q(\datamem.data_ram[22][29] ));
 sky130_fd_sc_hd__dfxtp_1 _32559_ (.CLK(clk),
    .D(_03981_),
    .Q(\datamem.data_ram[22][30] ));
 sky130_fd_sc_hd__dfxtp_1 _32560_ (.CLK(clk),
    .D(_03982_),
    .Q(\datamem.data_ram[22][31] ));
 sky130_fd_sc_hd__dfxtp_1 _32561_ (.CLK(clk),
    .D(_03983_),
    .Q(\datamem.data_ram[22][16] ));
 sky130_fd_sc_hd__dfxtp_1 _32562_ (.CLK(clk),
    .D(_03984_),
    .Q(\datamem.data_ram[22][17] ));
 sky130_fd_sc_hd__dfxtp_1 _32563_ (.CLK(clk),
    .D(_03985_),
    .Q(\datamem.data_ram[22][18] ));
 sky130_fd_sc_hd__dfxtp_1 _32564_ (.CLK(clk),
    .D(_03986_),
    .Q(\datamem.data_ram[22][19] ));
 sky130_fd_sc_hd__dfxtp_1 _32565_ (.CLK(clk),
    .D(_03987_),
    .Q(\datamem.data_ram[22][20] ));
 sky130_fd_sc_hd__dfxtp_1 _32566_ (.CLK(clk),
    .D(_03988_),
    .Q(\datamem.data_ram[22][21] ));
 sky130_fd_sc_hd__dfxtp_1 _32567_ (.CLK(clk),
    .D(_03989_),
    .Q(\datamem.data_ram[22][22] ));
 sky130_fd_sc_hd__dfxtp_1 _32568_ (.CLK(clk),
    .D(_03990_),
    .Q(\datamem.data_ram[22][23] ));
 sky130_fd_sc_hd__dfxtp_1 _32569_ (.CLK(clk),
    .D(_03991_),
    .Q(\datamem.data_ram[22][8] ));
 sky130_fd_sc_hd__dfxtp_1 _32570_ (.CLK(clk),
    .D(_03992_),
    .Q(\datamem.data_ram[22][9] ));
 sky130_fd_sc_hd__dfxtp_1 _32571_ (.CLK(clk),
    .D(_03993_),
    .Q(\datamem.data_ram[22][10] ));
 sky130_fd_sc_hd__dfxtp_1 _32572_ (.CLK(clk),
    .D(_03994_),
    .Q(\datamem.data_ram[22][11] ));
 sky130_fd_sc_hd__dfxtp_1 _32573_ (.CLK(clk),
    .D(_03995_),
    .Q(\datamem.data_ram[22][12] ));
 sky130_fd_sc_hd__dfxtp_1 _32574_ (.CLK(clk),
    .D(_03996_),
    .Q(\datamem.data_ram[22][13] ));
 sky130_fd_sc_hd__dfxtp_1 _32575_ (.CLK(clk),
    .D(_03997_),
    .Q(\datamem.data_ram[22][14] ));
 sky130_fd_sc_hd__dfxtp_1 _32576_ (.CLK(clk),
    .D(_03998_),
    .Q(\datamem.data_ram[22][15] ));
 sky130_fd_sc_hd__dfxtp_1 _32577_ (.CLK(clk),
    .D(_03999_),
    .Q(\datamem.data_ram[21][24] ));
 sky130_fd_sc_hd__dfxtp_1 _32578_ (.CLK(clk),
    .D(_04000_),
    .Q(\datamem.data_ram[21][25] ));
 sky130_fd_sc_hd__dfxtp_1 _32579_ (.CLK(clk),
    .D(_04001_),
    .Q(\datamem.data_ram[21][26] ));
 sky130_fd_sc_hd__dfxtp_1 _32580_ (.CLK(clk),
    .D(_04002_),
    .Q(\datamem.data_ram[21][27] ));
 sky130_fd_sc_hd__dfxtp_1 _32581_ (.CLK(clk),
    .D(_04003_),
    .Q(\datamem.data_ram[21][28] ));
 sky130_fd_sc_hd__dfxtp_1 _32582_ (.CLK(clk),
    .D(_04004_),
    .Q(\datamem.data_ram[21][29] ));
 sky130_fd_sc_hd__dfxtp_1 _32583_ (.CLK(clk),
    .D(_04005_),
    .Q(\datamem.data_ram[21][30] ));
 sky130_fd_sc_hd__dfxtp_1 _32584_ (.CLK(clk),
    .D(_04006_),
    .Q(\datamem.data_ram[21][31] ));
 sky130_fd_sc_hd__dfxtp_1 _32585_ (.CLK(clk),
    .D(_04007_),
    .Q(\datamem.data_ram[21][16] ));
 sky130_fd_sc_hd__dfxtp_1 _32586_ (.CLK(clk),
    .D(_04008_),
    .Q(\datamem.data_ram[21][17] ));
 sky130_fd_sc_hd__dfxtp_1 _32587_ (.CLK(clk),
    .D(_04009_),
    .Q(\datamem.data_ram[21][18] ));
 sky130_fd_sc_hd__dfxtp_1 _32588_ (.CLK(clk),
    .D(_04010_),
    .Q(\datamem.data_ram[21][19] ));
 sky130_fd_sc_hd__dfxtp_1 _32589_ (.CLK(clk),
    .D(_04011_),
    .Q(\datamem.data_ram[21][20] ));
 sky130_fd_sc_hd__dfxtp_1 _32590_ (.CLK(clk),
    .D(_04012_),
    .Q(\datamem.data_ram[21][21] ));
 sky130_fd_sc_hd__dfxtp_1 _32591_ (.CLK(clk),
    .D(_04013_),
    .Q(\datamem.data_ram[21][22] ));
 sky130_fd_sc_hd__dfxtp_1 _32592_ (.CLK(clk),
    .D(_04014_),
    .Q(\datamem.data_ram[21][23] ));
 sky130_fd_sc_hd__dfxtp_1 _32593_ (.CLK(clk),
    .D(_04015_),
    .Q(\datamem.data_ram[21][8] ));
 sky130_fd_sc_hd__dfxtp_1 _32594_ (.CLK(clk),
    .D(_04016_),
    .Q(\datamem.data_ram[21][9] ));
 sky130_fd_sc_hd__dfxtp_1 _32595_ (.CLK(clk),
    .D(_04017_),
    .Q(\datamem.data_ram[21][10] ));
 sky130_fd_sc_hd__dfxtp_1 _32596_ (.CLK(clk),
    .D(_04018_),
    .Q(\datamem.data_ram[21][11] ));
 sky130_fd_sc_hd__dfxtp_1 _32597_ (.CLK(clk),
    .D(_04019_),
    .Q(\datamem.data_ram[21][12] ));
 sky130_fd_sc_hd__dfxtp_1 _32598_ (.CLK(clk),
    .D(_04020_),
    .Q(\datamem.data_ram[21][13] ));
 sky130_fd_sc_hd__dfxtp_1 _32599_ (.CLK(clk),
    .D(_04021_),
    .Q(\datamem.data_ram[21][14] ));
 sky130_fd_sc_hd__dfxtp_1 _32600_ (.CLK(clk),
    .D(_04022_),
    .Q(\datamem.data_ram[21][15] ));
 sky130_fd_sc_hd__dfxtp_1 _32601_ (.CLK(clk),
    .D(_04023_),
    .Q(\datamem.data_ram[20][24] ));
 sky130_fd_sc_hd__dfxtp_1 _32602_ (.CLK(clk),
    .D(_04024_),
    .Q(\datamem.data_ram[20][25] ));
 sky130_fd_sc_hd__dfxtp_1 _32603_ (.CLK(clk),
    .D(_04025_),
    .Q(\datamem.data_ram[20][26] ));
 sky130_fd_sc_hd__dfxtp_1 _32604_ (.CLK(clk),
    .D(_04026_),
    .Q(\datamem.data_ram[20][27] ));
 sky130_fd_sc_hd__dfxtp_1 _32605_ (.CLK(clk),
    .D(_04027_),
    .Q(\datamem.data_ram[20][28] ));
 sky130_fd_sc_hd__dfxtp_1 _32606_ (.CLK(clk),
    .D(_04028_),
    .Q(\datamem.data_ram[20][29] ));
 sky130_fd_sc_hd__dfxtp_1 _32607_ (.CLK(clk),
    .D(_04029_),
    .Q(\datamem.data_ram[20][30] ));
 sky130_fd_sc_hd__dfxtp_1 _32608_ (.CLK(clk),
    .D(_04030_),
    .Q(\datamem.data_ram[20][31] ));
 sky130_fd_sc_hd__dfxtp_1 _32609_ (.CLK(clk),
    .D(_04031_),
    .Q(\datamem.data_ram[20][16] ));
 sky130_fd_sc_hd__dfxtp_1 _32610_ (.CLK(clk),
    .D(_04032_),
    .Q(\datamem.data_ram[20][17] ));
 sky130_fd_sc_hd__dfxtp_1 _32611_ (.CLK(clk),
    .D(_04033_),
    .Q(\datamem.data_ram[20][18] ));
 sky130_fd_sc_hd__dfxtp_1 _32612_ (.CLK(clk),
    .D(_04034_),
    .Q(\datamem.data_ram[20][19] ));
 sky130_fd_sc_hd__dfxtp_1 _32613_ (.CLK(clk),
    .D(_04035_),
    .Q(\datamem.data_ram[20][20] ));
 sky130_fd_sc_hd__dfxtp_1 _32614_ (.CLK(clk),
    .D(_04036_),
    .Q(\datamem.data_ram[20][21] ));
 sky130_fd_sc_hd__dfxtp_1 _32615_ (.CLK(clk),
    .D(_04037_),
    .Q(\datamem.data_ram[20][22] ));
 sky130_fd_sc_hd__dfxtp_1 _32616_ (.CLK(clk),
    .D(_04038_),
    .Q(\datamem.data_ram[20][23] ));
 sky130_fd_sc_hd__dfxtp_1 _32617_ (.CLK(clk),
    .D(_04039_),
    .Q(\datamem.data_ram[20][8] ));
 sky130_fd_sc_hd__dfxtp_1 _32618_ (.CLK(clk),
    .D(_04040_),
    .Q(\datamem.data_ram[20][9] ));
 sky130_fd_sc_hd__dfxtp_1 _32619_ (.CLK(clk),
    .D(_04041_),
    .Q(\datamem.data_ram[20][10] ));
 sky130_fd_sc_hd__dfxtp_1 _32620_ (.CLK(clk),
    .D(_04042_),
    .Q(\datamem.data_ram[20][11] ));
 sky130_fd_sc_hd__dfxtp_1 _32621_ (.CLK(clk),
    .D(_04043_),
    .Q(\datamem.data_ram[20][12] ));
 sky130_fd_sc_hd__dfxtp_1 _32622_ (.CLK(clk),
    .D(_04044_),
    .Q(\datamem.data_ram[20][13] ));
 sky130_fd_sc_hd__dfxtp_1 _32623_ (.CLK(clk),
    .D(_04045_),
    .Q(\datamem.data_ram[20][14] ));
 sky130_fd_sc_hd__dfxtp_1 _32624_ (.CLK(clk),
    .D(_04046_),
    .Q(\datamem.data_ram[20][15] ));
 sky130_fd_sc_hd__dfxtp_1 _32625_ (.CLK(clk),
    .D(_04047_),
    .Q(\datamem.data_ram[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _32626_ (.CLK(clk),
    .D(_04048_),
    .Q(\datamem.data_ram[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _32627_ (.CLK(clk),
    .D(_04049_),
    .Q(\datamem.data_ram[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _32628_ (.CLK(clk),
    .D(_04050_),
    .Q(\datamem.data_ram[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _32629_ (.CLK(clk),
    .D(_04051_),
    .Q(\datamem.data_ram[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _32630_ (.CLK(clk),
    .D(_04052_),
    .Q(\datamem.data_ram[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _32631_ (.CLK(clk),
    .D(_04053_),
    .Q(\datamem.data_ram[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _32632_ (.CLK(clk),
    .D(_04054_),
    .Q(\datamem.data_ram[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _32633_ (.CLK(clk),
    .D(_04055_),
    .Q(\datamem.data_ram[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _32634_ (.CLK(clk),
    .D(_04056_),
    .Q(\datamem.data_ram[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _32635_ (.CLK(clk),
    .D(_04057_),
    .Q(\datamem.data_ram[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _32636_ (.CLK(clk),
    .D(_04058_),
    .Q(\datamem.data_ram[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _32637_ (.CLK(clk),
    .D(_04059_),
    .Q(\datamem.data_ram[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _32638_ (.CLK(clk),
    .D(_04060_),
    .Q(\datamem.data_ram[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _32639_ (.CLK(clk),
    .D(_04061_),
    .Q(\datamem.data_ram[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _32640_ (.CLK(clk),
    .D(_04062_),
    .Q(\datamem.data_ram[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _32641_ (.CLK(clk),
    .D(_04063_),
    .Q(\datamem.data_ram[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _32642_ (.CLK(clk),
    .D(_04064_),
    .Q(\datamem.data_ram[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _32643_ (.CLK(clk),
    .D(_04065_),
    .Q(\datamem.data_ram[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _32644_ (.CLK(clk),
    .D(_04066_),
    .Q(\datamem.data_ram[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _32645_ (.CLK(clk),
    .D(_04067_),
    .Q(\datamem.data_ram[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _32646_ (.CLK(clk),
    .D(_04068_),
    .Q(\datamem.data_ram[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _32647_ (.CLK(clk),
    .D(_04069_),
    .Q(\datamem.data_ram[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _32648_ (.CLK(clk),
    .D(_04070_),
    .Q(\datamem.data_ram[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _32649_ (.CLK(clk),
    .D(_04071_),
    .Q(\datamem.data_ram[19][24] ));
 sky130_fd_sc_hd__dfxtp_1 _32650_ (.CLK(clk),
    .D(_04072_),
    .Q(\datamem.data_ram[19][25] ));
 sky130_fd_sc_hd__dfxtp_1 _32651_ (.CLK(clk),
    .D(_04073_),
    .Q(\datamem.data_ram[19][26] ));
 sky130_fd_sc_hd__dfxtp_1 _32652_ (.CLK(clk),
    .D(_04074_),
    .Q(\datamem.data_ram[19][27] ));
 sky130_fd_sc_hd__dfxtp_1 _32653_ (.CLK(clk),
    .D(_04075_),
    .Q(\datamem.data_ram[19][28] ));
 sky130_fd_sc_hd__dfxtp_1 _32654_ (.CLK(clk),
    .D(_04076_),
    .Q(\datamem.data_ram[19][29] ));
 sky130_fd_sc_hd__dfxtp_1 _32655_ (.CLK(clk),
    .D(_04077_),
    .Q(\datamem.data_ram[19][30] ));
 sky130_fd_sc_hd__dfxtp_1 _32656_ (.CLK(clk),
    .D(_04078_),
    .Q(\datamem.data_ram[19][31] ));
 sky130_fd_sc_hd__dfxtp_1 _32657_ (.CLK(clk),
    .D(_04079_),
    .Q(\datamem.data_ram[19][16] ));
 sky130_fd_sc_hd__dfxtp_1 _32658_ (.CLK(clk),
    .D(_04080_),
    .Q(\datamem.data_ram[19][17] ));
 sky130_fd_sc_hd__dfxtp_1 _32659_ (.CLK(clk),
    .D(_04081_),
    .Q(\datamem.data_ram[19][18] ));
 sky130_fd_sc_hd__dfxtp_1 _32660_ (.CLK(clk),
    .D(_04082_),
    .Q(\datamem.data_ram[19][19] ));
 sky130_fd_sc_hd__dfxtp_1 _32661_ (.CLK(clk),
    .D(_04083_),
    .Q(\datamem.data_ram[19][20] ));
 sky130_fd_sc_hd__dfxtp_1 _32662_ (.CLK(clk),
    .D(_04084_),
    .Q(\datamem.data_ram[19][21] ));
 sky130_fd_sc_hd__dfxtp_1 _32663_ (.CLK(clk),
    .D(_04085_),
    .Q(\datamem.data_ram[19][22] ));
 sky130_fd_sc_hd__dfxtp_1 _32664_ (.CLK(clk),
    .D(_04086_),
    .Q(\datamem.data_ram[19][23] ));
 sky130_fd_sc_hd__dfxtp_1 _32665_ (.CLK(clk),
    .D(_04087_),
    .Q(\datamem.data_ram[19][8] ));
 sky130_fd_sc_hd__dfxtp_1 _32666_ (.CLK(clk),
    .D(_04088_),
    .Q(\datamem.data_ram[19][9] ));
 sky130_fd_sc_hd__dfxtp_1 _32667_ (.CLK(clk),
    .D(_04089_),
    .Q(\datamem.data_ram[19][10] ));
 sky130_fd_sc_hd__dfxtp_1 _32668_ (.CLK(clk),
    .D(_04090_),
    .Q(\datamem.data_ram[19][11] ));
 sky130_fd_sc_hd__dfxtp_1 _32669_ (.CLK(clk),
    .D(_04091_),
    .Q(\datamem.data_ram[19][12] ));
 sky130_fd_sc_hd__dfxtp_1 _32670_ (.CLK(clk),
    .D(_04092_),
    .Q(\datamem.data_ram[19][13] ));
 sky130_fd_sc_hd__dfxtp_1 _32671_ (.CLK(clk),
    .D(_04093_),
    .Q(\datamem.data_ram[19][14] ));
 sky130_fd_sc_hd__dfxtp_1 _32672_ (.CLK(clk),
    .D(_04094_),
    .Q(\datamem.data_ram[19][15] ));
 sky130_fd_sc_hd__dfxtp_1 _32673_ (.CLK(clk),
    .D(_04095_),
    .Q(\datamem.data_ram[18][24] ));
 sky130_fd_sc_hd__dfxtp_1 _32674_ (.CLK(clk),
    .D(_04096_),
    .Q(\datamem.data_ram[18][25] ));
 sky130_fd_sc_hd__dfxtp_1 _32675_ (.CLK(clk),
    .D(_04097_),
    .Q(\datamem.data_ram[18][26] ));
 sky130_fd_sc_hd__dfxtp_1 _32676_ (.CLK(clk),
    .D(_04098_),
    .Q(\datamem.data_ram[18][27] ));
 sky130_fd_sc_hd__dfxtp_1 _32677_ (.CLK(clk),
    .D(_04099_),
    .Q(\datamem.data_ram[18][28] ));
 sky130_fd_sc_hd__dfxtp_1 _32678_ (.CLK(clk),
    .D(_04100_),
    .Q(\datamem.data_ram[18][29] ));
 sky130_fd_sc_hd__dfxtp_1 _32679_ (.CLK(clk),
    .D(_04101_),
    .Q(\datamem.data_ram[18][30] ));
 sky130_fd_sc_hd__dfxtp_1 _32680_ (.CLK(clk),
    .D(_04102_),
    .Q(\datamem.data_ram[18][31] ));
 sky130_fd_sc_hd__dfxtp_1 _32681_ (.CLK(clk),
    .D(_04103_),
    .Q(\datamem.data_ram[18][16] ));
 sky130_fd_sc_hd__dfxtp_1 _32682_ (.CLK(clk),
    .D(_04104_),
    .Q(\datamem.data_ram[18][17] ));
 sky130_fd_sc_hd__dfxtp_1 _32683_ (.CLK(clk),
    .D(_04105_),
    .Q(\datamem.data_ram[18][18] ));
 sky130_fd_sc_hd__dfxtp_1 _32684_ (.CLK(clk),
    .D(_04106_),
    .Q(\datamem.data_ram[18][19] ));
 sky130_fd_sc_hd__dfxtp_1 _32685_ (.CLK(clk),
    .D(_04107_),
    .Q(\datamem.data_ram[18][20] ));
 sky130_fd_sc_hd__dfxtp_1 _32686_ (.CLK(clk),
    .D(_04108_),
    .Q(\datamem.data_ram[18][21] ));
 sky130_fd_sc_hd__dfxtp_1 _32687_ (.CLK(clk),
    .D(_04109_),
    .Q(\datamem.data_ram[18][22] ));
 sky130_fd_sc_hd__dfxtp_1 _32688_ (.CLK(clk),
    .D(_04110_),
    .Q(\datamem.data_ram[18][23] ));
 sky130_fd_sc_hd__dfxtp_1 _32689_ (.CLK(clk),
    .D(_04111_),
    .Q(\datamem.data_ram[18][8] ));
 sky130_fd_sc_hd__dfxtp_1 _32690_ (.CLK(clk),
    .D(_04112_),
    .Q(\datamem.data_ram[18][9] ));
 sky130_fd_sc_hd__dfxtp_1 _32691_ (.CLK(clk),
    .D(_04113_),
    .Q(\datamem.data_ram[18][10] ));
 sky130_fd_sc_hd__dfxtp_1 _32692_ (.CLK(clk),
    .D(_04114_),
    .Q(\datamem.data_ram[18][11] ));
 sky130_fd_sc_hd__dfxtp_1 _32693_ (.CLK(clk),
    .D(_04115_),
    .Q(\datamem.data_ram[18][12] ));
 sky130_fd_sc_hd__dfxtp_1 _32694_ (.CLK(clk),
    .D(_04116_),
    .Q(\datamem.data_ram[18][13] ));
 sky130_fd_sc_hd__dfxtp_1 _32695_ (.CLK(clk),
    .D(_04117_),
    .Q(\datamem.data_ram[18][14] ));
 sky130_fd_sc_hd__dfxtp_1 _32696_ (.CLK(clk),
    .D(_04118_),
    .Q(\datamem.data_ram[18][15] ));
 sky130_fd_sc_hd__dfxtp_1 _32697_ (.CLK(clk),
    .D(_04119_),
    .Q(\datamem.data_ram[17][24] ));
 sky130_fd_sc_hd__dfxtp_1 _32698_ (.CLK(clk),
    .D(_04120_),
    .Q(\datamem.data_ram[17][25] ));
 sky130_fd_sc_hd__dfxtp_1 _32699_ (.CLK(clk),
    .D(_04121_),
    .Q(\datamem.data_ram[17][26] ));
 sky130_fd_sc_hd__dfxtp_1 _32700_ (.CLK(clk),
    .D(_04122_),
    .Q(\datamem.data_ram[17][27] ));
 sky130_fd_sc_hd__dfxtp_1 _32701_ (.CLK(clk),
    .D(_04123_),
    .Q(\datamem.data_ram[17][28] ));
 sky130_fd_sc_hd__dfxtp_1 _32702_ (.CLK(clk),
    .D(_04124_),
    .Q(\datamem.data_ram[17][29] ));
 sky130_fd_sc_hd__dfxtp_1 _32703_ (.CLK(clk),
    .D(_04125_),
    .Q(\datamem.data_ram[17][30] ));
 sky130_fd_sc_hd__dfxtp_1 _32704_ (.CLK(clk),
    .D(_04126_),
    .Q(\datamem.data_ram[17][31] ));
 sky130_fd_sc_hd__dfxtp_1 _32705_ (.CLK(clk),
    .D(_04127_),
    .Q(\datamem.data_ram[17][16] ));
 sky130_fd_sc_hd__dfxtp_1 _32706_ (.CLK(clk),
    .D(_04128_),
    .Q(\datamem.data_ram[17][17] ));
 sky130_fd_sc_hd__dfxtp_1 _32707_ (.CLK(clk),
    .D(_04129_),
    .Q(\datamem.data_ram[17][18] ));
 sky130_fd_sc_hd__dfxtp_1 _32708_ (.CLK(clk),
    .D(_04130_),
    .Q(\datamem.data_ram[17][19] ));
 sky130_fd_sc_hd__dfxtp_1 _32709_ (.CLK(clk),
    .D(_04131_),
    .Q(\datamem.data_ram[17][20] ));
 sky130_fd_sc_hd__dfxtp_1 _32710_ (.CLK(clk),
    .D(_04132_),
    .Q(\datamem.data_ram[17][21] ));
 sky130_fd_sc_hd__dfxtp_1 _32711_ (.CLK(clk),
    .D(_04133_),
    .Q(\datamem.data_ram[17][22] ));
 sky130_fd_sc_hd__dfxtp_1 _32712_ (.CLK(clk),
    .D(_04134_),
    .Q(\datamem.data_ram[17][23] ));
 sky130_fd_sc_hd__dfxtp_1 _32713_ (.CLK(clk),
    .D(_04135_),
    .Q(\datamem.data_ram[17][8] ));
 sky130_fd_sc_hd__dfxtp_1 _32714_ (.CLK(clk),
    .D(_04136_),
    .Q(\datamem.data_ram[17][9] ));
 sky130_fd_sc_hd__dfxtp_1 _32715_ (.CLK(clk),
    .D(_04137_),
    .Q(\datamem.data_ram[17][10] ));
 sky130_fd_sc_hd__dfxtp_1 _32716_ (.CLK(clk),
    .D(_04138_),
    .Q(\datamem.data_ram[17][11] ));
 sky130_fd_sc_hd__dfxtp_1 _32717_ (.CLK(clk),
    .D(_04139_),
    .Q(\datamem.data_ram[17][12] ));
 sky130_fd_sc_hd__dfxtp_1 _32718_ (.CLK(clk),
    .D(_04140_),
    .Q(\datamem.data_ram[17][13] ));
 sky130_fd_sc_hd__dfxtp_1 _32719_ (.CLK(clk),
    .D(_04141_),
    .Q(\datamem.data_ram[17][14] ));
 sky130_fd_sc_hd__dfxtp_1 _32720_ (.CLK(clk),
    .D(_04142_),
    .Q(\datamem.data_ram[17][15] ));
 sky130_fd_sc_hd__dfxtp_1 _32721_ (.CLK(clk),
    .D(_04143_),
    .Q(\datamem.data_ram[16][24] ));
 sky130_fd_sc_hd__dfxtp_1 _32722_ (.CLK(clk),
    .D(_04144_),
    .Q(\datamem.data_ram[16][25] ));
 sky130_fd_sc_hd__dfxtp_1 _32723_ (.CLK(clk),
    .D(_04145_),
    .Q(\datamem.data_ram[16][26] ));
 sky130_fd_sc_hd__dfxtp_1 _32724_ (.CLK(clk),
    .D(_04146_),
    .Q(\datamem.data_ram[16][27] ));
 sky130_fd_sc_hd__dfxtp_1 _32725_ (.CLK(clk),
    .D(_04147_),
    .Q(\datamem.data_ram[16][28] ));
 sky130_fd_sc_hd__dfxtp_1 _32726_ (.CLK(clk),
    .D(_04148_),
    .Q(\datamem.data_ram[16][29] ));
 sky130_fd_sc_hd__dfxtp_1 _32727_ (.CLK(clk),
    .D(_04149_),
    .Q(\datamem.data_ram[16][30] ));
 sky130_fd_sc_hd__dfxtp_1 _32728_ (.CLK(clk),
    .D(_04150_),
    .Q(\datamem.data_ram[16][31] ));
 sky130_fd_sc_hd__dfxtp_1 _32729_ (.CLK(clk),
    .D(_04151_),
    .Q(\datamem.data_ram[16][16] ));
 sky130_fd_sc_hd__dfxtp_1 _32730_ (.CLK(clk),
    .D(_04152_),
    .Q(\datamem.data_ram[16][17] ));
 sky130_fd_sc_hd__dfxtp_1 _32731_ (.CLK(clk),
    .D(_04153_),
    .Q(\datamem.data_ram[16][18] ));
 sky130_fd_sc_hd__dfxtp_1 _32732_ (.CLK(clk),
    .D(_04154_),
    .Q(\datamem.data_ram[16][19] ));
 sky130_fd_sc_hd__dfxtp_1 _32733_ (.CLK(clk),
    .D(_04155_),
    .Q(\datamem.data_ram[16][20] ));
 sky130_fd_sc_hd__dfxtp_1 _32734_ (.CLK(clk),
    .D(_04156_),
    .Q(\datamem.data_ram[16][21] ));
 sky130_fd_sc_hd__dfxtp_1 _32735_ (.CLK(clk),
    .D(_04157_),
    .Q(\datamem.data_ram[16][22] ));
 sky130_fd_sc_hd__dfxtp_1 _32736_ (.CLK(clk),
    .D(_04158_),
    .Q(\datamem.data_ram[16][23] ));
 sky130_fd_sc_hd__dfxtp_1 _32737_ (.CLK(clk),
    .D(_04159_),
    .Q(\datamem.data_ram[16][8] ));
 sky130_fd_sc_hd__dfxtp_1 _32738_ (.CLK(clk),
    .D(_04160_),
    .Q(\datamem.data_ram[16][9] ));
 sky130_fd_sc_hd__dfxtp_1 _32739_ (.CLK(clk),
    .D(_04161_),
    .Q(\datamem.data_ram[16][10] ));
 sky130_fd_sc_hd__dfxtp_1 _32740_ (.CLK(clk),
    .D(_04162_),
    .Q(\datamem.data_ram[16][11] ));
 sky130_fd_sc_hd__dfxtp_1 _32741_ (.CLK(clk),
    .D(_04163_),
    .Q(\datamem.data_ram[16][12] ));
 sky130_fd_sc_hd__dfxtp_1 _32742_ (.CLK(clk),
    .D(_04164_),
    .Q(\datamem.data_ram[16][13] ));
 sky130_fd_sc_hd__dfxtp_1 _32743_ (.CLK(clk),
    .D(_04165_),
    .Q(\datamem.data_ram[16][14] ));
 sky130_fd_sc_hd__dfxtp_1 _32744_ (.CLK(clk),
    .D(_04166_),
    .Q(\datamem.data_ram[16][15] ));
 sky130_fd_sc_hd__dfxtp_1 _32745_ (.CLK(clk),
    .D(_04167_),
    .Q(\datamem.data_ram[15][24] ));
 sky130_fd_sc_hd__dfxtp_1 _32746_ (.CLK(clk),
    .D(_04168_),
    .Q(\datamem.data_ram[15][25] ));
 sky130_fd_sc_hd__dfxtp_1 _32747_ (.CLK(clk),
    .D(_04169_),
    .Q(\datamem.data_ram[15][26] ));
 sky130_fd_sc_hd__dfxtp_1 _32748_ (.CLK(clk),
    .D(_04170_),
    .Q(\datamem.data_ram[15][27] ));
 sky130_fd_sc_hd__dfxtp_1 _32749_ (.CLK(clk),
    .D(_04171_),
    .Q(\datamem.data_ram[15][28] ));
 sky130_fd_sc_hd__dfxtp_1 _32750_ (.CLK(clk),
    .D(_04172_),
    .Q(\datamem.data_ram[15][29] ));
 sky130_fd_sc_hd__dfxtp_1 _32751_ (.CLK(clk),
    .D(_04173_),
    .Q(\datamem.data_ram[15][30] ));
 sky130_fd_sc_hd__dfxtp_1 _32752_ (.CLK(clk),
    .D(_04174_),
    .Q(\datamem.data_ram[15][31] ));
 sky130_fd_sc_hd__dfxtp_1 _32753_ (.CLK(clk),
    .D(_04175_),
    .Q(\datamem.data_ram[15][16] ));
 sky130_fd_sc_hd__dfxtp_1 _32754_ (.CLK(clk),
    .D(_04176_),
    .Q(\datamem.data_ram[15][17] ));
 sky130_fd_sc_hd__dfxtp_1 _32755_ (.CLK(clk),
    .D(_04177_),
    .Q(\datamem.data_ram[15][18] ));
 sky130_fd_sc_hd__dfxtp_1 _32756_ (.CLK(clk),
    .D(_04178_),
    .Q(\datamem.data_ram[15][19] ));
 sky130_fd_sc_hd__dfxtp_1 _32757_ (.CLK(clk),
    .D(_04179_),
    .Q(\datamem.data_ram[15][20] ));
 sky130_fd_sc_hd__dfxtp_1 _32758_ (.CLK(clk),
    .D(_04180_),
    .Q(\datamem.data_ram[15][21] ));
 sky130_fd_sc_hd__dfxtp_1 _32759_ (.CLK(clk),
    .D(_04181_),
    .Q(\datamem.data_ram[15][22] ));
 sky130_fd_sc_hd__dfxtp_1 _32760_ (.CLK(clk),
    .D(_04182_),
    .Q(\datamem.data_ram[15][23] ));
 sky130_fd_sc_hd__dfxtp_1 _32761_ (.CLK(clk),
    .D(_04183_),
    .Q(\datamem.data_ram[15][8] ));
 sky130_fd_sc_hd__dfxtp_1 _32762_ (.CLK(clk),
    .D(_04184_),
    .Q(\datamem.data_ram[15][9] ));
 sky130_fd_sc_hd__dfxtp_1 _32763_ (.CLK(clk),
    .D(_04185_),
    .Q(\datamem.data_ram[15][10] ));
 sky130_fd_sc_hd__dfxtp_1 _32764_ (.CLK(clk),
    .D(_04186_),
    .Q(\datamem.data_ram[15][11] ));
 sky130_fd_sc_hd__dfxtp_1 _32765_ (.CLK(clk),
    .D(_04187_),
    .Q(\datamem.data_ram[15][12] ));
 sky130_fd_sc_hd__dfxtp_1 _32766_ (.CLK(clk),
    .D(_04188_),
    .Q(\datamem.data_ram[15][13] ));
 sky130_fd_sc_hd__dfxtp_1 _32767_ (.CLK(clk),
    .D(_04189_),
    .Q(\datamem.data_ram[15][14] ));
 sky130_fd_sc_hd__dfxtp_1 _32768_ (.CLK(clk),
    .D(_04190_),
    .Q(\datamem.data_ram[15][15] ));
 sky130_fd_sc_hd__dfxtp_1 _32769_ (.CLK(clk),
    .D(_04191_),
    .Q(\datamem.data_ram[14][24] ));
 sky130_fd_sc_hd__dfxtp_1 _32770_ (.CLK(clk),
    .D(_04192_),
    .Q(\datamem.data_ram[14][25] ));
 sky130_fd_sc_hd__dfxtp_1 _32771_ (.CLK(clk),
    .D(_04193_),
    .Q(\datamem.data_ram[14][26] ));
 sky130_fd_sc_hd__dfxtp_1 _32772_ (.CLK(clk),
    .D(_04194_),
    .Q(\datamem.data_ram[14][27] ));
 sky130_fd_sc_hd__dfxtp_1 _32773_ (.CLK(clk),
    .D(_04195_),
    .Q(\datamem.data_ram[14][28] ));
 sky130_fd_sc_hd__dfxtp_1 _32774_ (.CLK(clk),
    .D(_04196_),
    .Q(\datamem.data_ram[14][29] ));
 sky130_fd_sc_hd__dfxtp_1 _32775_ (.CLK(clk),
    .D(_04197_),
    .Q(\datamem.data_ram[14][30] ));
 sky130_fd_sc_hd__dfxtp_1 _32776_ (.CLK(clk),
    .D(_04198_),
    .Q(\datamem.data_ram[14][31] ));
 sky130_fd_sc_hd__dfxtp_1 _32777_ (.CLK(clk),
    .D(_04199_),
    .Q(\datamem.data_ram[14][16] ));
 sky130_fd_sc_hd__dfxtp_1 _32778_ (.CLK(clk),
    .D(_04200_),
    .Q(\datamem.data_ram[14][17] ));
 sky130_fd_sc_hd__dfxtp_1 _32779_ (.CLK(clk),
    .D(_04201_),
    .Q(\datamem.data_ram[14][18] ));
 sky130_fd_sc_hd__dfxtp_1 _32780_ (.CLK(clk),
    .D(_04202_),
    .Q(\datamem.data_ram[14][19] ));
 sky130_fd_sc_hd__dfxtp_1 _32781_ (.CLK(clk),
    .D(_04203_),
    .Q(\datamem.data_ram[14][20] ));
 sky130_fd_sc_hd__dfxtp_1 _32782_ (.CLK(clk),
    .D(_04204_),
    .Q(\datamem.data_ram[14][21] ));
 sky130_fd_sc_hd__dfxtp_1 _32783_ (.CLK(clk),
    .D(_04205_),
    .Q(\datamem.data_ram[14][22] ));
 sky130_fd_sc_hd__dfxtp_1 _32784_ (.CLK(clk),
    .D(_04206_),
    .Q(\datamem.data_ram[14][23] ));
 sky130_fd_sc_hd__dfxtp_1 _32785_ (.CLK(clk),
    .D(_04207_),
    .Q(\datamem.data_ram[14][8] ));
 sky130_fd_sc_hd__dfxtp_1 _32786_ (.CLK(clk),
    .D(_04208_),
    .Q(\datamem.data_ram[14][9] ));
 sky130_fd_sc_hd__dfxtp_1 _32787_ (.CLK(clk),
    .D(_04209_),
    .Q(\datamem.data_ram[14][10] ));
 sky130_fd_sc_hd__dfxtp_1 _32788_ (.CLK(clk),
    .D(_04210_),
    .Q(\datamem.data_ram[14][11] ));
 sky130_fd_sc_hd__dfxtp_1 _32789_ (.CLK(clk),
    .D(_04211_),
    .Q(\datamem.data_ram[14][12] ));
 sky130_fd_sc_hd__dfxtp_1 _32790_ (.CLK(clk),
    .D(_04212_),
    .Q(\datamem.data_ram[14][13] ));
 sky130_fd_sc_hd__dfxtp_1 _32791_ (.CLK(clk),
    .D(_04213_),
    .Q(\datamem.data_ram[14][14] ));
 sky130_fd_sc_hd__dfxtp_1 _32792_ (.CLK(clk),
    .D(_04214_),
    .Q(\datamem.data_ram[14][15] ));
 sky130_fd_sc_hd__dfxtp_1 _32793_ (.CLK(clk),
    .D(_04215_),
    .Q(\datamem.data_ram[13][24] ));
 sky130_fd_sc_hd__dfxtp_1 _32794_ (.CLK(clk),
    .D(_04216_),
    .Q(\datamem.data_ram[13][25] ));
 sky130_fd_sc_hd__dfxtp_1 _32795_ (.CLK(clk),
    .D(_04217_),
    .Q(\datamem.data_ram[13][26] ));
 sky130_fd_sc_hd__dfxtp_1 _32796_ (.CLK(clk),
    .D(_04218_),
    .Q(\datamem.data_ram[13][27] ));
 sky130_fd_sc_hd__dfxtp_1 _32797_ (.CLK(clk),
    .D(_04219_),
    .Q(\datamem.data_ram[13][28] ));
 sky130_fd_sc_hd__dfxtp_1 _32798_ (.CLK(clk),
    .D(_04220_),
    .Q(\datamem.data_ram[13][29] ));
 sky130_fd_sc_hd__dfxtp_1 _32799_ (.CLK(clk),
    .D(_04221_),
    .Q(\datamem.data_ram[13][30] ));
 sky130_fd_sc_hd__dfxtp_1 _32800_ (.CLK(clk),
    .D(_04222_),
    .Q(\datamem.data_ram[13][31] ));
 sky130_fd_sc_hd__dfxtp_1 _32801_ (.CLK(clk),
    .D(_04223_),
    .Q(\datamem.data_ram[13][16] ));
 sky130_fd_sc_hd__dfxtp_1 _32802_ (.CLK(clk),
    .D(_04224_),
    .Q(\datamem.data_ram[13][17] ));
 sky130_fd_sc_hd__dfxtp_1 _32803_ (.CLK(clk),
    .D(_04225_),
    .Q(\datamem.data_ram[13][18] ));
 sky130_fd_sc_hd__dfxtp_1 _32804_ (.CLK(clk),
    .D(_04226_),
    .Q(\datamem.data_ram[13][19] ));
 sky130_fd_sc_hd__dfxtp_1 _32805_ (.CLK(clk),
    .D(_04227_),
    .Q(\datamem.data_ram[13][20] ));
 sky130_fd_sc_hd__dfxtp_1 _32806_ (.CLK(clk),
    .D(_04228_),
    .Q(\datamem.data_ram[13][21] ));
 sky130_fd_sc_hd__dfxtp_1 _32807_ (.CLK(clk),
    .D(_04229_),
    .Q(\datamem.data_ram[13][22] ));
 sky130_fd_sc_hd__dfxtp_1 _32808_ (.CLK(clk),
    .D(_04230_),
    .Q(\datamem.data_ram[13][23] ));
 sky130_fd_sc_hd__dfxtp_1 _32809_ (.CLK(clk),
    .D(_04231_),
    .Q(\datamem.data_ram[13][8] ));
 sky130_fd_sc_hd__dfxtp_1 _32810_ (.CLK(clk),
    .D(_04232_),
    .Q(\datamem.data_ram[13][9] ));
 sky130_fd_sc_hd__dfxtp_1 _32811_ (.CLK(clk),
    .D(_04233_),
    .Q(\datamem.data_ram[13][10] ));
 sky130_fd_sc_hd__dfxtp_1 _32812_ (.CLK(clk),
    .D(_04234_),
    .Q(\datamem.data_ram[13][11] ));
 sky130_fd_sc_hd__dfxtp_1 _32813_ (.CLK(clk),
    .D(_04235_),
    .Q(\datamem.data_ram[13][12] ));
 sky130_fd_sc_hd__dfxtp_1 _32814_ (.CLK(clk),
    .D(_04236_),
    .Q(\datamem.data_ram[13][13] ));
 sky130_fd_sc_hd__dfxtp_1 _32815_ (.CLK(clk),
    .D(_04237_),
    .Q(\datamem.data_ram[13][14] ));
 sky130_fd_sc_hd__dfxtp_1 _32816_ (.CLK(clk),
    .D(_04238_),
    .Q(\datamem.data_ram[13][15] ));
 sky130_fd_sc_hd__dfxtp_1 _32817_ (.CLK(clk),
    .D(_04239_),
    .Q(\datamem.data_ram[12][24] ));
 sky130_fd_sc_hd__dfxtp_1 _32818_ (.CLK(clk),
    .D(_04240_),
    .Q(\datamem.data_ram[12][25] ));
 sky130_fd_sc_hd__dfxtp_1 _32819_ (.CLK(clk),
    .D(_04241_),
    .Q(\datamem.data_ram[12][26] ));
 sky130_fd_sc_hd__dfxtp_1 _32820_ (.CLK(clk),
    .D(_04242_),
    .Q(\datamem.data_ram[12][27] ));
 sky130_fd_sc_hd__dfxtp_1 _32821_ (.CLK(clk),
    .D(_04243_),
    .Q(\datamem.data_ram[12][28] ));
 sky130_fd_sc_hd__dfxtp_1 _32822_ (.CLK(clk),
    .D(_04244_),
    .Q(\datamem.data_ram[12][29] ));
 sky130_fd_sc_hd__dfxtp_1 _32823_ (.CLK(clk),
    .D(_04245_),
    .Q(\datamem.data_ram[12][30] ));
 sky130_fd_sc_hd__dfxtp_1 _32824_ (.CLK(clk),
    .D(_04246_),
    .Q(\datamem.data_ram[12][31] ));
 sky130_fd_sc_hd__dfxtp_1 _32825_ (.CLK(clk),
    .D(_04247_),
    .Q(\datamem.data_ram[12][16] ));
 sky130_fd_sc_hd__dfxtp_1 _32826_ (.CLK(clk),
    .D(_04248_),
    .Q(\datamem.data_ram[12][17] ));
 sky130_fd_sc_hd__dfxtp_1 _32827_ (.CLK(clk),
    .D(_04249_),
    .Q(\datamem.data_ram[12][18] ));
 sky130_fd_sc_hd__dfxtp_1 _32828_ (.CLK(clk),
    .D(_04250_),
    .Q(\datamem.data_ram[12][19] ));
 sky130_fd_sc_hd__dfxtp_1 _32829_ (.CLK(clk),
    .D(_04251_),
    .Q(\datamem.data_ram[12][20] ));
 sky130_fd_sc_hd__dfxtp_1 _32830_ (.CLK(clk),
    .D(_04252_),
    .Q(\datamem.data_ram[12][21] ));
 sky130_fd_sc_hd__dfxtp_1 _32831_ (.CLK(clk),
    .D(_04253_),
    .Q(\datamem.data_ram[12][22] ));
 sky130_fd_sc_hd__dfxtp_1 _32832_ (.CLK(clk),
    .D(_04254_),
    .Q(\datamem.data_ram[12][23] ));
 sky130_fd_sc_hd__dfxtp_1 _32833_ (.CLK(clk),
    .D(_04255_),
    .Q(\datamem.data_ram[12][8] ));
 sky130_fd_sc_hd__dfxtp_1 _32834_ (.CLK(clk),
    .D(_04256_),
    .Q(\datamem.data_ram[12][9] ));
 sky130_fd_sc_hd__dfxtp_1 _32835_ (.CLK(clk),
    .D(_04257_),
    .Q(\datamem.data_ram[12][10] ));
 sky130_fd_sc_hd__dfxtp_1 _32836_ (.CLK(clk),
    .D(_04258_),
    .Q(\datamem.data_ram[12][11] ));
 sky130_fd_sc_hd__dfxtp_1 _32837_ (.CLK(clk),
    .D(_04259_),
    .Q(\datamem.data_ram[12][12] ));
 sky130_fd_sc_hd__dfxtp_1 _32838_ (.CLK(clk),
    .D(_04260_),
    .Q(\datamem.data_ram[12][13] ));
 sky130_fd_sc_hd__dfxtp_1 _32839_ (.CLK(clk),
    .D(_04261_),
    .Q(\datamem.data_ram[12][14] ));
 sky130_fd_sc_hd__dfxtp_1 _32840_ (.CLK(clk),
    .D(_04262_),
    .Q(\datamem.data_ram[12][15] ));
 sky130_fd_sc_hd__dfxtp_1 _32841_ (.CLK(clk),
    .D(_04263_),
    .Q(\datamem.data_ram[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _32842_ (.CLK(clk),
    .D(_04264_),
    .Q(\datamem.data_ram[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _32843_ (.CLK(clk),
    .D(_04265_),
    .Q(\datamem.data_ram[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _32844_ (.CLK(clk),
    .D(_04266_),
    .Q(\datamem.data_ram[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _32845_ (.CLK(clk),
    .D(_04267_),
    .Q(\datamem.data_ram[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _32846_ (.CLK(clk),
    .D(_04268_),
    .Q(\datamem.data_ram[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _32847_ (.CLK(clk),
    .D(_04269_),
    .Q(\datamem.data_ram[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _32848_ (.CLK(clk),
    .D(_04270_),
    .Q(\datamem.data_ram[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _32849_ (.CLK(clk),
    .D(_04271_),
    .Q(\datamem.data_ram[11][24] ));
 sky130_fd_sc_hd__dfxtp_1 _32850_ (.CLK(clk),
    .D(_04272_),
    .Q(\datamem.data_ram[11][25] ));
 sky130_fd_sc_hd__dfxtp_1 _32851_ (.CLK(clk),
    .D(_04273_),
    .Q(\datamem.data_ram[11][26] ));
 sky130_fd_sc_hd__dfxtp_1 _32852_ (.CLK(clk),
    .D(_04274_),
    .Q(\datamem.data_ram[11][27] ));
 sky130_fd_sc_hd__dfxtp_1 _32853_ (.CLK(clk),
    .D(_04275_),
    .Q(\datamem.data_ram[11][28] ));
 sky130_fd_sc_hd__dfxtp_1 _32854_ (.CLK(clk),
    .D(_04276_),
    .Q(\datamem.data_ram[11][29] ));
 sky130_fd_sc_hd__dfxtp_1 _32855_ (.CLK(clk),
    .D(_04277_),
    .Q(\datamem.data_ram[11][30] ));
 sky130_fd_sc_hd__dfxtp_1 _32856_ (.CLK(clk),
    .D(_04278_),
    .Q(\datamem.data_ram[11][31] ));
 sky130_fd_sc_hd__dfxtp_1 _32857_ (.CLK(clk),
    .D(_04279_),
    .Q(\datamem.data_ram[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _32858_ (.CLK(clk),
    .D(_04280_),
    .Q(\datamem.data_ram[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _32859_ (.CLK(clk),
    .D(_04281_),
    .Q(\datamem.data_ram[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _32860_ (.CLK(clk),
    .D(_04282_),
    .Q(\datamem.data_ram[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _32861_ (.CLK(clk),
    .D(_04283_),
    .Q(\datamem.data_ram[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _32862_ (.CLK(clk),
    .D(_04284_),
    .Q(\datamem.data_ram[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _32863_ (.CLK(clk),
    .D(_04285_),
    .Q(\datamem.data_ram[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _32864_ (.CLK(clk),
    .D(_04286_),
    .Q(\datamem.data_ram[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _32865_ (.CLK(clk),
    .D(_04287_),
    .Q(\datamem.data_ram[11][8] ));
 sky130_fd_sc_hd__dfxtp_1 _32866_ (.CLK(clk),
    .D(_04288_),
    .Q(\datamem.data_ram[11][9] ));
 sky130_fd_sc_hd__dfxtp_1 _32867_ (.CLK(clk),
    .D(_04289_),
    .Q(\datamem.data_ram[11][10] ));
 sky130_fd_sc_hd__dfxtp_1 _32868_ (.CLK(clk),
    .D(_04290_),
    .Q(\datamem.data_ram[11][11] ));
 sky130_fd_sc_hd__dfxtp_1 _32869_ (.CLK(clk),
    .D(_04291_),
    .Q(\datamem.data_ram[11][12] ));
 sky130_fd_sc_hd__dfxtp_1 _32870_ (.CLK(clk),
    .D(_04292_),
    .Q(\datamem.data_ram[11][13] ));
 sky130_fd_sc_hd__dfxtp_1 _32871_ (.CLK(clk),
    .D(_04293_),
    .Q(\datamem.data_ram[11][14] ));
 sky130_fd_sc_hd__dfxtp_1 _32872_ (.CLK(clk),
    .D(_04294_),
    .Q(\datamem.data_ram[11][15] ));
 sky130_fd_sc_hd__dfxtp_1 _32873_ (.CLK(clk),
    .D(_04295_),
    .Q(\datamem.data_ram[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _32874_ (.CLK(clk),
    .D(_04296_),
    .Q(\datamem.data_ram[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _32875_ (.CLK(clk),
    .D(_04297_),
    .Q(\datamem.data_ram[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _32876_ (.CLK(clk),
    .D(_04298_),
    .Q(\datamem.data_ram[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _32877_ (.CLK(clk),
    .D(_04299_),
    .Q(\datamem.data_ram[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _32878_ (.CLK(clk),
    .D(_04300_),
    .Q(\datamem.data_ram[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _32879_ (.CLK(clk),
    .D(_04301_),
    .Q(\datamem.data_ram[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _32880_ (.CLK(clk),
    .D(_04302_),
    .Q(\datamem.data_ram[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _32881_ (.CLK(clk),
    .D(_04303_),
    .Q(\datamem.data_ram[10][8] ));
 sky130_fd_sc_hd__dfxtp_1 _32882_ (.CLK(clk),
    .D(_04304_),
    .Q(\datamem.data_ram[10][9] ));
 sky130_fd_sc_hd__dfxtp_1 _32883_ (.CLK(clk),
    .D(_04305_),
    .Q(\datamem.data_ram[10][10] ));
 sky130_fd_sc_hd__dfxtp_1 _32884_ (.CLK(clk),
    .D(_04306_),
    .Q(\datamem.data_ram[10][11] ));
 sky130_fd_sc_hd__dfxtp_1 _32885_ (.CLK(clk),
    .D(_04307_),
    .Q(\datamem.data_ram[10][12] ));
 sky130_fd_sc_hd__dfxtp_1 _32886_ (.CLK(clk),
    .D(_04308_),
    .Q(\datamem.data_ram[10][13] ));
 sky130_fd_sc_hd__dfxtp_1 _32887_ (.CLK(clk),
    .D(_04309_),
    .Q(\datamem.data_ram[10][14] ));
 sky130_fd_sc_hd__dfxtp_1 _32888_ (.CLK(clk),
    .D(_04310_),
    .Q(\datamem.data_ram[10][15] ));
 sky130_fd_sc_hd__dfxtp_1 _32889_ (.CLK(clk),
    .D(_04311_),
    .Q(\datamem.data_ram[10][16] ));
 sky130_fd_sc_hd__dfxtp_1 _32890_ (.CLK(clk),
    .D(_04312_),
    .Q(\datamem.data_ram[10][17] ));
 sky130_fd_sc_hd__dfxtp_1 _32891_ (.CLK(clk),
    .D(_04313_),
    .Q(\datamem.data_ram[10][18] ));
 sky130_fd_sc_hd__dfxtp_1 _32892_ (.CLK(clk),
    .D(_04314_),
    .Q(\datamem.data_ram[10][19] ));
 sky130_fd_sc_hd__dfxtp_1 _32893_ (.CLK(clk),
    .D(_04315_),
    .Q(\datamem.data_ram[10][20] ));
 sky130_fd_sc_hd__dfxtp_1 _32894_ (.CLK(clk),
    .D(_04316_),
    .Q(\datamem.data_ram[10][21] ));
 sky130_fd_sc_hd__dfxtp_1 _32895_ (.CLK(clk),
    .D(_04317_),
    .Q(\datamem.data_ram[10][22] ));
 sky130_fd_sc_hd__dfxtp_1 _32896_ (.CLK(clk),
    .D(_04318_),
    .Q(\datamem.data_ram[10][23] ));
 sky130_fd_sc_hd__dfxtp_1 _32897_ (.CLK(clk),
    .D(_04319_),
    .Q(\datamem.data_ram[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _32898_ (.CLK(clk),
    .D(_04320_),
    .Q(\datamem.data_ram[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _32899_ (.CLK(clk),
    .D(_04321_),
    .Q(\datamem.data_ram[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _32900_ (.CLK(clk),
    .D(_04322_),
    .Q(\datamem.data_ram[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _32901_ (.CLK(clk),
    .D(_04323_),
    .Q(\datamem.data_ram[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _32902_ (.CLK(clk),
    .D(_04324_),
    .Q(\datamem.data_ram[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _32903_ (.CLK(clk),
    .D(_04325_),
    .Q(\datamem.data_ram[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _32904_ (.CLK(clk),
    .D(_04326_),
    .Q(\datamem.data_ram[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _32905_ (.CLK(clk),
    .D(_04327_),
    .Q(\datamem.data_ram[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _32906_ (.CLK(clk),
    .D(_04328_),
    .Q(\datamem.data_ram[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _32907_ (.CLK(clk),
    .D(_04329_),
    .Q(\datamem.data_ram[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _32908_ (.CLK(clk),
    .D(_04330_),
    .Q(\datamem.data_ram[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _32909_ (.CLK(clk),
    .D(_04331_),
    .Q(\datamem.data_ram[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _32910_ (.CLK(clk),
    .D(_04332_),
    .Q(\datamem.data_ram[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _32911_ (.CLK(clk),
    .D(_04333_),
    .Q(\datamem.data_ram[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _32912_ (.CLK(clk),
    .D(_04334_),
    .Q(\datamem.data_ram[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 _32913_ (.CLK(clk),
    .D(_04335_),
    .Q(\datamem.data_ram[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _32914_ (.CLK(clk),
    .D(_04336_),
    .Q(\datamem.data_ram[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _32915_ (.CLK(clk),
    .D(_04337_),
    .Q(\datamem.data_ram[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _32916_ (.CLK(clk),
    .D(_04338_),
    .Q(\datamem.data_ram[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _32917_ (.CLK(clk),
    .D(_04339_),
    .Q(\datamem.data_ram[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _32918_ (.CLK(clk),
    .D(_04340_),
    .Q(\datamem.data_ram[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _32919_ (.CLK(clk),
    .D(_04341_),
    .Q(\datamem.data_ram[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _32920_ (.CLK(clk),
    .D(_04342_),
    .Q(\datamem.data_ram[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _32921_ (.CLK(clk),
    .D(_04343_),
    .Q(\datamem.data_ram[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _32922_ (.CLK(clk),
    .D(_04344_),
    .Q(\datamem.data_ram[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _32923_ (.CLK(clk),
    .D(_04345_),
    .Q(\datamem.data_ram[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _32924_ (.CLK(clk),
    .D(_04346_),
    .Q(\datamem.data_ram[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _32925_ (.CLK(clk),
    .D(_04347_),
    .Q(\datamem.data_ram[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _32926_ (.CLK(clk),
    .D(_04348_),
    .Q(\datamem.data_ram[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _32927_ (.CLK(clk),
    .D(_04349_),
    .Q(\datamem.data_ram[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _32928_ (.CLK(clk),
    .D(_04350_),
    .Q(\datamem.data_ram[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _32929_ (.CLK(clk),
    .D(_04351_),
    .Q(\datamem.data_ram[7][16] ));
 sky130_fd_sc_hd__dfxtp_1 _32930_ (.CLK(clk),
    .D(_04352_),
    .Q(\datamem.data_ram[7][17] ));
 sky130_fd_sc_hd__dfxtp_1 _32931_ (.CLK(clk),
    .D(_04353_),
    .Q(\datamem.data_ram[7][18] ));
 sky130_fd_sc_hd__dfxtp_1 _32932_ (.CLK(clk),
    .D(_04354_),
    .Q(\datamem.data_ram[7][19] ));
 sky130_fd_sc_hd__dfxtp_1 _32933_ (.CLK(clk),
    .D(_04355_),
    .Q(\datamem.data_ram[7][20] ));
 sky130_fd_sc_hd__dfxtp_1 _32934_ (.CLK(clk),
    .D(_04356_),
    .Q(\datamem.data_ram[7][21] ));
 sky130_fd_sc_hd__dfxtp_1 _32935_ (.CLK(clk),
    .D(_04357_),
    .Q(\datamem.data_ram[7][22] ));
 sky130_fd_sc_hd__dfxtp_1 _32936_ (.CLK(clk),
    .D(_04358_),
    .Q(\datamem.data_ram[7][23] ));
 sky130_fd_sc_hd__dfxtp_1 _32937_ (.CLK(clk),
    .D(_04359_),
    .Q(\datamem.data_ram[6][16] ));
 sky130_fd_sc_hd__dfxtp_1 _32938_ (.CLK(clk),
    .D(_04360_),
    .Q(\datamem.data_ram[6][17] ));
 sky130_fd_sc_hd__dfxtp_1 _32939_ (.CLK(clk),
    .D(_04361_),
    .Q(\datamem.data_ram[6][18] ));
 sky130_fd_sc_hd__dfxtp_1 _32940_ (.CLK(clk),
    .D(_04362_),
    .Q(\datamem.data_ram[6][19] ));
 sky130_fd_sc_hd__dfxtp_1 _32941_ (.CLK(clk),
    .D(_04363_),
    .Q(\datamem.data_ram[6][20] ));
 sky130_fd_sc_hd__dfxtp_1 _32942_ (.CLK(clk),
    .D(_04364_),
    .Q(\datamem.data_ram[6][21] ));
 sky130_fd_sc_hd__dfxtp_1 _32943_ (.CLK(clk),
    .D(_04365_),
    .Q(\datamem.data_ram[6][22] ));
 sky130_fd_sc_hd__dfxtp_1 _32944_ (.CLK(clk),
    .D(_04366_),
    .Q(\datamem.data_ram[6][23] ));
 sky130_fd_sc_hd__dfxtp_1 _32945_ (.CLK(clk),
    .D(_04367_),
    .Q(\datamem.data_ram[6][24] ));
 sky130_fd_sc_hd__dfxtp_1 _32946_ (.CLK(clk),
    .D(_04368_),
    .Q(\datamem.data_ram[6][25] ));
 sky130_fd_sc_hd__dfxtp_1 _32947_ (.CLK(clk),
    .D(_04369_),
    .Q(\datamem.data_ram[6][26] ));
 sky130_fd_sc_hd__dfxtp_1 _32948_ (.CLK(clk),
    .D(_04370_),
    .Q(\datamem.data_ram[6][27] ));
 sky130_fd_sc_hd__dfxtp_1 _32949_ (.CLK(clk),
    .D(_04371_),
    .Q(\datamem.data_ram[6][28] ));
 sky130_fd_sc_hd__dfxtp_1 _32950_ (.CLK(clk),
    .D(_04372_),
    .Q(\datamem.data_ram[6][29] ));
 sky130_fd_sc_hd__dfxtp_1 _32951_ (.CLK(clk),
    .D(_04373_),
    .Q(\datamem.data_ram[6][30] ));
 sky130_fd_sc_hd__dfxtp_1 _32952_ (.CLK(clk),
    .D(_04374_),
    .Q(\datamem.data_ram[6][31] ));
 sky130_fd_sc_hd__dfxtp_1 _32953_ (.CLK(clk),
    .D(_04375_),
    .Q(\datamem.data_ram[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _32954_ (.CLK(clk),
    .D(_04376_),
    .Q(\datamem.data_ram[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _32955_ (.CLK(clk),
    .D(_04377_),
    .Q(\datamem.data_ram[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _32956_ (.CLK(clk),
    .D(_04378_),
    .Q(\datamem.data_ram[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _32957_ (.CLK(clk),
    .D(_04379_),
    .Q(\datamem.data_ram[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _32958_ (.CLK(clk),
    .D(_04380_),
    .Q(\datamem.data_ram[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _32959_ (.CLK(clk),
    .D(_04381_),
    .Q(\datamem.data_ram[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _32960_ (.CLK(clk),
    .D(_04382_),
    .Q(\datamem.data_ram[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _32961_ (.CLK(clk),
    .D(_04383_),
    .Q(\datamem.data_ram[63][24] ));
 sky130_fd_sc_hd__dfxtp_1 _32962_ (.CLK(clk),
    .D(_04384_),
    .Q(\datamem.data_ram[63][25] ));
 sky130_fd_sc_hd__dfxtp_1 _32963_ (.CLK(clk),
    .D(_04385_),
    .Q(\datamem.data_ram[63][26] ));
 sky130_fd_sc_hd__dfxtp_1 _32964_ (.CLK(clk),
    .D(_04386_),
    .Q(\datamem.data_ram[63][27] ));
 sky130_fd_sc_hd__dfxtp_1 _32965_ (.CLK(clk),
    .D(_04387_),
    .Q(\datamem.data_ram[63][28] ));
 sky130_fd_sc_hd__dfxtp_1 _32966_ (.CLK(clk),
    .D(_04388_),
    .Q(\datamem.data_ram[63][29] ));
 sky130_fd_sc_hd__dfxtp_1 _32967_ (.CLK(clk),
    .D(_04389_),
    .Q(\datamem.data_ram[63][30] ));
 sky130_fd_sc_hd__dfxtp_1 _32968_ (.CLK(clk),
    .D(_04390_),
    .Q(\datamem.data_ram[63][31] ));
 sky130_fd_sc_hd__dfxtp_1 _32969_ (.CLK(clk),
    .D(_04391_),
    .Q(\datamem.data_ram[63][16] ));
 sky130_fd_sc_hd__dfxtp_1 _32970_ (.CLK(clk),
    .D(_04392_),
    .Q(\datamem.data_ram[63][17] ));
 sky130_fd_sc_hd__dfxtp_1 _32971_ (.CLK(clk),
    .D(_04393_),
    .Q(\datamem.data_ram[63][18] ));
 sky130_fd_sc_hd__dfxtp_1 _32972_ (.CLK(clk),
    .D(_04394_),
    .Q(\datamem.data_ram[63][19] ));
 sky130_fd_sc_hd__dfxtp_1 _32973_ (.CLK(clk),
    .D(_04395_),
    .Q(\datamem.data_ram[63][20] ));
 sky130_fd_sc_hd__dfxtp_1 _32974_ (.CLK(clk),
    .D(_04396_),
    .Q(\datamem.data_ram[63][21] ));
 sky130_fd_sc_hd__dfxtp_1 _32975_ (.CLK(clk),
    .D(_04397_),
    .Q(\datamem.data_ram[63][22] ));
 sky130_fd_sc_hd__dfxtp_1 _32976_ (.CLK(clk),
    .D(_04398_),
    .Q(\datamem.data_ram[63][23] ));
 sky130_fd_sc_hd__dfxtp_1 _32977_ (.CLK(clk),
    .D(_04399_),
    .Q(\datamem.data_ram[63][8] ));
 sky130_fd_sc_hd__dfxtp_1 _32978_ (.CLK(clk),
    .D(_04400_),
    .Q(\datamem.data_ram[63][9] ));
 sky130_fd_sc_hd__dfxtp_1 _32979_ (.CLK(clk),
    .D(_04401_),
    .Q(\datamem.data_ram[63][10] ));
 sky130_fd_sc_hd__dfxtp_1 _32980_ (.CLK(clk),
    .D(_04402_),
    .Q(\datamem.data_ram[63][11] ));
 sky130_fd_sc_hd__dfxtp_1 _32981_ (.CLK(clk),
    .D(_04403_),
    .Q(\datamem.data_ram[63][12] ));
 sky130_fd_sc_hd__dfxtp_1 _32982_ (.CLK(clk),
    .D(_04404_),
    .Q(\datamem.data_ram[63][13] ));
 sky130_fd_sc_hd__dfxtp_1 _32983_ (.CLK(clk),
    .D(_04405_),
    .Q(\datamem.data_ram[63][14] ));
 sky130_fd_sc_hd__dfxtp_1 _32984_ (.CLK(clk),
    .D(_04406_),
    .Q(\datamem.data_ram[63][15] ));
 sky130_fd_sc_hd__dfxtp_1 _32985_ (.CLK(clk),
    .D(_04407_),
    .Q(\datamem.data_ram[62][24] ));
 sky130_fd_sc_hd__dfxtp_1 _32986_ (.CLK(clk),
    .D(_04408_),
    .Q(\datamem.data_ram[62][25] ));
 sky130_fd_sc_hd__dfxtp_1 _32987_ (.CLK(clk),
    .D(_04409_),
    .Q(\datamem.data_ram[62][26] ));
 sky130_fd_sc_hd__dfxtp_1 _32988_ (.CLK(clk),
    .D(_04410_),
    .Q(\datamem.data_ram[62][27] ));
 sky130_fd_sc_hd__dfxtp_1 _32989_ (.CLK(clk),
    .D(_04411_),
    .Q(\datamem.data_ram[62][28] ));
 sky130_fd_sc_hd__dfxtp_1 _32990_ (.CLK(clk),
    .D(_04412_),
    .Q(\datamem.data_ram[62][29] ));
 sky130_fd_sc_hd__dfxtp_1 _32991_ (.CLK(clk),
    .D(_04413_),
    .Q(\datamem.data_ram[62][30] ));
 sky130_fd_sc_hd__dfxtp_1 _32992_ (.CLK(clk),
    .D(_04414_),
    .Q(\datamem.data_ram[62][31] ));
 sky130_fd_sc_hd__buf_1 _32994_ (.A(net13),
    .X(net2));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Right_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Right_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Right_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Right_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Right_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Right_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Right_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Right_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Right_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Right_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Right_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Right_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Right_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Right_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Right_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Right_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Right_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Right_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Right_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Right_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Right_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Right_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Right_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Right_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Right_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Right_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Right_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Right_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Right_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Right_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Right_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Right_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Right_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Right_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Right_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Right_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Right_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Right_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Right_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Right_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Right_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Right_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Right_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Right_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Right_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Right_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Right_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Right_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Right_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Right_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Right_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_Right_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_Right_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_Right_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_Right_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_Right_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_Right_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_Right_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_Right_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_Right_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_Right_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_Right_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_Right_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_Right_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_Right_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_Right_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_Right_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_Right_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_Right_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_171_Right_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_172_Right_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_173_Right_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_174_Right_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_175_Right_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_176_Right_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_177_Right_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_178_Right_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_179_Right_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_180_Right_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_181_Right_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_182_Right_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_183_Right_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_184_Right_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_185_Right_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_186_Right_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_187_Right_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_188_Right_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_189_Right_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_190_Right_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_191_Right_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_192_Right_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_193_Right_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_194_Right_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_195_Right_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_196_Right_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_197_Right_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_198_Right_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_199_Right_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_200_Right_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_201_Right_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_202_Right_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_203_Right_203 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_204_Right_204 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_205_Right_205 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_206_Right_206 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_207_Right_207 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_208_Right_208 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_209_Right_209 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_210_Right_210 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_211_Right_211 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_212_Right_212 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_213_Right_213 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_214_Right_214 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_215_Right_215 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_216_Right_216 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_217_Right_217 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_218_Right_218 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_219_Right_219 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_220_Right_220 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_221_Right_221 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_222_Right_222 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_223_Right_223 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_224_Right_224 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_225_Right_225 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_226_Right_226 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_227_Right_227 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_228_Right_228 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_229_Right_229 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_230 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_231 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_232 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_233 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_234 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_235 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_236 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_237 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_238 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_239 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_240 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_241 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_242 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_243 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_244 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_245 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_246 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_247 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_248 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_249 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_250 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_251 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_252 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_253 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_254 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_255 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_256 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_257 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_258 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_259 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_260 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_261 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_262 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_263 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_264 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_265 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_266 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_267 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_268 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_269 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_270 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_271 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_272 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_273 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_274 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_275 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_276 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_277 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_278 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_279 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_280 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_281 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_282 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_283 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_284 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_285 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_286 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_287 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_288 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_289 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_290 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_291 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_292 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_293 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_294 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_295 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_296 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_297 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_298 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_299 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_300 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_301 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_302 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_303 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_304 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_305 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_306 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_307 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_308 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_309 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_310 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_311 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_312 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_313 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_314 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_315 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_316 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_317 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_318 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_319 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_320 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_321 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_322 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_323 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_324 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_325 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_326 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_327 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_328 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_329 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_330 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_331 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Left_332 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Left_333 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Left_334 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Left_335 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Left_336 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Left_337 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Left_338 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Left_339 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Left_340 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Left_341 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Left_342 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Left_343 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Left_344 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Left_345 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Left_346 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Left_347 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Left_348 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Left_349 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Left_350 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Left_351 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Left_352 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Left_353 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Left_354 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Left_355 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Left_356 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Left_357 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Left_358 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Left_359 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Left_360 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Left_361 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Left_362 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Left_363 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Left_364 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Left_365 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Left_366 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Left_367 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Left_368 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Left_369 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Left_370 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Left_371 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Left_372 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Left_373 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Left_374 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Left_375 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Left_376 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Left_377 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Left_378 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Left_379 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Left_380 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Left_381 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Left_382 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_Left_383 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_Left_384 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_Left_385 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_Left_386 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_Left_387 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_Left_388 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_Left_389 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_Left_390 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_Left_391 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_Left_392 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_Left_393 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_Left_394 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_Left_395 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_Left_396 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_Left_397 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_Left_398 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_Left_399 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_Left_400 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_171_Left_401 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_172_Left_402 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_173_Left_403 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_174_Left_404 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_175_Left_405 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_176_Left_406 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_177_Left_407 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_178_Left_408 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_179_Left_409 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_180_Left_410 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_181_Left_411 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_182_Left_412 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_183_Left_413 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_184_Left_414 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_185_Left_415 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_186_Left_416 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_187_Left_417 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_188_Left_418 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_189_Left_419 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_190_Left_420 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_191_Left_421 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_192_Left_422 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_193_Left_423 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_194_Left_424 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_195_Left_425 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_196_Left_426 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_197_Left_427 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_198_Left_428 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_199_Left_429 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_200_Left_430 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_201_Left_431 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_202_Left_432 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_203_Left_433 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_204_Left_434 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_205_Left_435 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_206_Left_436 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_207_Left_437 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_208_Left_438 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_209_Left_439 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_210_Left_440 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_211_Left_441 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_212_Left_442 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_213_Left_443 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_214_Left_444 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_215_Left_445 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_216_Left_446 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_217_Left_447 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_218_Left_448 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_219_Left_449 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_220_Left_450 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_221_Left_451 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_222_Left_452 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_223_Left_453 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_224_Left_454 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_225_Left_455 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_226_Left_456 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_227_Left_457 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_228_Left_458 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_229_Left_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6027 ();
 sky130_fd_sc_hd__buf_4 input1 (.A(reset),
    .X(net1));
 sky130_fd_sc_hd__buf_2 output2 (.A(net2),
    .X(Instr[0]));
 sky130_fd_sc_hd__buf_2 output3 (.A(net3),
    .X(Instr[10]));
 sky130_fd_sc_hd__buf_2 output4 (.A(net4),
    .X(Instr[11]));
 sky130_fd_sc_hd__buf_2 output5 (.A(net5),
    .X(Instr[12]));
 sky130_fd_sc_hd__buf_2 output6 (.A(net6),
    .X(Instr[13]));
 sky130_fd_sc_hd__buf_2 output7 (.A(net7),
    .X(Instr[14]));
 sky130_fd_sc_hd__buf_2 output8 (.A(net8),
    .X(Instr[15]));
 sky130_fd_sc_hd__buf_2 output9 (.A(net9),
    .X(Instr[16]));
 sky130_fd_sc_hd__buf_2 output10 (.A(net10),
    .X(Instr[17]));
 sky130_fd_sc_hd__buf_2 output11 (.A(net11),
    .X(Instr[18]));
 sky130_fd_sc_hd__buf_2 output12 (.A(net12),
    .X(Instr[19]));
 sky130_fd_sc_hd__buf_2 output13 (.A(net13),
    .X(Instr[1]));
 sky130_fd_sc_hd__buf_2 output14 (.A(net14),
    .X(Instr[20]));
 sky130_fd_sc_hd__buf_2 output15 (.A(net15),
    .X(Instr[21]));
 sky130_fd_sc_hd__buf_2 output16 (.A(net16),
    .X(Instr[22]));
 sky130_fd_sc_hd__buf_2 output17 (.A(net17),
    .X(Instr[23]));
 sky130_fd_sc_hd__buf_2 output18 (.A(net18),
    .X(Instr[24]));
 sky130_fd_sc_hd__buf_2 output19 (.A(net19),
    .X(Instr[25]));
 sky130_fd_sc_hd__buf_2 output20 (.A(net20),
    .X(Instr[26]));
 sky130_fd_sc_hd__buf_2 output21 (.A(net21),
    .X(Instr[27]));
 sky130_fd_sc_hd__buf_2 output22 (.A(net22),
    .X(Instr[28]));
 sky130_fd_sc_hd__buf_2 output23 (.A(net23),
    .X(Instr[29]));
 sky130_fd_sc_hd__buf_2 output24 (.A(net24),
    .X(Instr[2]));
 sky130_fd_sc_hd__buf_2 output25 (.A(net25),
    .X(Instr[30]));
 sky130_fd_sc_hd__buf_2 output26 (.A(net26),
    .X(Instr[31]));
 sky130_fd_sc_hd__buf_2 output27 (.A(net27),
    .X(Instr[3]));
 sky130_fd_sc_hd__buf_2 output28 (.A(net28),
    .X(Instr[4]));
 sky130_fd_sc_hd__buf_2 output29 (.A(net29),
    .X(Instr[5]));
 sky130_fd_sc_hd__buf_2 output30 (.A(net30),
    .X(Instr[6]));
 sky130_fd_sc_hd__buf_2 output31 (.A(net31),
    .X(Instr[7]));
 sky130_fd_sc_hd__buf_2 output32 (.A(net32),
    .X(Instr[8]));
 sky130_fd_sc_hd__buf_2 output33 (.A(net33),
    .X(Instr[9]));
 sky130_fd_sc_hd__buf_2 output34 (.A(net113),
    .X(correct));
 sky130_fd_sc_hd__buf_2 max_cap35 (.A(_10995_),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_4 wire36 (.A(_07964_),
    .X(net36));
 sky130_fd_sc_hd__buf_2 wire37 (.A(_07505_),
    .X(net37));
 sky130_fd_sc_hd__buf_1 wire38 (.A(_06472_),
    .X(net38));
 sky130_fd_sc_hd__buf_4 max_cap39 (.A(_13085_),
    .X(net39));
 sky130_fd_sc_hd__buf_4 max_cap40 (.A(_13058_),
    .X(net40));
 sky130_fd_sc_hd__buf_4 wire41 (.A(_12868_),
    .X(net41));
 sky130_fd_sc_hd__buf_4 wire42 (.A(_12841_),
    .X(net42));
 sky130_fd_sc_hd__buf_4 max_cap43 (.A(_12735_),
    .X(net43));
 sky130_fd_sc_hd__buf_4 max_cap44 (.A(_12592_),
    .X(net44));
 sky130_fd_sc_hd__buf_4 max_cap45 (.A(_12574_),
    .X(net45));
 sky130_fd_sc_hd__buf_4 max_cap46 (.A(_12564_),
    .X(net46));
 sky130_fd_sc_hd__buf_4 wire47 (.A(_12403_),
    .X(net47));
 sky130_fd_sc_hd__buf_4 max_cap48 (.A(_12316_),
    .X(net48));
 sky130_fd_sc_hd__buf_4 max_cap49 (.A(_12298_),
    .X(net49));
 sky130_fd_sc_hd__buf_4 max_cap50 (.A(_12289_),
    .X(net50));
 sky130_fd_sc_hd__buf_4 max_cap51 (.A(_12270_),
    .X(net51));
 sky130_fd_sc_hd__buf_2 max_cap52 (.A(_12041_),
    .X(net52));
 sky130_fd_sc_hd__buf_4 wire53 (.A(_11066_),
    .X(net53));
 sky130_fd_sc_hd__buf_4 max_cap54 (.A(_11021_),
    .X(net54));
 sky130_fd_sc_hd__buf_4 max_cap55 (.A(_10857_),
    .X(net55));
 sky130_fd_sc_hd__buf_4 max_cap56 (.A(_10839_),
    .X(net56));
 sky130_fd_sc_hd__buf_4 max_cap57 (.A(_10829_),
    .X(net57));
 sky130_fd_sc_hd__buf_4 wire58 (.A(_10812_),
    .X(net58));
 sky130_fd_sc_hd__buf_4 max_cap59 (.A(_10561_),
    .X(net59));
 sky130_fd_sc_hd__buf_4 max_cap60 (.A(_10466_),
    .X(net60));
 sky130_fd_sc_hd__buf_4 max_cap61 (.A(_10357_),
    .X(net61));
 sky130_fd_sc_hd__buf_4 wire62 (.A(_09341_),
    .X(net62));
 sky130_fd_sc_hd__buf_4 max_cap63 (.A(_13103_),
    .X(net63));
 sky130_fd_sc_hd__buf_4 max_cap64 (.A(_13094_),
    .X(net64));
 sky130_fd_sc_hd__buf_4 max_cap65 (.A(_13040_),
    .X(net65));
 sky130_fd_sc_hd__buf_4 max_cap66 (.A(_13020_),
    .X(net66));
 sky130_fd_sc_hd__buf_4 max_cap67 (.A(_12978_),
    .X(net67));
 sky130_fd_sc_hd__buf_4 wire68 (.A(_12950_),
    .X(net68));
 sky130_fd_sc_hd__buf_4 max_cap69 (.A(_12923_),
    .X(net69));
 sky130_fd_sc_hd__buf_4 max_cap70 (.A(_12896_),
    .X(net70));
 sky130_fd_sc_hd__buf_4 max_cap71 (.A(_12814_),
    .X(net71));
 sky130_fd_sc_hd__buf_4 max_cap72 (.A(_12623_),
    .X(net72));
 sky130_fd_sc_hd__buf_4 max_cap73 (.A(_12537_),
    .X(net73));
 sky130_fd_sc_hd__buf_4 max_cap74 (.A(_12519_),
    .X(net74));
 sky130_fd_sc_hd__buf_4 max_cap75 (.A(_12510_),
    .X(net75));
 sky130_fd_sc_hd__buf_4 max_cap76 (.A(_12448_),
    .X(net76));
 sky130_fd_sc_hd__buf_4 max_cap77 (.A(_12382_),
    .X(net77));
 sky130_fd_sc_hd__buf_4 wire78 (.A(_12346_),
    .X(net78));
 sky130_fd_sc_hd__buf_4 max_cap79 (.A(_12261_),
    .X(net79));
 sky130_fd_sc_hd__buf_4 max_cap80 (.A(_12242_),
    .X(net80));
 sky130_fd_sc_hd__buf_4 max_cap81 (.A(_12233_),
    .X(net81));
 sky130_fd_sc_hd__buf_4 wire82 (.A(_12215_),
    .X(net82));
 sky130_fd_sc_hd__buf_4 max_cap83 (.A(_12159_),
    .X(net83));
 sky130_fd_sc_hd__buf_4 max_cap84 (.A(_12143_),
    .X(net84));
 sky130_fd_sc_hd__buf_4 max_cap85 (.A(_12116_),
    .X(net85));
 sky130_fd_sc_hd__buf_4 max_cap86 (.A(_12107_),
    .X(net86));
 sky130_fd_sc_hd__buf_4 max_cap87 (.A(_10793_),
    .X(net87));
 sky130_fd_sc_hd__buf_4 max_cap88 (.A(_10784_),
    .X(net88));
 sky130_fd_sc_hd__buf_4 max_cap89 (.A(_10768_),
    .X(net89));
 sky130_fd_sc_hd__buf_4 wire90 (.A(_10742_),
    .X(net90));
 sky130_fd_sc_hd__buf_4 wire91 (.A(_10678_),
    .X(net91));
 sky130_fd_sc_hd__buf_4 max_cap92 (.A(_10650_),
    .X(net92));
 sky130_fd_sc_hd__buf_4 max_cap93 (.A(_10641_),
    .X(net93));
 sky130_fd_sc_hd__buf_4 wire94 (.A(_10602_),
    .X(net94));
 sky130_fd_sc_hd__buf_4 max_cap95 (.A(_12650_),
    .X(net95));
 sky130_fd_sc_hd__buf_4 max_cap96 (.A(_12483_),
    .X(net96));
 sky130_fd_sc_hd__buf_4 max_cap97 (.A(_12464_),
    .X(net97));
 sky130_fd_sc_hd__buf_4 max_cap98 (.A(_12206_),
    .X(net98));
 sky130_fd_sc_hd__buf_4 max_cap99 (.A(_12188_),
    .X(net99));
 sky130_fd_sc_hd__buf_4 max_cap100 (.A(_10725_),
    .X(net100));
 sky130_fd_sc_hd__buf_4 wire101 (.A(_10706_),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_2 max_cap102 (.A(_05429_),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_2 max_cap103 (.A(_05408_),
    .X(net103));
 sky130_fd_sc_hd__buf_8 max_cap104 (.A(_09228_),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_2 max_cap105 (.A(_05307_),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_2 max_cap106 (.A(net111),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_2 max_cap107 (.A(net108),
    .X(net107));
 sky130_fd_sc_hd__buf_2 wire108 (.A(net109),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_2 max_cap109 (.A(net110),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_2 max_cap110 (.A(net111),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_2 max_cap111 (.A(_09300_),
    .X(net111));
 sky130_fd_sc_hd__buf_8 load_slew112 (.A(_09268_),
    .X(net112));
 sky130_fd_sc_hd__buf_1 wire113 (.A(net34),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_2 max_cap114 (.A(net115),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_2 wire115 (.A(_05171_),
    .X(net115));
 sky130_fd_sc_hd__buf_1 max_cap116 (.A(_11377_),
    .X(net116));
 sky130_fd_sc_hd__buf_1 max_cap117 (.A(_08470_),
    .X(net117));
 sky130_fd_sc_hd__buf_2 fanout118 (.A(_00000_),
    .X(net118));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout119 (.A(_00000_),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_2 fanout120 (.A(_00000_),
    .X(net120));
 sky130_fd_sc_hd__buf_1 fanout121 (.A(_00000_),
    .X(net121));
 sky130_fd_sc_hd__buf_12 max_cap122 (.A(\rvcpu.dp.plem.ALUResultM[2] ),
    .X(net122));
 sky130_fd_sc_hd__conb_1 _31746__123 (.LO(net123));
 sky130_fd_sc_hd__conb_1 _31747__124 (.LO(net124));
 sky130_fd_sc_hd__conb_1 _31748__125 (.LO(net125));
 sky130_fd_sc_hd__conb_1 _31749__126 (.LO(net126));
endmodule
